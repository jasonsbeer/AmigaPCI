-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 14 2025 17:39:38

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    TM : in std_logic_vector(1 downto 0);
    TT : in std_logic_vector(1 downto 0);
    D : out std_logic_vector(7 downto 0);
    A : in std_logic_vector(31 downto 1);
    TICK60 : out std_logic;
    CIACS0n : out std_logic;
    CLK6 : in std_logic;
    CLK_CIA : out std_logic;
    BUFENn : out std_logic;
    CIACS1n : out std_logic;
    TICK50 : out std_logic;
    RAMSPACEn : out std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    REGSPACEn : out std_logic;
    TSn : in std_logic;
    RTC_ENn : out std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    TACKn : inout std_logic;
    ROMENn : out std_logic;
    PORTSIZE : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__7448\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2857\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_28\ : std_logic;
signal \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_7_cascade_\ : std_logic;
signal \A_c_29\ : std_logic;
signal \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_8\ : std_logic;
signal \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_9_cascade_\ : std_logic;
signal \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_10\ : std_logic;
signal \N_31_i\ : std_logic;
signal \A_c_31\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_25\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_8_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_10\ : std_logic;
signal \N_69_i\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_13\ : std_logic;
signal \N_101_cascade_\ : std_logic;
signal \N_105\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_17\ : std_logic;
signal \N_74_1_cascade_\ : std_logic;
signal \N_33_cascade_\ : std_logic;
signal \N_99\ : std_logic;
signal \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_5\ : std_logic;
signal \N_99_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_4\ : std_logic;
signal \A_c_18\ : std_logic;
signal \N_74_1\ : std_logic;
signal \N_101\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_9\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U409_ADDRESS_DECODE.HIROMZ0Z_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_94\ : std_logic;
signal \U409_DATA_BUFFERS.un1_BUFENn_iZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_\ : std_logic;
signal \CIA_SPACE_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.N_69\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \U409_ADDRESS_DECODE.un5_RAMSPACEn_cascade_\ : std_logic;
signal \A_c_21\ : std_logic;
signal \A_c_23\ : std_logic;
signal \A_c_22\ : std_logic;
signal \TM_c_0\ : std_logic;
signal \U409_ADDRESS_DECODE_HIROM\ : std_logic;
signal \U409_ADDRESS_DECODE_LOWROM_cascade_\ : std_logic;
signal \TM_c_1\ : std_logic;
signal \N_107\ : std_logic;
signal \N_33\ : std_logic;
signal \N_68_i\ : std_logic;
signal \U409_TRANSFER_ACK.N_71\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \N_67_i\ : std_logic;
signal \N_100\ : std_logic;
signal \OVL_c\ : std_logic;
signal \N_67\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_106\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER15Z0Z_1\ : std_logic;
signal \U409_ADDRESS_DECODE_Z2_SPACE\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\ : std_logic;
signal \ROMENn_c\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_EN_iC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_70_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_55\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U409_TRANSFER_ACK.CO1\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_EN_e_1\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_17_mux\ : std_logic;
signal \U409_TRANSFER_ACK.N_3_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_3_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_6_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \TSn_c\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \U409_TRANSFER_ACK.N_70\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \CIA_ENABLE\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_0C_net\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U409_TICK.TICK603_8_cascade_\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \bfn_15_3_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \bfn_15_4_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \bfn_15_6_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_6\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_7\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_2_0_a4_1_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_6\ : std_logic;
signal \U409_CIA.CLK_CIA_RNOZ0Z_1_cascade_\ : std_logic;
signal \CLK_CIA_c\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_3_0_a4_0_cascade_\ : std_logic;
signal \CIA_SPACE\ : std_logic;
signal \U409_CIA.VMA_RNOZ0Z_0_cascade_\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a4_2_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CLK_CIA6_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CLK_CIA6_1_cascade_\ : std_logic;
signal \U409_CIA.N_104\ : std_logic;
signal \U409_CIA.CLK_CIA6\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \TACK_EN_i\ : std_logic;
signal \N_465_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \D_wire\ : std_logic_vector(7 downto 0);
signal \RTC_ENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \TM_wire\ : std_logic_vector(1 downto 0);
signal \CLK_CIA_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    \TT_wire\ <= TT;
    D <= \D_wire\;
    RTC_ENn <= \RTC_ENn_wire\;
    \A_wire\ <= A;
    \TM_wire\ <= TM;
    CLK_CIA <= \CLK_CIA_wire\;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    \TSn_wire\ <= TSn;
    BUFENn <= \BUFENn_wire\;
    PORTSIZE <= \PORTSIZE_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TICK60 <= \TICK60_wire\;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__4882\,
            RESETB => \N__4759\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__7446\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7448\,
            DIN => \N__7447\,
            DOUT => \N__7446\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7448\,
            PADOUT => \N__7447\,
            PADIN => \N__7446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__7436\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7438\,
            DIN => \N__7437\,
            DOUT => \N__7436\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7438\,
            PADOUT => \N__7437\,
            PADIN => \N__7436\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7427\,
            DIN => \N__7426\,
            DOUT => \N__7425\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7427\,
            PADOUT => \N__7426\,
            PADIN => \N__7425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7418\,
            DIN => \N__7417\,
            DOUT => \N__7416\,
            PACKAGEPIN => \D_wire\(6)
        );

    \D_obuft_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7418\,
            PADOUT => \N__7417\,
            PADIN => \N__7416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RTC_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7409\,
            DIN => \N__7408\,
            DOUT => \N__7407\,
            PACKAGEPIN => \RTC_ENn_wire\
        );

    \RTC_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7409\,
            PADOUT => \N__7408\,
            PADIN => \N__7407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3226\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7400\,
            DIN => \N__7399\,
            DOUT => \N__7398\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7400\,
            PADOUT => \N__7399\,
            PADIN => \N__7398\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7391\,
            DIN => \N__7390\,
            DOUT => \N__7389\,
            PACKAGEPIN => \D_wire\(5)
        );

    \D_obuft_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7391\,
            PADOUT => \N__7390\,
            PADIN => \N__7389\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7382\,
            DIN => \N__7381\,
            DOUT => \N__7380\,
            PACKAGEPIN => \TM_wire\(1)
        );

    \TM_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7382\,
            PADOUT => \N__7381\,
            PADIN => \N__7380\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7373\,
            DIN => \N__7372\,
            DOUT => \N__7371\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7373\,
            PADOUT => \N__7372\,
            PADIN => \N__7371\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_CIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7364\,
            DIN => \N__7363\,
            DOUT => \N__7362\,
            PACKAGEPIN => \CLK_CIA_wire\
        );

    \CLK_CIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7364\,
            PADOUT => \N__7363\,
            PADIN => \N__7362\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6856\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7355\,
            DIN => \N__7354\,
            DOUT => \N__7353\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7355\,
            PADOUT => \N__7354\,
            PADIN => \N__7353\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7346\,
            DIN => \N__7345\,
            DOUT => \N__7344\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7346\,
            PADOUT => \N__7345\,
            PADIN => \N__7344\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4228\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7337\,
            DIN => \N__7336\,
            DOUT => \N__7335\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7337\,
            PADOUT => \N__7336\,
            PADIN => \N__7335\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6910\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__4519\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7328\,
            DIN => \N__7327\,
            DOUT => \N__7326\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7328\,
            PADOUT => \N__7327\,
            PADIN => \N__7326\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7319\,
            DIN => \N__7318\,
            DOUT => \N__7317\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7319\,
            PADOUT => \N__7318\,
            PADIN => \N__7317\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4348\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7310\,
            DIN => \N__7309\,
            DOUT => \N__7308\,
            PACKAGEPIN => \D_wire\(0)
        );

    \D_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7310\,
            PADOUT => \N__7309\,
            PADIN => \N__7308\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7301\,
            DIN => \N__7300\,
            DOUT => \N__7299\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7301\,
            PADOUT => \N__7300\,
            PADIN => \N__7299\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7292\,
            DIN => \N__7291\,
            DOUT => \N__7290\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7292\,
            PADOUT => \N__7291\,
            PADIN => \N__7290\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7283\,
            DIN => \N__7282\,
            DOUT => \N__7281\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7283\,
            PADOUT => \N__7282\,
            PADIN => \N__7281\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3004\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7274\,
            DIN => \N__7273\,
            DOUT => \N__7272\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7274\,
            PADOUT => \N__7273\,
            PADIN => \N__7272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3949\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7265\,
            DIN => \N__7264\,
            DOUT => \N__7263\,
            PACKAGEPIN => \D_wire\(7)
        );

    \D_obuft_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7265\,
            PADOUT => \N__7264\,
            PADIN => \N__7263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7256\,
            DIN => \N__7255\,
            DOUT => \N__7254\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7256\,
            PADOUT => \N__7255\,
            PADIN => \N__7254\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7247\,
            DIN => \N__7246\,
            DOUT => \N__7245\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7247\,
            PADOUT => \N__7246\,
            PADIN => \N__7245\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7238\,
            DIN => \N__7237\,
            DOUT => \N__7236\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7238\,
            PADOUT => \N__7237\,
            PADIN => \N__7236\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7229\,
            DIN => \N__7228\,
            DOUT => \N__7227\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7229\,
            PADOUT => \N__7228\,
            PADIN => \N__7227\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7220\,
            DIN => \N__7219\,
            DOUT => \N__7218\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7220\,
            PADOUT => \N__7219\,
            PADIN => \N__7218\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7211\,
            DIN => \N__7210\,
            DOUT => \N__7209\,
            PACKAGEPIN => \D_wire\(2)
        );

    \D_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7211\,
            PADOUT => \N__7210\,
            PADIN => \N__7209\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7202\,
            DIN => \N__7201\,
            DOUT => \N__7200\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7202\,
            PADOUT => \N__7201\,
            PADIN => \N__7200\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7193\,
            DIN => \N__7192\,
            DOUT => \N__7191\,
            PACKAGEPIN => \TM_wire\(0)
        );

    \TM_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7193\,
            PADOUT => \N__7192\,
            PADIN => \N__7191\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7184\,
            DIN => \N__7183\,
            DOUT => \N__7182\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7184\,
            PADOUT => \N__7183\,
            PADIN => \N__7182\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7175\,
            DIN => \N__7174\,
            DOUT => \N__7173\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7175\,
            PADOUT => \N__7174\,
            PADIN => \N__7173\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7166\,
            DIN => \N__7165\,
            DOUT => \N__7164\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7166\,
            PADOUT => \N__7165\,
            PADIN => \N__7164\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7157\,
            DIN => \N__7156\,
            DOUT => \N__7155\,
            PACKAGEPIN => \D_wire\(1)
        );

    \D_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7157\,
            PADOUT => \N__7156\,
            PADIN => \N__7155\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7148\,
            DIN => \N__7147\,
            DOUT => \N__7146\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7148\,
            PADOUT => \N__7147\,
            PADIN => \N__7146\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5371\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7139\,
            DIN => \N__7138\,
            DOUT => \N__7137\,
            PACKAGEPIN => \D_wire\(4)
        );

    \D_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7139\,
            PADOUT => \N__7138\,
            PADIN => \N__7137\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7130\,
            DIN => \N__7129\,
            DOUT => \N__7128\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7130\,
            PADOUT => \N__7129\,
            PADIN => \N__7128\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5677\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7121\,
            DIN => \N__7120\,
            DOUT => \N__7119\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7121\,
            PADOUT => \N__7120\,
            PADIN => \N__7119\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7112\,
            DIN => \N__7111\,
            DOUT => \N__7110\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7112\,
            PADOUT => \N__7111\,
            PADIN => \N__7110\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7103\,
            DIN => \N__7102\,
            DOUT => \N__7101\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7103\,
            PADOUT => \N__7102\,
            PADIN => \N__7101\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7094\,
            DIN => \N__7093\,
            DOUT => \N__7092\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7094\,
            PADOUT => \N__7093\,
            PADIN => \N__7092\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7085\,
            DIN => \N__7084\,
            DOUT => \N__7083\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7085\,
            PADOUT => \N__7084\,
            PADIN => \N__7083\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7076\,
            DIN => \N__7075\,
            DOUT => \N__7074\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7076\,
            PADOUT => \N__7075\,
            PADIN => \N__7074\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5806\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7067\,
            DIN => \N__7066\,
            DOUT => \N__7065\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7067\,
            PADOUT => \N__7066\,
            PADIN => \N__7065\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7058\,
            DIN => \N__7057\,
            DOUT => \N__7056\,
            PACKAGEPIN => \D_wire\(3)
        );

    \D_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7058\,
            PADOUT => \N__7057\,
            PADIN => \N__7056\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7049\,
            DIN => \N__7048\,
            DOUT => \N__7047\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7049\,
            PADOUT => \N__7048\,
            PADIN => \N__7047\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7040\,
            DIN => \N__7039\,
            DOUT => \N__7038\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7040\,
            PADOUT => \N__7039\,
            PADIN => \N__7038\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7031\,
            DIN => \N__7030\,
            DOUT => \N__7029\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7031\,
            PADOUT => \N__7030\,
            PADIN => \N__7029\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5410\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7022\,
            DIN => \N__7021\,
            DOUT => \N__7020\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7022\,
            PADOUT => \N__7021\,
            PADIN => \N__7020\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3673\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__7003\,
            I => \N__6998\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6989\
        );

    \I__1630\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6989\
        );

    \I__1629\ : InMux
    port map (
            O => \N__6998\,
            I => \N__6986\
        );

    \I__1628\ : InMux
    port map (
            O => \N__6997\,
            I => \N__6977\
        );

    \I__1627\ : InMux
    port map (
            O => \N__6996\,
            I => \N__6977\
        );

    \I__1626\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6977\
        );

    \I__1625\ : InMux
    port map (
            O => \N__6994\,
            I => \N__6977\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__6989\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__6986\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__6977\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__6970\,
            I => \N__6965\
        );

    \I__1620\ : InMux
    port map (
            O => \N__6969\,
            I => \N__6959\
        );

    \I__1619\ : InMux
    port map (
            O => \N__6968\,
            I => \N__6954\
        );

    \I__1618\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6954\
        );

    \I__1617\ : InMux
    port map (
            O => \N__6964\,
            I => \N__6947\
        );

    \I__1616\ : InMux
    port map (
            O => \N__6963\,
            I => \N__6947\
        );

    \I__1615\ : InMux
    port map (
            O => \N__6962\,
            I => \N__6947\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__6959\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__6954\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__6947\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1611\ : ClkMux
    port map (
            O => \N__6940\,
            I => \N__6931\
        );

    \I__1610\ : ClkMux
    port map (
            O => \N__6939\,
            I => \N__6931\
        );

    \I__1609\ : ClkMux
    port map (
            O => \N__6938\,
            I => \N__6931\
        );

    \I__1608\ : GlobalMux
    port map (
            O => \N__6931\,
            I => \N__6928\
        );

    \I__1607\ : gio2CtrlBuf
    port map (
            O => \N__6928\,
            I => \CLK28_IN_c_g\
        );

    \I__1606\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6922\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__6922\,
            I => \N__6919\
        );

    \I__1604\ : Span4Mux_v
    port map (
            O => \N__6919\,
            I => \N__6916\
        );

    \I__1603\ : Span4Mux_h
    port map (
            O => \N__6916\,
            I => \N__6913\
        );

    \I__1602\ : Odrv4
    port map (
            O => \N__6913\,
            I => \TACK_EN_i\
        );

    \I__1601\ : IoInMux
    port map (
            O => \N__6910\,
            I => \N__6907\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__6907\,
            I => \N__6904\
        );

    \I__1599\ : Span4Mux_s2_v
    port map (
            O => \N__6904\,
            I => \N__6901\
        );

    \I__1598\ : Sp12to4
    port map (
            O => \N__6901\,
            I => \N__6898\
        );

    \I__1597\ : Span12Mux_h
    port map (
            O => \N__6898\,
            I => \N__6895\
        );

    \I__1596\ : Odrv12
    port map (
            O => \N__6895\,
            I => \N_465_i\
        );

    \I__1595\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6887\
        );

    \I__1594\ : InMux
    port map (
            O => \N__6891\,
            I => \N__6882\
        );

    \I__1593\ : InMux
    port map (
            O => \N__6890\,
            I => \N__6882\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__6887\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__6882\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__6877\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_2_0_a4_1_cascade_\
        );

    \I__1589\ : InMux
    port map (
            O => \N__6874\,
            I => \N__6869\
        );

    \I__1588\ : InMux
    port map (
            O => \N__6873\,
            I => \N__6864\
        );

    \I__1587\ : InMux
    port map (
            O => \N__6872\,
            I => \N__6864\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__6869\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__6864\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__6859\,
            I => \U409_CIA.CLK_CIA_RNOZ0Z_1_cascade_\
        );

    \I__1583\ : IoInMux
    port map (
            O => \N__6856\,
            I => \N__6853\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__6853\,
            I => \N__6850\
        );

    \I__1581\ : IoSpan4Mux
    port map (
            O => \N__6850\,
            I => \N__6847\
        );

    \I__1580\ : Span4Mux_s1_v
    port map (
            O => \N__6847\,
            I => \N__6844\
        );

    \I__1579\ : Sp12to4
    port map (
            O => \N__6844\,
            I => \N__6840\
        );

    \I__1578\ : InMux
    port map (
            O => \N__6843\,
            I => \N__6837\
        );

    \I__1577\ : Span12Mux_s9_v
    port map (
            O => \N__6840\,
            I => \N__6833\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__6837\,
            I => \N__6830\
        );

    \I__1575\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6827\
        );

    \I__1574\ : Odrv12
    port map (
            O => \N__6833\,
            I => \CLK_CIA_c\
        );

    \I__1573\ : Odrv4
    port map (
            O => \N__6830\,
            I => \CLK_CIA_c\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__6827\,
            I => \CLK_CIA_c\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__6820\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_3_0_a4_0_cascade_\
        );

    \I__1570\ : InMux
    port map (
            O => \N__6817\,
            I => \N__6814\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__6814\,
            I => \N__6811\
        );

    \I__1568\ : Span4Mux_v
    port map (
            O => \N__6811\,
            I => \N__6808\
        );

    \I__1567\ : Sp12to4
    port map (
            O => \N__6808\,
            I => \N__6805\
        );

    \I__1566\ : Span12Mux_h
    port map (
            O => \N__6805\,
            I => \N__6802\
        );

    \I__1565\ : Odrv12
    port map (
            O => \N__6802\,
            I => \CIA_SPACE\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__6799\,
            I => \U409_CIA.VMA_RNOZ0Z_0_cascade_\
        );

    \I__1563\ : InMux
    port map (
            O => \N__6796\,
            I => \N__6792\
        );

    \I__1562\ : InMux
    port map (
            O => \N__6795\,
            I => \N__6789\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__6792\,
            I => \N__6786\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__6789\,
            I => \N__6783\
        );

    \I__1559\ : Span4Mux_v
    port map (
            O => \N__6786\,
            I => \N__6777\
        );

    \I__1558\ : Span4Mux_v
    port map (
            O => \N__6783\,
            I => \N__6777\
        );

    \I__1557\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6774\
        );

    \I__1556\ : Odrv4
    port map (
            O => \N__6777\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__6774\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1554\ : CascadeMux
    port map (
            O => \N__6769\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a4_2_cascade_\
        );

    \I__1553\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6760\
        );

    \I__1552\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6760\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__6760\,
            I => \U409_CIA.CIA_CLK_COUNT11\
        );

    \I__1550\ : InMux
    port map (
            O => \N__6757\,
            I => \N__6754\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__6754\,
            I => \N__6748\
        );

    \I__1548\ : InMux
    port map (
            O => \N__6753\,
            I => \N__6745\
        );

    \I__1547\ : InMux
    port map (
            O => \N__6752\,
            I => \N__6742\
        );

    \I__1546\ : InMux
    port map (
            O => \N__6751\,
            I => \N__6739\
        );

    \I__1545\ : Odrv4
    port map (
            O => \N__6748\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__6745\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__6742\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__6739\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1541\ : InMux
    port map (
            O => \N__6730\,
            I => \N__6724\
        );

    \I__1540\ : InMux
    port map (
            O => \N__6729\,
            I => \N__6721\
        );

    \I__1539\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6716\
        );

    \I__1538\ : InMux
    port map (
            O => \N__6727\,
            I => \N__6716\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__6724\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__6721\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__6716\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1534\ : InMux
    port map (
            O => \N__6709\,
            I => \N__6706\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__6706\,
            I => \U409_CIA.CLK_CIA6_1\
        );

    \I__1532\ : InMux
    port map (
            O => \N__6703\,
            I => \N__6696\
        );

    \I__1531\ : InMux
    port map (
            O => \N__6702\,
            I => \N__6693\
        );

    \I__1530\ : InMux
    port map (
            O => \N__6701\,
            I => \N__6686\
        );

    \I__1529\ : InMux
    port map (
            O => \N__6700\,
            I => \N__6686\
        );

    \I__1528\ : InMux
    port map (
            O => \N__6699\,
            I => \N__6686\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__6696\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__6693\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__6686\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1524\ : CascadeMux
    port map (
            O => \N__6679\,
            I => \U409_CIA.CLK_CIA6_1_cascade_\
        );

    \I__1523\ : InMux
    port map (
            O => \N__6676\,
            I => \N__6671\
        );

    \I__1522\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6666\
        );

    \I__1521\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6666\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__6671\,
            I => \U409_CIA.N_104\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__6666\,
            I => \U409_CIA.N_104\
        );

    \I__1518\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6658\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__6658\,
            I => \U409_CIA.CLK_CIA6\
        );

    \I__1516\ : InMux
    port map (
            O => \N__6655\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__1515\ : InMux
    port map (
            O => \N__6652\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__1514\ : InMux
    port map (
            O => \N__6649\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__1513\ : InMux
    port map (
            O => \N__6646\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__1512\ : InMux
    port map (
            O => \N__6643\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\
        );

    \I__1511\ : InMux
    port map (
            O => \N__6640\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__6637\,
            I => \N__6633\
        );

    \I__1509\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6629\
        );

    \I__1508\ : InMux
    port map (
            O => \N__6633\,
            I => \N__6624\
        );

    \I__1507\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6624\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__6629\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__6624\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1504\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6615\
        );

    \I__1503\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6612\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__6615\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__6612\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__1500\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6604\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__6604\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__1498\ : InMux
    port map (
            O => \N__6601\,
            I => \bfn_15_4_0_\
        );

    \I__1497\ : InMux
    port map (
            O => \N__6598\,
            I => \N__6594\
        );

    \I__1496\ : InMux
    port map (
            O => \N__6597\,
            I => \N__6591\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__6594\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__6591\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__1493\ : InMux
    port map (
            O => \N__6586\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__1492\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6579\
        );

    \I__1491\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6576\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__6579\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__6576\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__1488\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6568\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__6568\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__1486\ : InMux
    port map (
            O => \N__6565\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__1485\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6558\
        );

    \I__1484\ : InMux
    port map (
            O => \N__6561\,
            I => \N__6555\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__6558\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__6555\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__1481\ : InMux
    port map (
            O => \N__6550\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__1480\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6543\
        );

    \I__1479\ : InMux
    port map (
            O => \N__6546\,
            I => \N__6540\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__6543\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__6540\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1476\ : InMux
    port map (
            O => \N__6535\,
            I => \N__6532\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__6532\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__1474\ : InMux
    port map (
            O => \N__6529\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__1473\ : InMux
    port map (
            O => \N__6526\,
            I => \N__6522\
        );

    \I__1472\ : InMux
    port map (
            O => \N__6525\,
            I => \N__6519\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__6522\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__6519\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__6514\,
            I => \N__6511\
        );

    \I__1468\ : InMux
    port map (
            O => \N__6511\,
            I => \N__6508\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__6508\,
            I => \N__6505\
        );

    \I__1466\ : Odrv4
    port map (
            O => \N__6505\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__1465\ : InMux
    port map (
            O => \N__6502\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__1464\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6495\
        );

    \I__1463\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6492\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__6495\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__6492\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1460\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6484\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__6484\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__1458\ : InMux
    port map (
            O => \N__6481\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__1457\ : InMux
    port map (
            O => \N__6478\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6471\
        );

    \I__1455\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6468\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__6471\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__6468\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__1452\ : ClkMux
    port map (
            O => \N__6463\,
            I => \N__6439\
        );

    \I__1451\ : ClkMux
    port map (
            O => \N__6462\,
            I => \N__6439\
        );

    \I__1450\ : ClkMux
    port map (
            O => \N__6461\,
            I => \N__6439\
        );

    \I__1449\ : ClkMux
    port map (
            O => \N__6460\,
            I => \N__6439\
        );

    \I__1448\ : ClkMux
    port map (
            O => \N__6459\,
            I => \N__6439\
        );

    \I__1447\ : ClkMux
    port map (
            O => \N__6458\,
            I => \N__6439\
        );

    \I__1446\ : ClkMux
    port map (
            O => \N__6457\,
            I => \N__6439\
        );

    \I__1445\ : ClkMux
    port map (
            O => \N__6456\,
            I => \N__6439\
        );

    \I__1444\ : GlobalMux
    port map (
            O => \N__6439\,
            I => \N__6436\
        );

    \I__1443\ : gio2CtrlBuf
    port map (
            O => \N__6436\,
            I => \CLK6_c_g\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__6433\,
            I => \N__6429\
        );

    \I__1441\ : InMux
    port map (
            O => \N__6432\,
            I => \N__6423\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6429\,
            I => \N__6423\
        );

    \I__1439\ : InMux
    port map (
            O => \N__6428\,
            I => \N__6420\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__6423\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__6420\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1436\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6410\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__6414\,
            I => \N__6406\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6413\,
            I => \N__6403\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__6410\,
            I => \N__6400\
        );

    \I__1432\ : InMux
    port map (
            O => \N__6409\,
            I => \N__6397\
        );

    \I__1431\ : InMux
    port map (
            O => \N__6406\,
            I => \N__6394\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6403\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__6400\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__6397\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__6394\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6381\
        );

    \I__1425\ : InMux
    port map (
            O => \N__6384\,
            I => \N__6378\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__6381\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__6378\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6373\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6370\,
            I => \N__6366\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6369\,
            I => \N__6363\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__6366\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__6363\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__1417\ : InMux
    port map (
            O => \N__6358\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__6355\,
            I => \N__6352\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6348\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6351\,
            I => \N__6345\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__6348\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6345\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1411\ : InMux
    port map (
            O => \N__6340\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__6337\,
            I => \N__6333\
        );

    \I__1409\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6330\
        );

    \I__1408\ : InMux
    port map (
            O => \N__6333\,
            I => \N__6327\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__6330\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__6327\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__1404\ : InMux
    port map (
            O => \N__6319\,
            I => \N__6316\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__6316\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6313\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__6310\,
            I => \N__6307\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6303\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6300\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6303\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__6300\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__6295\,
            I => \N__6292\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6292\,
            I => \N__6289\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6289\,
            I => \N__6286\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__6286\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6283\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__1391\ : InMux
    port map (
            O => \N__6280\,
            I => \N__6276\
        );

    \I__1390\ : InMux
    port map (
            O => \N__6279\,
            I => \N__6273\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__6276\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6273\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6268\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__1386\ : InMux
    port map (
            O => \N__6265\,
            I => \N__6261\
        );

    \I__1385\ : InMux
    port map (
            O => \N__6264\,
            I => \N__6258\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__6261\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__6258\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6253\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6250\,
            I => \N__6246\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6243\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6246\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6243\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6235\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__6235\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6232\,
            I => \bfn_14_9_0_\
        );

    \I__1374\ : InMux
    port map (
            O => \N__6229\,
            I => \N__6225\
        );

    \I__1373\ : InMux
    port map (
            O => \N__6228\,
            I => \N__6222\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__6225\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6222\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1370\ : InMux
    port map (
            O => \N__6217\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6210\
        );

    \I__1368\ : InMux
    port map (
            O => \N__6213\,
            I => \N__6207\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__6210\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__6207\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6202\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6195\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6192\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__6195\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6192\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__1360\ : InMux
    port map (
            O => \N__6187\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__1359\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6180\
        );

    \I__1358\ : InMux
    port map (
            O => \N__6183\,
            I => \N__6177\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__6180\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__6177\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6172\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__1354\ : InMux
    port map (
            O => \N__6169\,
            I => \N__6165\
        );

    \I__1353\ : InMux
    port map (
            O => \N__6168\,
            I => \N__6162\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__6165\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6162\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__1350\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6154\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6154\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6151\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6148\,
            I => \N__6144\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6141\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__6144\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__6141\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6136\,
            I => \N__6133\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6133\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6130\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6127\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6124\,
            I => \N__6120\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6123\,
            I => \N__6117\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6120\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__6117\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__1335\ : CascadeMux
    port map (
            O => \N__6112\,
            I => \N__6108\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6104\
        );

    \I__1333\ : InMux
    port map (
            O => \N__6108\,
            I => \N__6101\
        );

    \I__1332\ : InMux
    port map (
            O => \N__6107\,
            I => \N__6098\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__6104\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__6101\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6098\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__6091\,
            I => \N__6087\
        );

    \I__1327\ : CascadeMux
    port map (
            O => \N__6090\,
            I => \N__6082\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6087\,
            I => \N__6079\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6086\,
            I => \N__6076\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6073\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6070\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6079\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6076\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6073\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6070\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6061\,
            I => \N__6057\
        );

    \I__1317\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6054\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6057\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__6054\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6049\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6046\,
            I => \N__6042\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6039\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6042\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6039\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6034\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6027\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6030\,
            I => \N__6024\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6027\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6024\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6019\,
            I => \N__6016\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6016\,
            I => \N__6013\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__6013\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6010\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6007\,
            I => \N__6003\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6006\,
            I => \N__6000\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__6003\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6000\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__1296\ : InMux
    port map (
            O => \N__5995\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__5992\,
            I => \N__5988\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__5991\,
            I => \N__5985\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5988\,
            I => \N__5982\
        );

    \I__1292\ : InMux
    port map (
            O => \N__5985\,
            I => \N__5979\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5982\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__5979\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__1289\ : InMux
    port map (
            O => \N__5974\,
            I => \N__5971\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__5971\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__1287\ : InMux
    port map (
            O => \N__5968\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__5965\,
            I => \N__5962\
        );

    \I__1285\ : InMux
    port map (
            O => \N__5962\,
            I => \N__5959\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__5959\,
            I => \N__5955\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5952\
        );

    \I__1282\ : Odrv4
    port map (
            O => \N__5955\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__5952\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5947\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5940\
        );

    \I__1278\ : InMux
    port map (
            O => \N__5943\,
            I => \N__5937\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5940\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__5937\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__1275\ : InMux
    port map (
            O => \N__5932\,
            I => \N__5929\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5929\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__1273\ : InMux
    port map (
            O => \N__5926\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5923\,
            I => \N__5920\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__5920\,
            I => \U409_TICK.TICK503_11\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__5917\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__5914\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5895\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5910\,
            I => \N__5895\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5909\,
            I => \N__5895\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5908\,
            I => \N__5895\
        );

    \I__1264\ : InMux
    port map (
            O => \N__5907\,
            I => \N__5886\
        );

    \I__1263\ : InMux
    port map (
            O => \N__5906\,
            I => \N__5886\
        );

    \I__1262\ : InMux
    port map (
            O => \N__5905\,
            I => \N__5886\
        );

    \I__1261\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5886\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5895\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5886\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5881\,
            I => \N__5863\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5880\,
            I => \N__5863\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5879\,
            I => \N__5863\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5878\,
            I => \N__5863\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5863\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5856\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5856\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5856\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5863\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5856\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__5851\,
            I => \N__5846\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5850\,
            I => \N__5833\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5849\,
            I => \N__5833\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5846\,
            I => \N__5833\
        );

    \I__1244\ : InMux
    port map (
            O => \N__5845\,
            I => \N__5833\
        );

    \I__1243\ : CascadeMux
    port map (
            O => \N__5844\,
            I => \N__5829\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__5843\,
            I => \N__5826\
        );

    \I__1241\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5823\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__5833\,
            I => \N__5820\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5832\,
            I => \N__5813\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5813\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5826\,
            I => \N__5813\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__5823\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__5820\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5813\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1233\ : IoInMux
    port map (
            O => \N__5806\,
            I => \N__5803\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__5803\,
            I => \N__5800\
        );

    \I__1231\ : Span4Mux_s0_v
    port map (
            O => \N__5800\,
            I => \N__5797\
        );

    \I__1230\ : Span4Mux_v
    port map (
            O => \N__5797\,
            I => \N__5794\
        );

    \I__1229\ : Span4Mux_v
    port map (
            O => \N__5794\,
            I => \N__5791\
        );

    \I__1228\ : Span4Mux_v
    port map (
            O => \N__5791\,
            I => \N__5787\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5790\,
            I => \N__5784\
        );

    \I__1226\ : Odrv4
    port map (
            O => \N__5787\,
            I => \TICK60_c\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__5784\,
            I => \TICK60_c\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__5779\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__5776\,
            I => \N__5770\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__5775\,
            I => \N__5767\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5774\,
            I => \N__5755\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5755\
        );

    \I__1219\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5755\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5755\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5766\,
            I => \N__5748\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5765\,
            I => \N__5748\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5764\,
            I => \N__5748\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__5755\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5748\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__5743\,
            I => \N__5740\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5740\,
            I => \N__5737\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__5737\,
            I => \N__5728\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5736\,
            I => \N__5721\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5735\,
            I => \N__5721\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5721\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5714\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5732\,
            I => \N__5714\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5714\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__5728\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5721\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__5714\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__5707\,
            I => \N__5703\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5689\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5689\
        );

    \I__1197\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5689\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5689\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5700\,
            I => \N__5682\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5682\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5698\,
            I => \N__5682\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5689\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__5682\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1190\ : IoInMux
    port map (
            O => \N__5677\,
            I => \N__5674\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5674\,
            I => \N__5671\
        );

    \I__1188\ : Span4Mux_s1_v
    port map (
            O => \N__5671\,
            I => \N__5668\
        );

    \I__1187\ : Sp12to4
    port map (
            O => \N__5668\,
            I => \N__5665\
        );

    \I__1186\ : Span12Mux_h
    port map (
            O => \N__5665\,
            I => \N__5661\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5658\
        );

    \I__1184\ : Odrv12
    port map (
            O => \N__5661\,
            I => \TICK50_c\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5658\,
            I => \TICK50_c\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__5653\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__1181\ : SRMux
    port map (
            O => \N__5650\,
            I => \N__5646\
        );

    \I__1180\ : SRMux
    port map (
            O => \N__5649\,
            I => \N__5642\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5646\,
            I => \N__5637\
        );

    \I__1178\ : SRMux
    port map (
            O => \N__5645\,
            I => \N__5634\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5642\,
            I => \N__5631\
        );

    \I__1176\ : SRMux
    port map (
            O => \N__5641\,
            I => \N__5628\
        );

    \I__1175\ : SRMux
    port map (
            O => \N__5640\,
            I => \N__5625\
        );

    \I__1174\ : Span4Mux_v
    port map (
            O => \N__5637\,
            I => \N__5621\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5634\,
            I => \N__5618\
        );

    \I__1172\ : Span4Mux_v
    port map (
            O => \N__5631\,
            I => \N__5615\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__5628\,
            I => \N__5612\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5625\,
            I => \N__5609\
        );

    \I__1169\ : SRMux
    port map (
            O => \N__5624\,
            I => \N__5606\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__5621\,
            I => \RESETn_c_i\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__5618\,
            I => \RESETn_c_i\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__5615\,
            I => \RESETn_c_i\
        );

    \I__1165\ : Odrv12
    port map (
            O => \N__5612\,
            I => \RESETn_c_i\
        );

    \I__1164\ : Odrv12
    port map (
            O => \N__5609\,
            I => \RESETn_c_i\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5606\,
            I => \RESETn_c_i\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__5593\,
            I => \U409_TICK.TICK603_8_cascade_\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__5590\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5584\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5584\,
            I => \U409_TICK.TICK603_11\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__5581\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__5578\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__5575\,
            I => \N__5570\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5565\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5573\,
            I => \N__5562\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5570\,
            I => \N__5555\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5569\,
            I => \N__5555\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5568\,
            I => \N__5555\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5565\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5562\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5555\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__5548\,
            I => \N__5541\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5547\,
            I => \N__5536\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5536\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5545\,
            I => \N__5533\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5528\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5528\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5536\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5533\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5528\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5508\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5508\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5519\,
            I => \N__5508\
        );

    \I__1135\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5505\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5502\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5516\,
            I => \N__5497\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5515\,
            I => \N__5497\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__5508\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__5505\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__5502\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5497\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5482\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5479\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5486\,
            I => \N__5474\
        );

    \I__1124\ : InMux
    port map (
            O => \N__5485\,
            I => \N__5474\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__5482\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__5479\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__5474\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1120\ : SRMux
    port map (
            O => \N__5467\,
            I => \N__5463\
        );

    \I__1119\ : SRMux
    port map (
            O => \N__5466\,
            I => \N__5459\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5463\,
            I => \N__5456\
        );

    \I__1117\ : SRMux
    port map (
            O => \N__5462\,
            I => \N__5453\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5459\,
            I => \N__5449\
        );

    \I__1115\ : Span4Mux_v
    port map (
            O => \N__5456\,
            I => \N__5444\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__5453\,
            I => \N__5444\
        );

    \I__1113\ : SRMux
    port map (
            O => \N__5452\,
            I => \N__5441\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__5449\,
            I => \N__5436\
        );

    \I__1111\ : Span4Mux_h
    port map (
            O => \N__5444\,
            I => \N__5436\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5441\,
            I => \N__5433\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__5436\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__5433\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5428\,
            I => \N__5425\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__5425\,
            I => \N__5422\
        );

    \I__1105\ : Span4Mux_v
    port map (
            O => \N__5422\,
            I => \N__5419\
        );

    \I__1104\ : Sp12to4
    port map (
            O => \N__5419\,
            I => \N__5416\
        );

    \I__1103\ : Span12Mux_h
    port map (
            O => \N__5416\,
            I => \N__5413\
        );

    \I__1102\ : Odrv12
    port map (
            O => \N__5413\,
            I => \A_c_13\
        );

    \I__1101\ : IoInMux
    port map (
            O => \N__5410\,
            I => \N__5407\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5407\,
            I => \N__5404\
        );

    \I__1099\ : IoSpan4Mux
    port map (
            O => \N__5404\,
            I => \N__5401\
        );

    \I__1098\ : IoSpan4Mux
    port map (
            O => \N__5401\,
            I => \N__5398\
        );

    \I__1097\ : Sp12to4
    port map (
            O => \N__5398\,
            I => \N__5395\
        );

    \I__1096\ : Span12Mux_s7_h
    port map (
            O => \N__5395\,
            I => \N__5392\
        );

    \I__1095\ : Odrv12
    port map (
            O => \N__5392\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5389\,
            I => \N__5386\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5386\,
            I => \N__5383\
        );

    \I__1092\ : Span4Mux_v
    port map (
            O => \N__5383\,
            I => \N__5380\
        );

    \I__1091\ : Sp12to4
    port map (
            O => \N__5380\,
            I => \N__5377\
        );

    \I__1090\ : Span12Mux_h
    port map (
            O => \N__5377\,
            I => \N__5374\
        );

    \I__1089\ : Odrv12
    port map (
            O => \N__5374\,
            I => \A_c_12\
        );

    \I__1088\ : IoInMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__5368\,
            I => \N__5365\
        );

    \I__1086\ : IoSpan4Mux
    port map (
            O => \N__5365\,
            I => \N__5362\
        );

    \I__1085\ : IoSpan4Mux
    port map (
            O => \N__5362\,
            I => \N__5359\
        );

    \I__1084\ : Span4Mux_s2_h
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__1083\ : Sp12to4
    port map (
            O => \N__5356\,
            I => \N__5353\
        );

    \I__1082\ : Odrv12
    port map (
            O => \N__5353\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__1081\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5344\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5344\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5344\,
            I => \CIA_ENABLE\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__5341\,
            I => \N__5336\
        );

    \I__1077\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5332\
        );

    \I__1076\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5329\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5325\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5322\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5332\,
            I => \N__5319\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5329\,
            I => \N__5316\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5328\,
            I => \N__5313\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__5325\,
            I => \N__5307\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5322\,
            I => \N__5307\
        );

    \I__1068\ : Span4Mux_h
    port map (
            O => \N__5319\,
            I => \N__5304\
        );

    \I__1067\ : Span4Mux_v
    port map (
            O => \N__5316\,
            I => \N__5301\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5313\,
            I => \N__5298\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__5312\,
            I => \N__5295\
        );

    \I__1064\ : Span4Mux_v
    port map (
            O => \N__5307\,
            I => \N__5292\
        );

    \I__1063\ : Span4Mux_h
    port map (
            O => \N__5304\,
            I => \N__5288\
        );

    \I__1062\ : Span4Mux_h
    port map (
            O => \N__5301\,
            I => \N__5283\
        );

    \I__1061\ : Span4Mux_v
    port map (
            O => \N__5298\,
            I => \N__5283\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5295\,
            I => \N__5280\
        );

    \I__1059\ : Span4Mux_h
    port map (
            O => \N__5292\,
            I => \N__5273\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5270\
        );

    \I__1057\ : Span4Mux_h
    port map (
            O => \N__5288\,
            I => \N__5264\
        );

    \I__1056\ : Span4Mux_h
    port map (
            O => \N__5283\,
            I => \N__5259\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__5280\,
            I => \N__5259\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5250\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5278\,
            I => \N__5250\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5277\,
            I => \N__5250\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5250\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__5273\,
            I => \N__5244\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5270\,
            I => \N__5244\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5241\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5238\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5235\
        );

    \I__1045\ : Span4Mux_v
    port map (
            O => \N__5264\,
            I => \N__5232\
        );

    \I__1044\ : Span4Mux_v
    port map (
            O => \N__5259\,
            I => \N__5227\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5250\,
            I => \N__5227\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5249\,
            I => \N__5224\
        );

    \I__1041\ : Span4Mux_h
    port map (
            O => \N__5244\,
            I => \N__5219\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5241\,
            I => \N__5219\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5238\,
            I => \N__5214\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__5235\,
            I => \N__5214\
        );

    \I__1037\ : Sp12to4
    port map (
            O => \N__5232\,
            I => \N__5207\
        );

    \I__1036\ : Sp12to4
    port map (
            O => \N__5227\,
            I => \N__5207\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5224\,
            I => \N__5207\
        );

    \I__1034\ : Span4Mux_v
    port map (
            O => \N__5219\,
            I => \N__5202\
        );

    \I__1033\ : Span4Mux_v
    port map (
            O => \N__5214\,
            I => \N__5202\
        );

    \I__1032\ : Span12Mux_v
    port map (
            O => \N__5207\,
            I => \N__5199\
        );

    \I__1031\ : Sp12to4
    port map (
            O => \N__5202\,
            I => \N__5196\
        );

    \I__1030\ : Span12Mux_h
    port map (
            O => \N__5199\,
            I => \N__5193\
        );

    \I__1029\ : Span12Mux_h
    port map (
            O => \N__5196\,
            I => \N__5190\
        );

    \I__1028\ : Odrv12
    port map (
            O => \N__5193\,
            I => \RESETn_c\
        );

    \I__1027\ : Odrv12
    port map (
            O => \N__5190\,
            I => \RESETn_c\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5180\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5175\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5175\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5180\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__5175\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5164\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5169\,
            I => \N__5164\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5164\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1018\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5158\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5158\,
            I => \U409_TRANSFER_ACK.N_3_0\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__5155\,
            I => \U409_TRANSFER_ACK.N_3_0_cascade_\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__5152\,
            I => \N__5147\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5144\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5141\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5138\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5144\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__5141\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5138\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__5131\,
            I => \U409_TRANSFER_ACK.N_6_0_cascade_\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__5128\,
            I => \N__5125\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5125\,
            I => \N__5120\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__5124\,
            I => \N__5116\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5123\,
            I => \N__5112\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5120\,
            I => \N__5109\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5119\,
            I => \N__5102\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5116\,
            I => \N__5102\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5102\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5112\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__998\ : Odrv4
    port map (
            O => \N__5109\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5102\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__996\ : InMux
    port map (
            O => \N__5095\,
            I => \N__5089\
        );

    \I__995\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5086\
        );

    \I__994\ : InMux
    port map (
            O => \N__5093\,
            I => \N__5081\
        );

    \I__993\ : InMux
    port map (
            O => \N__5092\,
            I => \N__5081\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5089\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5086\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5081\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__989\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5069\
        );

    \I__988\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5066\
        );

    \I__987\ : InMux
    port map (
            O => \N__5072\,
            I => \N__5063\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5069\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5066\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5063\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__983\ : InMux
    port map (
            O => \N__5056\,
            I => \N__5050\
        );

    \I__982\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5050\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5050\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__980\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5041\
        );

    \I__979\ : InMux
    port map (
            O => \N__5046\,
            I => \N__5038\
        );

    \I__978\ : InMux
    port map (
            O => \N__5045\,
            I => \N__5035\
        );

    \I__977\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5032\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5041\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__5038\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5035\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__5032\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__5023\,
            I => \N__5016\
        );

    \I__971\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5013\
        );

    \I__970\ : InMux
    port map (
            O => \N__5021\,
            I => \N__5010\
        );

    \I__969\ : InMux
    port map (
            O => \N__5020\,
            I => \N__5007\
        );

    \I__968\ : InMux
    port map (
            O => \N__5019\,
            I => \N__5002\
        );

    \I__967\ : InMux
    port map (
            O => \N__5016\,
            I => \N__5002\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5013\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__5010\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5007\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__5002\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__4993\,
            I => \N__4987\
        );

    \I__961\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4980\
        );

    \I__960\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4980\
        );

    \I__959\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4977\
        );

    \I__958\ : InMux
    port map (
            O => \N__4987\,
            I => \N__4974\
        );

    \I__957\ : InMux
    port map (
            O => \N__4986\,
            I => \N__4971\
        );

    \I__956\ : InMux
    port map (
            O => \N__4985\,
            I => \N__4968\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4980\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4977\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4974\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4971\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4968\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__4957\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_\
        );

    \I__949\ : CascadeMux
    port map (
            O => \N__4954\,
            I => \N__4951\
        );

    \I__948\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4945\
        );

    \I__947\ : InMux
    port map (
            O => \N__4950\,
            I => \N__4945\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4945\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__945\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4939\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4939\,
            I => \N__4935\
        );

    \I__943\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4932\
        );

    \I__942\ : Span4Mux_v
    port map (
            O => \N__4935\,
            I => \N__4925\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__4932\,
            I => \N__4925\
        );

    \I__940\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4922\
        );

    \I__939\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4919\
        );

    \I__938\ : Span4Mux_h
    port map (
            O => \N__4925\,
            I => \N__4913\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4922\,
            I => \N__4913\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4919\,
            I => \N__4910\
        );

    \I__935\ : CascadeMux
    port map (
            O => \N__4918\,
            I => \N__4907\
        );

    \I__934\ : Span4Mux_v
    port map (
            O => \N__4913\,
            I => \N__4904\
        );

    \I__933\ : Span4Mux_v
    port map (
            O => \N__4910\,
            I => \N__4901\
        );

    \I__932\ : InMux
    port map (
            O => \N__4907\,
            I => \N__4898\
        );

    \I__931\ : Sp12to4
    port map (
            O => \N__4904\,
            I => \N__4891\
        );

    \I__930\ : Sp12to4
    port map (
            O => \N__4901\,
            I => \N__4891\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4898\,
            I => \N__4891\
        );

    \I__928\ : Span12Mux_h
    port map (
            O => \N__4891\,
            I => \N__4888\
        );

    \I__927\ : Span12Mux_v
    port map (
            O => \N__4888\,
            I => \N__4885\
        );

    \I__926\ : Odrv12
    port map (
            O => \N__4885\,
            I => \TSn_c\
        );

    \I__925\ : IoInMux
    port map (
            O => \N__4882\,
            I => \N__4879\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4879\,
            I => \N__4875\
        );

    \I__923\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4872\
        );

    \I__922\ : IoSpan4Mux
    port map (
            O => \N__4875\,
            I => \N__4868\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4872\,
            I => \N__4865\
        );

    \I__920\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4862\
        );

    \I__919\ : Span4Mux_s0_v
    port map (
            O => \N__4868\,
            I => \N__4856\
        );

    \I__918\ : Span4Mux_v
    port map (
            O => \N__4865\,
            I => \N__4853\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4862\,
            I => \N__4850\
        );

    \I__916\ : InMux
    port map (
            O => \N__4861\,
            I => \N__4847\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__4860\,
            I => \N__4844\
        );

    \I__914\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4841\
        );

    \I__913\ : Sp12to4
    port map (
            O => \N__4856\,
            I => \N__4837\
        );

    \I__912\ : Sp12to4
    port map (
            O => \N__4853\,
            I => \N__4834\
        );

    \I__911\ : Span4Mux_h
    port map (
            O => \N__4850\,
            I => \N__4829\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4847\,
            I => \N__4829\
        );

    \I__909\ : InMux
    port map (
            O => \N__4844\,
            I => \N__4826\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4841\,
            I => \N__4823\
        );

    \I__907\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4820\
        );

    \I__906\ : Span12Mux_v
    port map (
            O => \N__4837\,
            I => \N__4811\
        );

    \I__905\ : Span12Mux_h
    port map (
            O => \N__4834\,
            I => \N__4811\
        );

    \I__904\ : Sp12to4
    port map (
            O => \N__4829\,
            I => \N__4811\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4826\,
            I => \N__4811\
        );

    \I__902\ : Span12Mux_h
    port map (
            O => \N__4823\,
            I => \N__4808\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4820\,
            I => \N__4805\
        );

    \I__900\ : Span12Mux_v
    port map (
            O => \N__4811\,
            I => \N__4802\
        );

    \I__899\ : Span12Mux_v
    port map (
            O => \N__4808\,
            I => \N__4799\
        );

    \I__898\ : Span12Mux_v
    port map (
            O => \N__4805\,
            I => \N__4796\
        );

    \I__897\ : Odrv12
    port map (
            O => \N__4802\,
            I => \CLK40_IN_c\
        );

    \I__896\ : Odrv12
    port map (
            O => \N__4799\,
            I => \CLK40_IN_c\
        );

    \I__895\ : Odrv12
    port map (
            O => \N__4796\,
            I => \CLK40_IN_c\
        );

    \I__894\ : InMux
    port map (
            O => \N__4789\,
            I => \N__4785\
        );

    \I__893\ : InMux
    port map (
            O => \N__4788\,
            I => \N__4782\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4785\,
            I => \U409_TRANSFER_ACK.N_70\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__4782\,
            I => \U409_TRANSFER_ACK.N_70\
        );

    \I__890\ : InMux
    port map (
            O => \N__4777\,
            I => \N__4771\
        );

    \I__889\ : InMux
    port map (
            O => \N__4776\,
            I => \N__4771\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4771\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__4768\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\
        );

    \I__886\ : InMux
    port map (
            O => \N__4765\,
            I => \N__4762\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4762\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out\
        );

    \I__884\ : IoInMux
    port map (
            O => \N__4759\,
            I => \N__4756\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4756\,
            I => \N__4753\
        );

    \I__882\ : Span4Mux_s3_v
    port map (
            O => \N__4753\,
            I => \N__4750\
        );

    \I__881\ : Span4Mux_h
    port map (
            O => \N__4750\,
            I => \N__4747\
        );

    \I__880\ : Odrv4
    port map (
            O => \N__4747\,
            I => \CONSTANT_ONE_NET\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__4744\,
            I => \N__4741\
        );

    \I__878\ : InMux
    port map (
            O => \N__4741\,
            I => \N__4737\
        );

    \I__877\ : InMux
    port map (
            O => \N__4740\,
            I => \N__4734\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4737\,
            I => \N__4731\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4734\,
            I => \U409_TRANSFER_ACK.CO1\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__4731\,
            I => \U409_TRANSFER_ACK.CO1\
        );

    \I__873\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4723\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4723\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__4720\,
            I => \N__4714\
        );

    \I__870\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4711\
        );

    \I__869\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4708\
        );

    \I__868\ : InMux
    port map (
            O => \N__4717\,
            I => \N__4703\
        );

    \I__867\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4703\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4711\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4708\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4703\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__4696\,
            I => \N__4690\
        );

    \I__862\ : InMux
    port map (
            O => \N__4695\,
            I => \N__4686\
        );

    \I__861\ : InMux
    port map (
            O => \N__4694\,
            I => \N__4683\
        );

    \I__860\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4680\
        );

    \I__859\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4675\
        );

    \I__858\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4675\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4686\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4683\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4680\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4675\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__853\ : CascadeMux
    port map (
            O => \N__4666\,
            I => \N__4663\
        );

    \I__852\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4660\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4660\,
            I => \U409_TRANSFER_ACK.ROM_TACK_EN_e_1\
        );

    \I__850\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4654\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4654\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\
        );

    \I__848\ : InMux
    port map (
            O => \N__4651\,
            I => \N__4647\
        );

    \I__847\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4644\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4647\,
            I => \U409_TRANSFER_ACK.N_17_mux\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4644\,
            I => \U409_TRANSFER_ACK.N_17_mux\
        );

    \I__844\ : InMux
    port map (
            O => \N__4639\,
            I => \N__4635\
        );

    \I__843\ : InMux
    port map (
            O => \N__4638\,
            I => \N__4632\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4635\,
            I => \N__4629\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4632\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__4629\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__839\ : CascadeMux
    port map (
            O => \N__4624\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3_cascade_\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__4621\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_3_cascade_\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__4618\,
            I => \U409_TRANSFER_ACK.N_70_cascade_\
        );

    \I__836\ : InMux
    port map (
            O => \N__4615\,
            I => \N__4611\
        );

    \I__835\ : InMux
    port map (
            O => \N__4614\,
            I => \N__4608\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4611\,
            I => \U409_TRANSFER_ACK.N_55\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4608\,
            I => \U409_TRANSFER_ACK.N_55\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__4603\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__4600\,
            I => \N__4596\
        );

    \I__830\ : InMux
    port map (
            O => \N__4599\,
            I => \N__4589\
        );

    \I__829\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4589\
        );

    \I__828\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4584\
        );

    \I__827\ : InMux
    port map (
            O => \N__4594\,
            I => \N__4584\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4589\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4584\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__824\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4570\
        );

    \I__823\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4570\
        );

    \I__822\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4570\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4570\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__4567\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_\
        );

    \I__819\ : InMux
    port map (
            O => \N__4564\,
            I => \N__4560\
        );

    \I__818\ : InMux
    port map (
            O => \N__4563\,
            I => \N__4557\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4560\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4557\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__815\ : InMux
    port map (
            O => \N__4552\,
            I => \N__4548\
        );

    \I__814\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4545\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4548\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__4545\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__4540\,
            I => \N__4536\
        );

    \I__810\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4533\
        );

    \I__809\ : InMux
    port map (
            O => \N__4536\,
            I => \N__4530\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4533\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4530\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__4525\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__4522\,
            I => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\
        );

    \I__804\ : IoInMux
    port map (
            O => \N__4519\,
            I => \N__4516\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4516\,
            I => \N__4513\
        );

    \I__802\ : Span12Mux_s7_v
    port map (
            O => \N__4513\,
            I => \N__4510\
        );

    \I__801\ : Span12Mux_v
    port map (
            O => \N__4510\,
            I => \N__4507\
        );

    \I__800\ : Span12Mux_h
    port map (
            O => \N__4507\,
            I => \N__4502\
        );

    \I__799\ : InMux
    port map (
            O => \N__4506\,
            I => \N__4497\
        );

    \I__798\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4497\
        );

    \I__797\ : Odrv12
    port map (
            O => \N__4502\,
            I => \TACK_OUTn\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4497\,
            I => \TACK_OUTn\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__4492\,
            I => \N__4487\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__4491\,
            I => \N__4483\
        );

    \I__793\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4479\
        );

    \I__792\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4472\
        );

    \I__791\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4472\
        );

    \I__790\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4472\
        );

    \I__789\ : InMux
    port map (
            O => \N__4482\,
            I => \N__4469\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4479\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4472\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4469\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__785\ : InMux
    port map (
            O => \N__4462\,
            I => \N__4455\
        );

    \I__784\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4446\
        );

    \I__783\ : InMux
    port map (
            O => \N__4460\,
            I => \N__4446\
        );

    \I__782\ : InMux
    port map (
            O => \N__4459\,
            I => \N__4446\
        );

    \I__781\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4446\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4455\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4446\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__778\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4436\
        );

    \I__777\ : InMux
    port map (
            O => \N__4440\,
            I => \N__4431\
        );

    \I__776\ : InMux
    port map (
            O => \N__4439\,
            I => \N__4431\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4436\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4431\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__773\ : CEMux
    port map (
            O => \N__4426\,
            I => \N__4423\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__4423\,
            I => \N__4420\
        );

    \I__771\ : Span4Mux_v
    port map (
            O => \N__4420\,
            I => \N__4417\
        );

    \I__770\ : Span4Mux_h
    port map (
            O => \N__4417\,
            I => \N__4414\
        );

    \I__769\ : Odrv4
    port map (
            O => \N__4414\,
            I => \U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__4411\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_cascade_\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__4408\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_cascade_\
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__4405\,
            I => \N__4402\
        );

    \I__765\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4395\
        );

    \I__764\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4395\
        );

    \I__763\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4392\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4395\,
            I => \N__4389\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4392\,
            I => \N__4386\
        );

    \I__760\ : Span4Mux_h
    port map (
            O => \N__4389\,
            I => \N__4383\
        );

    \I__759\ : Span4Mux_v
    port map (
            O => \N__4386\,
            I => \N__4380\
        );

    \I__758\ : Span4Mux_v
    port map (
            O => \N__4383\,
            I => \N__4377\
        );

    \I__757\ : Odrv4
    port map (
            O => \N__4380\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__4377\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\
        );

    \I__755\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4368\
        );

    \I__754\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4365\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4368\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__4365\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\
        );

    \I__751\ : InMux
    port map (
            O => \N__4360\,
            I => \N__4356\
        );

    \I__750\ : InMux
    port map (
            O => \N__4359\,
            I => \N__4353\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4356\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4353\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\
        );

    \I__747\ : IoInMux
    port map (
            O => \N__4348\,
            I => \N__4345\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4345\,
            I => \N__4342\
        );

    \I__745\ : IoSpan4Mux
    port map (
            O => \N__4342\,
            I => \N__4339\
        );

    \I__744\ : IoSpan4Mux
    port map (
            O => \N__4339\,
            I => \N__4336\
        );

    \I__743\ : Span4Mux_s0_v
    port map (
            O => \N__4336\,
            I => \N__4333\
        );

    \I__742\ : Sp12to4
    port map (
            O => \N__4333\,
            I => \N__4329\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__4332\,
            I => \N__4326\
        );

    \I__740\ : Span12Mux_s11_v
    port map (
            O => \N__4329\,
            I => \N__4323\
        );

    \I__739\ : InMux
    port map (
            O => \N__4326\,
            I => \N__4320\
        );

    \I__738\ : Odrv12
    port map (
            O => \N__4323\,
            I => \ROMENn_c\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__4320\,
            I => \ROMENn_c\
        );

    \I__736\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4308\
        );

    \I__735\ : InMux
    port map (
            O => \N__4314\,
            I => \N__4305\
        );

    \I__734\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4298\
        );

    \I__733\ : InMux
    port map (
            O => \N__4312\,
            I => \N__4298\
        );

    \I__732\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4298\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4308\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4305\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__4298\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__728\ : InMux
    port map (
            O => \N__4291\,
            I => \N__4283\
        );

    \I__727\ : InMux
    port map (
            O => \N__4290\,
            I => \N__4280\
        );

    \I__726\ : InMux
    port map (
            O => \N__4289\,
            I => \N__4271\
        );

    \I__725\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4271\
        );

    \I__724\ : InMux
    port map (
            O => \N__4287\,
            I => \N__4271\
        );

    \I__723\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4271\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4283\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4280\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4271\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__719\ : InMux
    port map (
            O => \N__4264\,
            I => \N__4261\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__4261\,
            I => \N__4258\
        );

    \I__717\ : Odrv12
    port map (
            O => \N__4258\,
            I => \U409_TRANSFER_ACK.N_71\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__4255\,
            I => \N__4252\
        );

    \I__715\ : InMux
    port map (
            O => \N__4252\,
            I => \N__4249\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__4249\,
            I => \N__4246\
        );

    \I__713\ : Span4Mux_v
    port map (
            O => \N__4246\,
            I => \N__4243\
        );

    \I__712\ : Span4Mux_h
    port map (
            O => \N__4243\,
            I => \N__4240\
        );

    \I__711\ : Sp12to4
    port map (
            O => \N__4240\,
            I => \N__4237\
        );

    \I__710\ : Span12Mux_h
    port map (
            O => \N__4237\,
            I => \N__4234\
        );

    \I__709\ : Span12Mux_v
    port map (
            O => \N__4234\,
            I => \N__4231\
        );

    \I__708\ : Odrv12
    port map (
            O => \N__4231\,
            I => \TACKn_in\
        );

    \I__707\ : IoInMux
    port map (
            O => \N__4228\,
            I => \N__4225\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4225\,
            I => \N__4222\
        );

    \I__705\ : Span4Mux_s2_v
    port map (
            O => \N__4222\,
            I => \N__4219\
        );

    \I__704\ : Span4Mux_h
    port map (
            O => \N__4219\,
            I => \N__4216\
        );

    \I__703\ : Sp12to4
    port map (
            O => \N__4216\,
            I => \N__4213\
        );

    \I__702\ : Span12Mux_v
    port map (
            O => \N__4213\,
            I => \N__4210\
        );

    \I__701\ : Odrv12
    port map (
            O => \N__4210\,
            I => \N_67_i\
        );

    \I__700\ : InMux
    port map (
            O => \N__4207\,
            I => \N__4204\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__4204\,
            I => \N__4201\
        );

    \I__698\ : Span4Mux_v
    port map (
            O => \N__4201\,
            I => \N__4196\
        );

    \I__697\ : InMux
    port map (
            O => \N__4200\,
            I => \N__4193\
        );

    \I__696\ : InMux
    port map (
            O => \N__4199\,
            I => \N__4190\
        );

    \I__695\ : Span4Mux_h
    port map (
            O => \N__4196\,
            I => \N__4183\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4193\,
            I => \N__4183\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4190\,
            I => \N__4183\
        );

    \I__692\ : Odrv4
    port map (
            O => \N__4183\,
            I => \N_100\
        );

    \I__691\ : InMux
    port map (
            O => \N__4180\,
            I => \N__4177\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4177\,
            I => \N__4174\
        );

    \I__689\ : Span4Mux_h
    port map (
            O => \N__4174\,
            I => \N__4169\
        );

    \I__688\ : InMux
    port map (
            O => \N__4173\,
            I => \N__4164\
        );

    \I__687\ : InMux
    port map (
            O => \N__4172\,
            I => \N__4164\
        );

    \I__686\ : Span4Mux_v
    port map (
            O => \N__4169\,
            I => \N__4161\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4164\,
            I => \N__4158\
        );

    \I__684\ : Sp12to4
    port map (
            O => \N__4161\,
            I => \N__4153\
        );

    \I__683\ : Span12Mux_v
    port map (
            O => \N__4158\,
            I => \N__4153\
        );

    \I__682\ : Span12Mux_v
    port map (
            O => \N__4153\,
            I => \N__4150\
        );

    \I__681\ : Span12Mux_h
    port map (
            O => \N__4150\,
            I => \N__4147\
        );

    \I__680\ : Odrv12
    port map (
            O => \N__4147\,
            I => \OVL_c\
        );

    \I__679\ : InMux
    port map (
            O => \N__4144\,
            I => \N__4141\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__4141\,
            I => \N__4138\
        );

    \I__677\ : Span4Mux_v
    port map (
            O => \N__4138\,
            I => \N__4134\
        );

    \I__676\ : InMux
    port map (
            O => \N__4137\,
            I => \N__4131\
        );

    \I__675\ : Odrv4
    port map (
            O => \N__4134\,
            I => \N_67\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__4131\,
            I => \N_67\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__4126\,
            I => \N__4123\
        );

    \I__672\ : InMux
    port map (
            O => \N__4123\,
            I => \N__4119\
        );

    \I__671\ : CascadeMux
    port map (
            O => \N__4122\,
            I => \N__4116\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4119\,
            I => \N__4113\
        );

    \I__669\ : InMux
    port map (
            O => \N__4116\,
            I => \N__4110\
        );

    \I__668\ : Span4Mux_h
    port map (
            O => \N__4113\,
            I => \N__4105\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4110\,
            I => \N__4105\
        );

    \I__666\ : Span4Mux_v
    port map (
            O => \N__4105\,
            I => \N__4102\
        );

    \I__665\ : Span4Mux_h
    port map (
            O => \N__4102\,
            I => \N__4099\
        );

    \I__664\ : Odrv4
    port map (
            O => \N__4099\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\
        );

    \I__663\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4092\
        );

    \I__662\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4089\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4092\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4089\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__659\ : InMux
    port map (
            O => \N__4084\,
            I => \N__4081\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4081\,
            I => \N__4078\
        );

    \I__657\ : Odrv4
    port map (
            O => \N__4078\,
            I => \U409_TRANSFER_ACK.N_106\
        );

    \I__656\ : InMux
    port map (
            O => \N__4075\,
            I => \N__4072\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__4072\,
            I => \N__4069\
        );

    \I__654\ : Span4Mux_h
    port map (
            O => \N__4069\,
            I => \N__4066\
        );

    \I__653\ : Odrv4
    port map (
            O => \N__4066\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER15Z0Z_1\
        );

    \I__652\ : InMux
    port map (
            O => \N__4063\,
            I => \N__4058\
        );

    \I__651\ : InMux
    port map (
            O => \N__4062\,
            I => \N__4052\
        );

    \I__650\ : InMux
    port map (
            O => \N__4061\,
            I => \N__4052\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4058\,
            I => \N__4049\
        );

    \I__648\ : InMux
    port map (
            O => \N__4057\,
            I => \N__4046\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4052\,
            I => \N__4043\
        );

    \I__646\ : Span4Mux_h
    port map (
            O => \N__4049\,
            I => \N__4038\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4046\,
            I => \N__4038\
        );

    \I__644\ : Odrv12
    port map (
            O => \N__4043\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__643\ : Odrv4
    port map (
            O => \N__4038\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__642\ : InMux
    port map (
            O => \N__4033\,
            I => \N__4030\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__4030\,
            I => \N__4027\
        );

    \I__640\ : Odrv12
    port map (
            O => \N__4027\,
            I => \U409_DATA_BUFFERS.un1_BUFENn_iZ0Z_0\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__4024\,
            I => \N__4021\
        );

    \I__638\ : InMux
    port map (
            O => \N__4021\,
            I => \N__4018\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4018\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1\
        );

    \I__636\ : InMux
    port map (
            O => \N__4015\,
            I => \N__4011\
        );

    \I__635\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4008\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4011\,
            I => \N__4004\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4008\,
            I => \N__4001\
        );

    \I__632\ : InMux
    port map (
            O => \N__4007\,
            I => \N__3996\
        );

    \I__631\ : Span4Mux_v
    port map (
            O => \N__4004\,
            I => \N__3991\
        );

    \I__630\ : Span4Mux_v
    port map (
            O => \N__4001\,
            I => \N__3991\
        );

    \I__629\ : InMux
    port map (
            O => \N__4000\,
            I => \N__3988\
        );

    \I__628\ : InMux
    port map (
            O => \N__3999\,
            I => \N__3985\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3996\,
            I => \N__3982\
        );

    \I__626\ : Sp12to4
    port map (
            O => \N__3991\,
            I => \N__3977\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3988\,
            I => \N__3977\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3985\,
            I => \N__3974\
        );

    \I__623\ : Span12Mux_v
    port map (
            O => \N__3982\,
            I => \N__3971\
        );

    \I__622\ : Span12Mux_h
    port map (
            O => \N__3977\,
            I => \N__3966\
        );

    \I__621\ : Span12Mux_v
    port map (
            O => \N__3974\,
            I => \N__3966\
        );

    \I__620\ : Odrv12
    port map (
            O => \N__3971\,
            I => \A_c_20\
        );

    \I__619\ : Odrv12
    port map (
            O => \N__3966\,
            I => \A_c_20\
        );

    \I__618\ : CascadeMux
    port map (
            O => \N__3961\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__3958\,
            I => \CIA_SPACE_cascade_\
        );

    \I__616\ : InMux
    port map (
            O => \N__3955\,
            I => \N__3952\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3952\,
            I => \U409_ADDRESS_DECODE.N_69\
        );

    \I__614\ : IoInMux
    port map (
            O => \N__3949\,
            I => \N__3946\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3946\,
            I => \N__3943\
        );

    \I__612\ : IoSpan4Mux
    port map (
            O => \N__3943\,
            I => \N__3940\
        );

    \I__611\ : Span4Mux_s2_v
    port map (
            O => \N__3940\,
            I => \N__3937\
        );

    \I__610\ : Span4Mux_v
    port map (
            O => \N__3937\,
            I => \N__3934\
        );

    \I__609\ : Span4Mux_v
    port map (
            O => \N__3934\,
            I => \N__3931\
        );

    \I__608\ : Odrv4
    port map (
            O => \N__3931\,
            I => \PORTSIZE_0_i\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__3928\,
            I => \U409_ADDRESS_DECODE.un5_RAMSPACEn_cascade_\
        );

    \I__606\ : InMux
    port map (
            O => \N__3925\,
            I => \N__3914\
        );

    \I__605\ : InMux
    port map (
            O => \N__3924\,
            I => \N__3914\
        );

    \I__604\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3914\
        );

    \I__603\ : InMux
    port map (
            O => \N__3922\,
            I => \N__3909\
        );

    \I__602\ : InMux
    port map (
            O => \N__3921\,
            I => \N__3909\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3914\,
            I => \N__3906\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3909\,
            I => \N__3903\
        );

    \I__599\ : Span4Mux_v
    port map (
            O => \N__3906\,
            I => \N__3899\
        );

    \I__598\ : Span4Mux_v
    port map (
            O => \N__3903\,
            I => \N__3896\
        );

    \I__597\ : InMux
    port map (
            O => \N__3902\,
            I => \N__3893\
        );

    \I__596\ : Sp12to4
    port map (
            O => \N__3899\,
            I => \N__3886\
        );

    \I__595\ : Sp12to4
    port map (
            O => \N__3896\,
            I => \N__3886\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3893\,
            I => \N__3886\
        );

    \I__593\ : Odrv12
    port map (
            O => \N__3886\,
            I => \A_c_21\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__3883\,
            I => \N__3879\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__3882\,
            I => \N__3876\
        );

    \I__590\ : InMux
    port map (
            O => \N__3879\,
            I => \N__3871\
        );

    \I__589\ : InMux
    port map (
            O => \N__3876\,
            I => \N__3871\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3871\,
            I => \N__3865\
        );

    \I__587\ : InMux
    port map (
            O => \N__3870\,
            I => \N__3862\
        );

    \I__586\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3857\
        );

    \I__585\ : InMux
    port map (
            O => \N__3868\,
            I => \N__3857\
        );

    \I__584\ : Span4Mux_v
    port map (
            O => \N__3865\,
            I => \N__3854\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3862\,
            I => \N__3849\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__3857\,
            I => \N__3849\
        );

    \I__581\ : Span4Mux_h
    port map (
            O => \N__3854\,
            I => \N__3846\
        );

    \I__580\ : Span4Mux_v
    port map (
            O => \N__3849\,
            I => \N__3843\
        );

    \I__579\ : Sp12to4
    port map (
            O => \N__3846\,
            I => \N__3838\
        );

    \I__578\ : Sp12to4
    port map (
            O => \N__3843\,
            I => \N__3838\
        );

    \I__577\ : Odrv12
    port map (
            O => \N__3838\,
            I => \A_c_23\
        );

    \I__576\ : InMux
    port map (
            O => \N__3835\,
            I => \N__3824\
        );

    \I__575\ : InMux
    port map (
            O => \N__3834\,
            I => \N__3824\
        );

    \I__574\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3824\
        );

    \I__573\ : InMux
    port map (
            O => \N__3832\,
            I => \N__3819\
        );

    \I__572\ : InMux
    port map (
            O => \N__3831\,
            I => \N__3819\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3824\,
            I => \N__3814\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3819\,
            I => \N__3814\
        );

    \I__569\ : Sp12to4
    port map (
            O => \N__3814\,
            I => \N__3811\
        );

    \I__568\ : Span12Mux_v
    port map (
            O => \N__3811\,
            I => \N__3808\
        );

    \I__567\ : Odrv12
    port map (
            O => \N__3808\,
            I => \A_c_22\
        );

    \I__566\ : CascadeMux
    port map (
            O => \N__3805\,
            I => \N__3799\
        );

    \I__565\ : InMux
    port map (
            O => \N__3804\,
            I => \N__3792\
        );

    \I__564\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3792\
        );

    \I__563\ : InMux
    port map (
            O => \N__3802\,
            I => \N__3792\
        );

    \I__562\ : InMux
    port map (
            O => \N__3799\,
            I => \N__3789\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3792\,
            I => \N__3784\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3789\,
            I => \N__3784\
        );

    \I__559\ : Span12Mux_h
    port map (
            O => \N__3784\,
            I => \N__3781\
        );

    \I__558\ : Span12Mux_v
    port map (
            O => \N__3781\,
            I => \N__3778\
        );

    \I__557\ : Odrv12
    port map (
            O => \N__3778\,
            I => \TM_c_0\
        );

    \I__556\ : InMux
    port map (
            O => \N__3775\,
            I => \N__3772\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3772\,
            I => \U409_ADDRESS_DECODE_HIROM\
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__3769\,
            I => \U409_ADDRESS_DECODE_LOWROM_cascade_\
        );

    \I__553\ : InMux
    port map (
            O => \N__3766\,
            I => \N__3756\
        );

    \I__552\ : InMux
    port map (
            O => \N__3765\,
            I => \N__3756\
        );

    \I__551\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3756\
        );

    \I__550\ : InMux
    port map (
            O => \N__3763\,
            I => \N__3753\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3756\,
            I => \N__3748\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3753\,
            I => \N__3748\
        );

    \I__547\ : Span4Mux_h
    port map (
            O => \N__3748\,
            I => \N__3745\
        );

    \I__546\ : Sp12to4
    port map (
            O => \N__3745\,
            I => \N__3742\
        );

    \I__545\ : Odrv12
    port map (
            O => \N__3742\,
            I => \TM_c_1\
        );

    \I__544\ : InMux
    port map (
            O => \N__3739\,
            I => \N__3735\
        );

    \I__543\ : InMux
    port map (
            O => \N__3738\,
            I => \N__3731\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3735\,
            I => \N__3725\
        );

    \I__541\ : InMux
    port map (
            O => \N__3734\,
            I => \N__3722\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__3731\,
            I => \N__3719\
        );

    \I__539\ : InMux
    port map (
            O => \N__3730\,
            I => \N__3716\
        );

    \I__538\ : InMux
    port map (
            O => \N__3729\,
            I => \N__3713\
        );

    \I__537\ : InMux
    port map (
            O => \N__3728\,
            I => \N__3710\
        );

    \I__536\ : Odrv12
    port map (
            O => \N__3725\,
            I => \N_107\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3722\,
            I => \N_107\
        );

    \I__534\ : Odrv4
    port map (
            O => \N__3719\,
            I => \N_107\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3716\,
            I => \N_107\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3713\,
            I => \N_107\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3710\,
            I => \N_107\
        );

    \I__530\ : InMux
    port map (
            O => \N__3697\,
            I => \N__3693\
        );

    \I__529\ : InMux
    port map (
            O => \N__3696\,
            I => \N__3689\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3693\,
            I => \N__3686\
        );

    \I__527\ : InMux
    port map (
            O => \N__3692\,
            I => \N__3683\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3689\,
            I => \N__3680\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__3686\,
            I => \N_33\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3683\,
            I => \N_33\
        );

    \I__523\ : Odrv4
    port map (
            O => \N__3680\,
            I => \N_33\
        );

    \I__522\ : IoInMux
    port map (
            O => \N__3673\,
            I => \N__3670\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3670\,
            I => \N__3667\
        );

    \I__520\ : IoSpan4Mux
    port map (
            O => \N__3667\,
            I => \N__3664\
        );

    \I__519\ : IoSpan4Mux
    port map (
            O => \N__3664\,
            I => \N__3661\
        );

    \I__518\ : Sp12to4
    port map (
            O => \N__3661\,
            I => \N__3658\
        );

    \I__517\ : Span12Mux_v
    port map (
            O => \N__3658\,
            I => \N__3655\
        );

    \I__516\ : Odrv12
    port map (
            O => \N__3655\,
            I => \N_68_i\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__3652\,
            I => \N_74_1_cascade_\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__3649\,
            I => \N_33_cascade_\
        );

    \I__513\ : InMux
    port map (
            O => \N__3646\,
            I => \N__3643\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3643\,
            I => \N_99\
        );

    \I__511\ : InMux
    port map (
            O => \N__3640\,
            I => \N__3636\
        );

    \I__510\ : InMux
    port map (
            O => \N__3639\,
            I => \N__3633\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3636\,
            I => \N__3628\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3633\,
            I => \N__3628\
        );

    \I__507\ : Span4Mux_v
    port map (
            O => \N__3628\,
            I => \N__3624\
        );

    \I__506\ : InMux
    port map (
            O => \N__3627\,
            I => \N__3621\
        );

    \I__505\ : Odrv4
    port map (
            O => \N__3624\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_5\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3621\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_5\
        );

    \I__503\ : CascadeMux
    port map (
            O => \N__3616\,
            I => \N_99_cascade_\
        );

    \I__502\ : InMux
    port map (
            O => \N__3613\,
            I => \N__3610\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3610\,
            I => \N__3605\
        );

    \I__500\ : InMux
    port map (
            O => \N__3609\,
            I => \N__3602\
        );

    \I__499\ : InMux
    port map (
            O => \N__3608\,
            I => \N__3599\
        );

    \I__498\ : Span4Mux_v
    port map (
            O => \N__3605\,
            I => \N__3594\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3602\,
            I => \N__3594\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3599\,
            I => \N__3591\
        );

    \I__495\ : Span4Mux_h
    port map (
            O => \N__3594\,
            I => \N__3588\
        );

    \I__494\ : Span4Mux_v
    port map (
            O => \N__3591\,
            I => \N__3585\
        );

    \I__493\ : Odrv4
    port map (
            O => \N__3588\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_4\
        );

    \I__492\ : Odrv4
    port map (
            O => \N__3585\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_4\
        );

    \I__491\ : InMux
    port map (
            O => \N__3580\,
            I => \N__3574\
        );

    \I__490\ : InMux
    port map (
            O => \N__3579\,
            I => \N__3571\
        );

    \I__489\ : InMux
    port map (
            O => \N__3578\,
            I => \N__3568\
        );

    \I__488\ : InMux
    port map (
            O => \N__3577\,
            I => \N__3565\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3574\,
            I => \N__3558\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3571\,
            I => \N__3558\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3568\,
            I => \N__3558\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3565\,
            I => \N__3555\
        );

    \I__483\ : Span4Mux_v
    port map (
            O => \N__3558\,
            I => \N__3552\
        );

    \I__482\ : Span4Mux_v
    port map (
            O => \N__3555\,
            I => \N__3549\
        );

    \I__481\ : Sp12to4
    port map (
            O => \N__3552\,
            I => \N__3544\
        );

    \I__480\ : Sp12to4
    port map (
            O => \N__3549\,
            I => \N__3544\
        );

    \I__479\ : Span12Mux_h
    port map (
            O => \N__3544\,
            I => \N__3541\
        );

    \I__478\ : Span12Mux_v
    port map (
            O => \N__3541\,
            I => \N__3538\
        );

    \I__477\ : Odrv12
    port map (
            O => \N__3538\,
            I => \A_c_18\
        );

    \I__476\ : InMux
    port map (
            O => \N__3535\,
            I => \N__3532\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__3532\,
            I => \N__3528\
        );

    \I__474\ : CascadeMux
    port map (
            O => \N__3531\,
            I => \N__3525\
        );

    \I__473\ : Span4Mux_v
    port map (
            O => \N__3528\,
            I => \N__3522\
        );

    \I__472\ : InMux
    port map (
            O => \N__3525\,
            I => \N__3519\
        );

    \I__471\ : Odrv4
    port map (
            O => \N__3522\,
            I => \N_74_1\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3519\,
            I => \N_74_1\
        );

    \I__469\ : InMux
    port map (
            O => \N__3514\,
            I => \N__3509\
        );

    \I__468\ : InMux
    port map (
            O => \N__3513\,
            I => \N__3506\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__3512\,
            I => \N__3503\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3509\,
            I => \N__3500\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3506\,
            I => \N__3497\
        );

    \I__464\ : InMux
    port map (
            O => \N__3503\,
            I => \N__3494\
        );

    \I__463\ : Odrv4
    port map (
            O => \N__3500\,
            I => \N_101\
        );

    \I__462\ : Odrv4
    port map (
            O => \N__3497\,
            I => \N_101\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3494\,
            I => \N_101\
        );

    \I__460\ : InMux
    port map (
            O => \N__3487\,
            I => \N__3484\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3484\,
            I => \N__3481\
        );

    \I__458\ : Span12Mux_h
    port map (
            O => \N__3481\,
            I => \N__3478\
        );

    \I__457\ : Span12Mux_v
    port map (
            O => \N__3478\,
            I => \N__3475\
        );

    \I__456\ : Odrv12
    port map (
            O => \N__3475\,
            I => \TT_c_0\
        );

    \I__455\ : InMux
    port map (
            O => \N__3472\,
            I => \N__3469\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3469\,
            I => \N__3466\
        );

    \I__453\ : Span4Mux_h
    port map (
            O => \N__3466\,
            I => \N__3463\
        );

    \I__452\ : Odrv4
    port map (
            O => \N__3463\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_9\
        );

    \I__451\ : InMux
    port map (
            O => \N__3460\,
            I => \N__3452\
        );

    \I__450\ : InMux
    port map (
            O => \N__3459\,
            I => \N__3452\
        );

    \I__449\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3449\
        );

    \I__448\ : InMux
    port map (
            O => \N__3457\,
            I => \N__3446\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3452\,
            I => \N__3440\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__3449\,
            I => \N__3440\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3446\,
            I => \N__3437\
        );

    \I__444\ : InMux
    port map (
            O => \N__3445\,
            I => \N__3434\
        );

    \I__443\ : Span4Mux_v
    port map (
            O => \N__3440\,
            I => \N__3431\
        );

    \I__442\ : Span4Mux_h
    port map (
            O => \N__3437\,
            I => \N__3428\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3434\,
            I => \N__3425\
        );

    \I__440\ : Sp12to4
    port map (
            O => \N__3431\,
            I => \N__3422\
        );

    \I__439\ : Span4Mux_h
    port map (
            O => \N__3428\,
            I => \N__3419\
        );

    \I__438\ : Span4Mux_h
    port map (
            O => \N__3425\,
            I => \N__3416\
        );

    \I__437\ : Span12Mux_h
    port map (
            O => \N__3422\,
            I => \N__3409\
        );

    \I__436\ : Sp12to4
    port map (
            O => \N__3419\,
            I => \N__3409\
        );

    \I__435\ : Sp12to4
    port map (
            O => \N__3416\,
            I => \N__3409\
        );

    \I__434\ : Span12Mux_v
    port map (
            O => \N__3409\,
            I => \N__3406\
        );

    \I__433\ : Odrv12
    port map (
            O => \N__3406\,
            I => \A_c_19\
        );

    \I__432\ : CascadeMux
    port map (
            O => \N__3403\,
            I => \U409_ADDRESS_DECODE.HIROMZ0Z_1_cascade_\
        );

    \I__431\ : InMux
    port map (
            O => \N__3400\,
            I => \N__3394\
        );

    \I__430\ : InMux
    port map (
            O => \N__3399\,
            I => \N__3394\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3394\,
            I => \U409_TRANSFER_ACK.N_94\
        );

    \I__428\ : InMux
    port map (
            O => \N__3391\,
            I => \N__3387\
        );

    \I__427\ : InMux
    port map (
            O => \N__3390\,
            I => \N__3383\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__3387\,
            I => \N__3380\
        );

    \I__425\ : InMux
    port map (
            O => \N__3386\,
            I => \N__3377\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3383\,
            I => \N__3374\
        );

    \I__423\ : Span4Mux_v
    port map (
            O => \N__3380\,
            I => \N__3371\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3377\,
            I => \N__3368\
        );

    \I__421\ : Span4Mux_v
    port map (
            O => \N__3374\,
            I => \N__3365\
        );

    \I__420\ : Sp12to4
    port map (
            O => \N__3371\,
            I => \N__3360\
        );

    \I__419\ : Span12Mux_v
    port map (
            O => \N__3368\,
            I => \N__3360\
        );

    \I__418\ : Span4Mux_h
    port map (
            O => \N__3365\,
            I => \N__3357\
        );

    \I__417\ : Odrv12
    port map (
            O => \N__3360\,
            I => \A_c_27\
        );

    \I__416\ : Odrv4
    port map (
            O => \N__3357\,
            I => \A_c_27\
        );

    \I__415\ : InMux
    port map (
            O => \N__3352\,
            I => \N__3346\
        );

    \I__414\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3346\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__3346\,
            I => \N__3342\
        );

    \I__412\ : InMux
    port map (
            O => \N__3345\,
            I => \N__3339\
        );

    \I__411\ : Span4Mux_h
    port map (
            O => \N__3342\,
            I => \N__3334\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3339\,
            I => \N__3334\
        );

    \I__409\ : Span4Mux_h
    port map (
            O => \N__3334\,
            I => \N__3331\
        );

    \I__408\ : Span4Mux_v
    port map (
            O => \N__3331\,
            I => \N__3328\
        );

    \I__407\ : Span4Mux_v
    port map (
            O => \N__3328\,
            I => \N__3325\
        );

    \I__406\ : Odrv4
    port map (
            O => \N__3325\,
            I => \A_c_26\
        );

    \I__405\ : CascadeMux
    port map (
            O => \N__3322\,
            I => \N__3317\
        );

    \I__404\ : CascadeMux
    port map (
            O => \N__3321\,
            I => \N__3314\
        );

    \I__403\ : InMux
    port map (
            O => \N__3320\,
            I => \N__3311\
        );

    \I__402\ : InMux
    port map (
            O => \N__3317\,
            I => \N__3306\
        );

    \I__401\ : InMux
    port map (
            O => \N__3314\,
            I => \N__3306\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3311\,
            I => \N__3303\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3306\,
            I => \N__3300\
        );

    \I__398\ : Span4Mux_v
    port map (
            O => \N__3303\,
            I => \N__3297\
        );

    \I__397\ : Sp12to4
    port map (
            O => \N__3300\,
            I => \N__3294\
        );

    \I__396\ : Span4Mux_v
    port map (
            O => \N__3297\,
            I => \N__3291\
        );

    \I__395\ : Span12Mux_v
    port map (
            O => \N__3294\,
            I => \N__3288\
        );

    \I__394\ : Span4Mux_h
    port map (
            O => \N__3291\,
            I => \N__3285\
        );

    \I__393\ : Odrv12
    port map (
            O => \N__3288\,
            I => \A_c_24\
        );

    \I__392\ : Odrv4
    port map (
            O => \N__3285\,
            I => \A_c_24\
        );

    \I__391\ : CascadeMux
    port map (
            O => \N__3280\,
            I => \N__3275\
        );

    \I__390\ : InMux
    port map (
            O => \N__3279\,
            I => \N__3270\
        );

    \I__389\ : InMux
    port map (
            O => \N__3278\,
            I => \N__3270\
        );

    \I__388\ : InMux
    port map (
            O => \N__3275\,
            I => \N__3267\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3270\,
            I => \N__3264\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__3267\,
            I => \N__3261\
        );

    \I__385\ : Span4Mux_v
    port map (
            O => \N__3264\,
            I => \N__3258\
        );

    \I__384\ : Span4Mux_v
    port map (
            O => \N__3261\,
            I => \N__3255\
        );

    \I__383\ : Sp12to4
    port map (
            O => \N__3258\,
            I => \N__3252\
        );

    \I__382\ : Span4Mux_h
    port map (
            O => \N__3255\,
            I => \N__3249\
        );

    \I__381\ : Odrv12
    port map (
            O => \N__3252\,
            I => \A_c_25\
        );

    \I__380\ : Odrv4
    port map (
            O => \N__3249\,
            I => \A_c_25\
        );

    \I__379\ : InMux
    port map (
            O => \N__3244\,
            I => \N__3241\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3241\,
            I => \N__3238\
        );

    \I__377\ : Odrv4
    port map (
            O => \N__3238\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_7\
        );

    \I__376\ : CascadeMux
    port map (
            O => \N__3235\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_8_cascade_\
        );

    \I__375\ : InMux
    port map (
            O => \N__3232\,
            I => \N__3229\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3229\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_10\
        );

    \I__373\ : IoInMux
    port map (
            O => \N__3226\,
            I => \N__3223\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3223\,
            I => \N__3220\
        );

    \I__371\ : IoSpan4Mux
    port map (
            O => \N__3220\,
            I => \N__3217\
        );

    \I__370\ : Span4Mux_s3_h
    port map (
            O => \N__3217\,
            I => \N__3214\
        );

    \I__369\ : Sp12to4
    port map (
            O => \N__3214\,
            I => \N__3211\
        );

    \I__368\ : Span12Mux_v
    port map (
            O => \N__3211\,
            I => \N__3208\
        );

    \I__367\ : Span12Mux_h
    port map (
            O => \N__3208\,
            I => \N__3205\
        );

    \I__366\ : Odrv12
    port map (
            O => \N__3205\,
            I => \N_69_i\
        );

    \I__365\ : InMux
    port map (
            O => \N__3202\,
            I => \N__3199\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3199\,
            I => \N__3196\
        );

    \I__363\ : Span4Mux_v
    port map (
            O => \N__3196\,
            I => \N__3193\
        );

    \I__362\ : Odrv4
    port map (
            O => \N__3193\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_13\
        );

    \I__361\ : CascadeMux
    port map (
            O => \N__3190\,
            I => \N_101_cascade_\
        );

    \I__360\ : InMux
    port map (
            O => \N__3187\,
            I => \N__3183\
        );

    \I__359\ : InMux
    port map (
            O => \N__3186\,
            I => \N__3180\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3183\,
            I => \N__3177\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__3180\,
            I => \N__3174\
        );

    \I__356\ : Odrv12
    port map (
            O => \N__3177\,
            I => \N_105\
        );

    \I__355\ : Odrv4
    port map (
            O => \N__3174\,
            I => \N_105\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__3169\,
            I => \N__3166\
        );

    \I__353\ : InMux
    port map (
            O => \N__3166\,
            I => \N__3161\
        );

    \I__352\ : InMux
    port map (
            O => \N__3165\,
            I => \N__3156\
        );

    \I__351\ : InMux
    port map (
            O => \N__3164\,
            I => \N__3156\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__3161\,
            I => \N__3153\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__3156\,
            I => \N__3150\
        );

    \I__348\ : Span4Mux_h
    port map (
            O => \N__3153\,
            I => \N__3146\
        );

    \I__347\ : Span4Mux_v
    port map (
            O => \N__3150\,
            I => \N__3143\
        );

    \I__346\ : InMux
    port map (
            O => \N__3149\,
            I => \N__3140\
        );

    \I__345\ : Span4Mux_h
    port map (
            O => \N__3146\,
            I => \N__3137\
        );

    \I__344\ : Sp12to4
    port map (
            O => \N__3143\,
            I => \N__3132\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3140\,
            I => \N__3132\
        );

    \I__342\ : Sp12to4
    port map (
            O => \N__3137\,
            I => \N__3127\
        );

    \I__341\ : Span12Mux_h
    port map (
            O => \N__3132\,
            I => \N__3127\
        );

    \I__340\ : Span12Mux_v
    port map (
            O => \N__3127\,
            I => \N__3124\
        );

    \I__339\ : Odrv12
    port map (
            O => \N__3124\,
            I => \A_c_16\
        );

    \I__338\ : InMux
    port map (
            O => \N__3121\,
            I => \N__3115\
        );

    \I__337\ : InMux
    port map (
            O => \N__3120\,
            I => \N__3115\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__3115\,
            I => \N__3110\
        );

    \I__335\ : InMux
    port map (
            O => \N__3114\,
            I => \N__3107\
        );

    \I__334\ : InMux
    port map (
            O => \N__3113\,
            I => \N__3104\
        );

    \I__333\ : Span4Mux_h
    port map (
            O => \N__3110\,
            I => \N__3099\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__3107\,
            I => \N__3099\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__3104\,
            I => \N__3096\
        );

    \I__330\ : Span4Mux_v
    port map (
            O => \N__3099\,
            I => \N__3093\
        );

    \I__329\ : Sp12to4
    port map (
            O => \N__3096\,
            I => \N__3090\
        );

    \I__328\ : Sp12to4
    port map (
            O => \N__3093\,
            I => \N__3087\
        );

    \I__327\ : Span12Mux_v
    port map (
            O => \N__3090\,
            I => \N__3084\
        );

    \I__326\ : Span12Mux_v
    port map (
            O => \N__3087\,
            I => \N__3081\
        );

    \I__325\ : Odrv12
    port map (
            O => \N__3084\,
            I => \A_c_17\
        );

    \I__324\ : Odrv12
    port map (
            O => \N__3081\,
            I => \A_c_17\
        );

    \I__323\ : CascadeMux
    port map (
            O => \N__3076\,
            I => \N__3071\
        );

    \I__322\ : CascadeMux
    port map (
            O => \N__3075\,
            I => \N__3068\
        );

    \I__321\ : InMux
    port map (
            O => \N__3074\,
            I => \N__3061\
        );

    \I__320\ : InMux
    port map (
            O => \N__3071\,
            I => \N__3061\
        );

    \I__319\ : InMux
    port map (
            O => \N__3068\,
            I => \N__3061\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__3061\,
            I => \N__3058\
        );

    \I__317\ : Span4Mux_h
    port map (
            O => \N__3058\,
            I => \N__3055\
        );

    \I__316\ : Sp12to4
    port map (
            O => \N__3055\,
            I => \N__3052\
        );

    \I__315\ : Span12Mux_v
    port map (
            O => \N__3052\,
            I => \N__3049\
        );

    \I__314\ : Odrv12
    port map (
            O => \N__3049\,
            I => \A_c_28\
        );

    \I__313\ : CascadeMux
    port map (
            O => \N__3046\,
            I => \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_7_cascade_\
        );

    \I__312\ : CascadeMux
    port map (
            O => \N__3043\,
            I => \N__3040\
        );

    \I__311\ : InMux
    port map (
            O => \N__3040\,
            I => \N__3031\
        );

    \I__310\ : InMux
    port map (
            O => \N__3039\,
            I => \N__3031\
        );

    \I__309\ : InMux
    port map (
            O => \N__3038\,
            I => \N__3031\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__3031\,
            I => \N__3028\
        );

    \I__307\ : Sp12to4
    port map (
            O => \N__3028\,
            I => \N__3025\
        );

    \I__306\ : Span12Mux_v
    port map (
            O => \N__3025\,
            I => \N__3022\
        );

    \I__305\ : Odrv12
    port map (
            O => \N__3022\,
            I => \A_c_29\
        );

    \I__304\ : InMux
    port map (
            O => \N__3019\,
            I => \N__3016\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__3016\,
            I => \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_8\
        );

    \I__302\ : CascadeMux
    port map (
            O => \N__3013\,
            I => \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_9_cascade_\
        );

    \I__301\ : InMux
    port map (
            O => \N__3010\,
            I => \N__3007\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__3007\,
            I => \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_10\
        );

    \I__299\ : IoInMux
    port map (
            O => \N__3004\,
            I => \N__3001\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__3001\,
            I => \N__2998\
        );

    \I__297\ : Span4Mux_s3_v
    port map (
            O => \N__2998\,
            I => \N__2995\
        );

    \I__296\ : Sp12to4
    port map (
            O => \N__2995\,
            I => \N__2992\
        );

    \I__295\ : Span12Mux_h
    port map (
            O => \N__2992\,
            I => \N__2989\
        );

    \I__294\ : Span12Mux_h
    port map (
            O => \N__2989\,
            I => \N__2986\
        );

    \I__293\ : Odrv12
    port map (
            O => \N__2986\,
            I => \N_31_i\
        );

    \I__292\ : InMux
    port map (
            O => \N__2983\,
            I => \N__2978\
        );

    \I__291\ : InMux
    port map (
            O => \N__2982\,
            I => \N__2973\
        );

    \I__290\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2973\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2978\,
            I => \N__2970\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2973\,
            I => \N__2967\
        );

    \I__287\ : Span4Mux_v
    port map (
            O => \N__2970\,
            I => \N__2964\
        );

    \I__286\ : Span4Mux_v
    port map (
            O => \N__2967\,
            I => \N__2961\
        );

    \I__285\ : Span4Mux_v
    port map (
            O => \N__2964\,
            I => \N__2958\
        );

    \I__284\ : Span4Mux_v
    port map (
            O => \N__2961\,
            I => \N__2955\
        );

    \I__283\ : Span4Mux_h
    port map (
            O => \N__2958\,
            I => \N__2952\
        );

    \I__282\ : Span4Mux_h
    port map (
            O => \N__2955\,
            I => \N__2949\
        );

    \I__281\ : Odrv4
    port map (
            O => \N__2952\,
            I => \A_c_31\
        );

    \I__280\ : Odrv4
    port map (
            O => \N__2949\,
            I => \A_c_31\
        );

    \I__279\ : CascadeMux
    port map (
            O => \N__2944\,
            I => \N__2941\
        );

    \I__278\ : InMux
    port map (
            O => \N__2941\,
            I => \N__2938\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2938\,
            I => \N__2935\
        );

    \I__276\ : Span12Mux_v
    port map (
            O => \N__2935\,
            I => \N__2932\
        );

    \I__275\ : Odrv12
    port map (
            O => \N__2932\,
            I => \TT_c_1\
        );

    \I__274\ : CascadeMux
    port map (
            O => \N__2929\,
            I => \N__2924\
        );

    \I__273\ : InMux
    port map (
            O => \N__2928\,
            I => \N__2921\
        );

    \I__272\ : InMux
    port map (
            O => \N__2927\,
            I => \N__2918\
        );

    \I__271\ : InMux
    port map (
            O => \N__2924\,
            I => \N__2915\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2921\,
            I => \N__2910\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__2918\,
            I => \N__2910\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2915\,
            I => \N__2905\
        );

    \I__267\ : Sp12to4
    port map (
            O => \N__2910\,
            I => \N__2905\
        );

    \I__266\ : Span12Mux_v
    port map (
            O => \N__2905\,
            I => \N__2902\
        );

    \I__265\ : Odrv12
    port map (
            O => \N__2902\,
            I => \A_c_30\
        );

    \I__264\ : ClkMux
    port map (
            O => \N__2899\,
            I => \N__2857\
        );

    \I__263\ : ClkMux
    port map (
            O => \N__2898\,
            I => \N__2857\
        );

    \I__262\ : ClkMux
    port map (
            O => \N__2897\,
            I => \N__2857\
        );

    \I__261\ : ClkMux
    port map (
            O => \N__2896\,
            I => \N__2857\
        );

    \I__260\ : ClkMux
    port map (
            O => \N__2895\,
            I => \N__2857\
        );

    \I__259\ : ClkMux
    port map (
            O => \N__2894\,
            I => \N__2857\
        );

    \I__258\ : ClkMux
    port map (
            O => \N__2893\,
            I => \N__2857\
        );

    \I__257\ : ClkMux
    port map (
            O => \N__2892\,
            I => \N__2857\
        );

    \I__256\ : ClkMux
    port map (
            O => \N__2891\,
            I => \N__2857\
        );

    \I__255\ : ClkMux
    port map (
            O => \N__2890\,
            I => \N__2857\
        );

    \I__254\ : ClkMux
    port map (
            O => \N__2889\,
            I => \N__2857\
        );

    \I__253\ : ClkMux
    port map (
            O => \N__2888\,
            I => \N__2857\
        );

    \I__252\ : ClkMux
    port map (
            O => \N__2887\,
            I => \N__2857\
        );

    \I__251\ : ClkMux
    port map (
            O => \N__2886\,
            I => \N__2857\
        );

    \I__250\ : GlobalMux
    port map (
            O => \N__2857\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            I => \N__2892\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            I => \N__2897\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            I => \N__2890\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            I => \N__2888\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            I => \N__2886\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            I => \N__2899\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            I => \N__2898\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            I => \N__2896\
        );

    \INVU409_TRANSFER_ACK.TACK_EN_iC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            I => \N__2894\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__2891\
        );

    \INVU409_TRANSFER_ACK.CIA_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            I => \N__2889\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\,
            I => \N__2887\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            I => \N__2895\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\,
            I => \N__2893\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_15_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_3_0_\
        );

    \IN_MUX_bfv_15_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_15_4_0_\
        );

    \IN_MUX_bfv_15_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_6_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3149\,
            in2 => \_gnd_net_\,
            in3 => \N__3114\,
            lcout => \N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_7_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__3074\,
            in1 => \_gnd_net_\,
            in2 => \N__3043\,
            in3 => \N__3390\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_4_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3039\,
            in1 => \N__2982\,
            in2 => \N__3076\,
            in3 => \N__2927\,
            lcout => \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.un1_BUFENn_i_a4_7_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3186\,
            in1 => \N__4207\,
            in2 => \N__3075\,
            in3 => \N__2981\,
            lcout => OPEN,
            ltout => \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.un1_BUFENn_i_a4_10_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__3345\,
            in1 => \_gnd_net_\,
            in2 => \N__3046\,
            in3 => \N__3038\,
            lcout => \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.un1_BUFENn_i_a4_8_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__3445\,
            in1 => \N__3577\,
            in2 => \N__2929\,
            in3 => \N__5340\,
            lcout => \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.un1_BUFENn_i_a4_9_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3999\,
            in1 => \N__3386\,
            in2 => \N__3280\,
            in3 => \N__3320\,
            lcout => OPEN,
            ltout => \U409_DATA_BUFFERS.un1_BUFENn_i_a4Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.N_31_i_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__4033\,
            in1 => \N__3019\,
            in2 => \N__3013\,
            in3 => \N__3010\,
            lcout => \N_31_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_10_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2983\,
            in1 => \N__3902\,
            in2 => \N__2944\,
            in3 => \N__2928\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3608\,
            in1 => \N__3627\,
            in2 => \_gnd_net_\,
            in3 => \N__5339\,
            lcout => \U409_ADDRESS_DECODE_Z2_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_5_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3391\,
            in1 => \N__3351\,
            in2 => \N__3321\,
            in3 => \N__3278\,
            lcout => \U409_TRANSFER_ACK_DELAYED_TACK_RST_1_i_a2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_8_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3535\,
            in1 => \N__3352\,
            in2 => \N__3322\,
            in3 => \N__3279\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_LC_3_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3244\,
            in1 => \N__3472\,
            in2 => \N__3235\,
            in3 => \N__3232\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.N_69_i_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__3513\,
            in1 => \N__3113\,
            in2 => \N__3169\,
            in3 => \N__3739\,
            lcout => \N_69_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3457\,
            in1 => \N__4015\,
            in2 => \_gnd_net_\,
            in3 => \N__3578\,
            lcout => \N_101\,
            ltout => \N_101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__3738\,
            in1 => \N__3202\,
            in2 => \N__3190\,
            in3 => \N__3187\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a4_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3120\,
            in1 => \N__3729\,
            in2 => \N__3512\,
            in3 => \N__3164\,
            lcout => \U409_ADDRESS_DECODE.N_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_1_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3165\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3121\,
            lcout => \N_74_1\,
            ltout => \N_74_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_o2_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001100110011"
        )
    port map (
            in0 => \N__3458\,
            in1 => \N__4000\,
            in2 => \N__3652\,
            in3 => \N__3579\,
            lcout => \N_33\,
            ltout => \N_33_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a4_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3646\,
            in1 => \N__3640\,
            in2 => \N__3649\,
            in3 => \N__3613\,
            lcout => \U409_TRANSFER_ACK.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_1_i_a2_0_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3922\,
            in1 => \N__3399\,
            in2 => \N__3805\,
            in3 => \N__3763\,
            lcout => \N_99\,
            ltout => \N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3639\,
            in1 => \N__5335\,
            in2 => \N__3616\,
            in3 => \N__3609\,
            lcout => \N_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3580\,
            in1 => \N__3459\,
            in2 => \N__3531\,
            in3 => \N__3868\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15_9_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3400\,
            in1 => \N__3514\,
            in2 => \N__5341\,
            in3 => \N__3487\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a4_0_15Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_1_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3831\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4014\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.HIROMZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3460\,
            in1 => \N__3870\,
            in2 => \N__3403\,
            in3 => \N__3921\,
            lcout => \U409_ADDRESS_DECODE_HIROM\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3832\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3869\,
            lcout => \U409_TRANSFER_ACK.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.un1_BUFENn_i_0_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__3730\,
            in1 => \N__3696\,
            in2 => \_gnd_net_\,
            in3 => \N__4144\,
            lcout => \U409_DATA_BUFFERS.un1_BUFENn_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3802\,
            in1 => \N__3923\,
            in2 => \N__4024\,
            in3 => \N__3764\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4057\,
            in1 => \N__4007\,
            in2 => \N__3961\,
            in3 => \N__3833\,
            lcout => \CIA_SPACE\,
            ltout => \CIA_SPACE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__3692\,
            in1 => \N__3728\,
            in2 => \N__3958\,
            in3 => \N__3955\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un5_RAMSPACEn_0_a2_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__3925\,
            in1 => \_gnd_net_\,
            in2 => \N__3883\,
            in3 => \N__3835\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.un5_RAMSPACEn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a2_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__3803\,
            in1 => \_gnd_net_\,
            in2 => \N__3928\,
            in3 => \N__3765\,
            lcout => \N_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.LOWROM_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__3924\,
            in1 => \N__4180\,
            in2 => \N__3882\,
            in3 => \N__3834\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE_LOWROM_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_1_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010010101000"
        )
    port map (
            in0 => \N__3804\,
            in1 => \N__3775\,
            in2 => \N__3769\,
            in3 => \N__3766\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER15Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.N_68_i_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__3734\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3697\,
            lcout => \N_68_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__4137\,
            in1 => \N__4264\,
            in2 => \N__4255\,
            in3 => \N__5328\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.N_67_i_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__4172\,
            in1 => \N__4061\,
            in2 => \_gnd_net_\,
            in3 => \N__4199\,
            lcout => \N_67_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a4_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4062\,
            in1 => \N__4200\,
            in2 => \_gnd_net_\,
            in3 => \N__4173\,
            lcout => \N_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4314\,
            in2 => \_gnd_net_\,
            in3 => \N__4290\,
            lcout => \U409_TRANSFER_ACK.CO1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__4084\,
            in1 => \N__4095\,
            in2 => \N__4126\,
            in3 => \N__4564\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5650\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4942\,
            in1 => \N__4096\,
            in2 => \N__4122\,
            in3 => \N__4878\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4938\,
            in2 => \_gnd_net_\,
            in3 => \N__4871\,
            lcout => \U409_TRANSFER_ACK.N_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4075\,
            in1 => \N__4063\,
            in2 => \N__4918\,
            in3 => \N__4859\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_3_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4287\,
            in1 => \N__4717\,
            in2 => \N__4696\,
            in3 => \N__4311\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\,
            ltout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIERIJ7_3_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4401\,
            in2 => \N__4411\,
            in3 => \N__4359\,
            lcout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0\,
            ltout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__4288\,
            in1 => \_gnd_net_\,
            in2 => \N__4408\,
            in3 => \N__4313\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__5640\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_3_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4312\,
            in1 => \N__4689\,
            in2 => \N__4720\,
            in3 => \N__4286\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010101"
        )
    port map (
            in0 => \N__4289\,
            in1 => \_gnd_net_\,
            in2 => \N__4405\,
            in3 => \N__4371\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__5640\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001001100"
        )
    port map (
            in0 => \N__5123\,
            in1 => \N__4552\,
            in2 => \N__5152\,
            in3 => \N__4651\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5649\
        );

    \U409_TRANSFER_ACK.ROMENn_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101101110000"
        )
    port map (
            in0 => \N__4400\,
            in1 => \N__4372\,
            in2 => \N__4332\,
            in3 => \N__4360\,
            lcout => \ROMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5649\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4740\,
            in2 => \_gnd_net_\,
            in3 => \N__4694\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5649\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101000101010"
        )
    port map (
            in0 => \N__4539\,
            in1 => \N__4315\,
            in2 => \N__4666\,
            in3 => \N__4291\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5649\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011111110111"
        )
    port map (
            in0 => \N__5074\,
            in1 => \N__5094\,
            in2 => \N__5128\,
            in3 => \N__4650\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001010001010"
        )
    port map (
            in0 => \N__5276\,
            in1 => \N__5151\,
            in2 => \N__4567\,
            in3 => \N__4657\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001000100"
        )
    port map (
            in0 => \N__4461\,
            in1 => \N__5277\,
            in2 => \N__4492\,
            in3 => \N__4440\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4563\,
            in1 => \N__4551\,
            in2 => \N__4540\,
            in3 => \N__4639\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER6\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100110111"
        )
    port map (
            in0 => \N__4459\,
            in1 => \N__5279\,
            in2 => \N__4525\,
            in3 => \N__4482\,
            lcout => \U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__5278\,
            in1 => \N__4486\,
            in2 => \_gnd_net_\,
            in3 => \N__4460\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100111"
        )
    port map (
            in0 => \N__4458\,
            in1 => \N__4505\,
            in2 => \N__4491\,
            in3 => \N__4439\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__4506\,
            in1 => \_gnd_net_\,
            in2 => \N__4522\,
            in3 => \N__5291\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__4490\,
            in1 => \N__4462\,
            in2 => \N__5312\,
            in3 => \N__4441\,
            lcout => \TACK_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            ce => \N__4426\,
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__4638\,
            in1 => \N__4788\,
            in2 => \_gnd_net_\,
            in3 => \N__4615\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5466\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4594\,
            in1 => \N__4577\,
            in2 => \N__5023\,
            in3 => \N__5044\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__5516\,
            in1 => \N__4986\,
            in2 => \N__4624\,
            in3 => \N__5055\,
            lcout => \U409_TRANSFER_ACK.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4578\,
            in1 => \N__5019\,
            in2 => \N__4600\,
            in3 => \N__5045\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5056\,
            in1 => \N__4985\,
            in2 => \N__4621\,
            in3 => \N__5515\,
            lcout => \U409_TRANSFER_ACK.N_70\,
            ltout => \U409_TRANSFER_ACK.N_70_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_3_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011111111"
        )
    port map (
            in0 => \N__4861\,
            in1 => \N__4931\,
            in2 => \N__4618\,
            in3 => \N__4614\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4599\,
            in2 => \N__4603\,
            in3 => \N__4950\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__5467\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__4579\,
            in1 => \N__4595\,
            in2 => \N__4954\,
            in3 => \N__5573\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__5467\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__4776\,
            in1 => \N__4991\,
            in2 => \_gnd_net_\,
            in3 => \N__5568\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__5452\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__4992\,
            in1 => \N__4777\,
            in2 => \N__5575\,
            in3 => \N__5022\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__5452\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5518\,
            in1 => \N__5487\,
            in2 => \_gnd_net_\,
            in3 => \N__5545\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__4765\,
            in1 => \N__5047\,
            in2 => \N__4768\,
            in3 => \N__5569\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__5452\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4990\,
            in2 => \_gnd_net_\,
            in3 => \N__5021\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__4719\,
            in1 => \N__4695\,
            in2 => \N__4744\,
            in3 => \N__4726\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__5624\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4718\,
            in2 => \_gnd_net_\,
            in3 => \N__4693\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_EN_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__5073\,
            in1 => \N__5092\,
            in2 => \N__5124\,
            in3 => \N__5161\,
            lcout => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIA48I_1_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4840\,
            in1 => \N__5170\,
            in2 => \_gnd_net_\,
            in3 => \N__5184\,
            lcout => \U409_TRANSFER_ACK.N_17_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5169\,
            in2 => \_gnd_net_\,
            in3 => \N__5183\,
            lcout => \U409_TRANSFER_ACK.N_3_0\,
            ltout => \U409_TRANSFER_ACK.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100100111"
        )
    port map (
            in0 => \N__5115\,
            in1 => \N__5093\,
            in2 => \N__5155\,
            in3 => \N__5072\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.N_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101000001000"
        )
    port map (
            in0 => \N__5269\,
            in1 => \N__5150\,
            in2 => \N__5131\,
            in3 => \N__5119\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5249\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6795\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__5645\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5095\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__5645\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5548\,
            in3 => \N__5485\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5046\,
            in1 => \N__5020\,
            in2 => \N__4993\,
            in3 => \N__5486\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5517\,
            in2 => \N__4957\,
            in3 => \N__5544\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110000110011"
        )
    port map (
            in0 => \N__4930\,
            in1 => \N__5519\,
            in2 => \N__4860\,
            in3 => \N__4789\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5462\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5520\,
            in1 => \N__5546\,
            in2 => \_gnd_net_\,
            in3 => \N__5574\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5462\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__5547\,
            in1 => \N__5521\,
            in2 => \_gnd_net_\,
            in3 => \N__5488\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5462\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5428\,
            in2 => \_gnd_net_\,
            in3 => \N__5350\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5349\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5389\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNI692L_0_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5267\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6796\,
            lcout => \CIA_ENABLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5268\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6843\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__5641\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5185\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__5641\
        );

    \U409_TICK.COUNTER60_9_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5699\,
            in1 => \N__5733\,
            in2 => \N__5776\,
            in3 => \N__6238\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6460\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6007\,
            in1 => \N__6031\,
            in2 => \_gnd_net_\,
            in3 => \N__6085\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6214\,
            in1 => \N__5587\,
            in2 => \N__5593\,
            in3 => \N__6046\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__6019\,
            in1 => \N__5700\,
            in2 => \N__5590\,
            in3 => \N__5774\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6460\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5698\,
            in1 => \N__5732\,
            in2 => \N__5775\,
            in3 => \N__6157\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6460\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6199\,
            in1 => \N__6061\,
            in2 => \N__6112\,
            in3 => \N__6123\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__6184\,
            in1 => \N__6229\,
            in2 => \N__5965\,
            in3 => \N__6148\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5731\,
            in1 => \N__5773\,
            in2 => \N__5581\,
            in3 => \N__6136\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6460\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__6526\,
            in1 => \N__6499\,
            in2 => \N__6355\,
            in3 => \N__6280\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_14_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5845\,
            in1 => \N__5908\,
            in2 => \N__5578\,
            in3 => \N__6487\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6456\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_14_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__5909\,
            in1 => \N__5874\,
            in2 => \N__6322\,
            in3 => \N__5849\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6456\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_14_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6432\,
            in2 => \_gnd_net_\,
            in3 => \N__6413\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6456\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6265\,
            in1 => \N__6385\,
            in2 => \N__6433\,
            in3 => \N__6474\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_14_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__5876\,
            in1 => \N__5664\,
            in2 => \N__5851\,
            in3 => \N__5911\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6456\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_14_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__5910\,
            in1 => \N__5875\,
            in2 => \N__6295\,
            in3 => \N__5850\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6456\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5878\,
            in1 => \N__5905\,
            in2 => \N__5843\,
            in3 => \N__6571\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6583\,
            in1 => \N__6619\,
            in2 => \N__6310\,
            in3 => \N__6547\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__5877\,
            in1 => \N__6415\,
            in2 => \N__5653\,
            in3 => \N__5904\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6370\,
            in1 => \N__6336\,
            in2 => \_gnd_net_\,
            in3 => \N__6409\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5923\,
            in1 => \N__6562\,
            in2 => \N__5917\,
            in3 => \N__6598\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5842\,
            in1 => \N__5881\,
            in2 => \N__5914\,
            in3 => \N__6607\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5879\,
            in1 => \N__5906\,
            in2 => \N__5844\,
            in3 => \N__6535\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__5907\,
            in1 => \N__5880\,
            in2 => \N__6514\,
            in3 => \N__5832\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5734\,
            in1 => \N__5766\,
            in2 => \N__5707\,
            in3 => \N__5932\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__5765\,
            in1 => \N__5790\,
            in2 => \N__5743\,
            in3 => \N__5702\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6250\,
            in1 => \N__5944\,
            in2 => \N__5992\,
            in3 => \N__6169\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__5974\,
            in1 => \N__5701\,
            in2 => \N__5779\,
            in3 => \N__5736\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__5764\,
            in1 => \N__5735\,
            in2 => \N__6091\,
            in3 => \N__5706\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6086\,
            in2 => \_gnd_net_\,
            in3 => \N__6111\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6461\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6107\,
            in2 => \N__6090\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6060\,
            in2 => \_gnd_net_\,
            in3 => \N__6049\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__6462\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6045\,
            in2 => \_gnd_net_\,
            in3 => \N__6034\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__6462\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6030\,
            in2 => \_gnd_net_\,
            in3 => \N__6010\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6006\,
            in2 => \_gnd_net_\,
            in3 => \N__5995\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__6462\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5991\,
            in3 => \N__5968\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5958\,
            in2 => \_gnd_net_\,
            in3 => \N__5947\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__6462\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5943\,
            in2 => \_gnd_net_\,
            in3 => \N__5926\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6249\,
            in2 => \_gnd_net_\,
            in3 => \N__6232\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6228\,
            in2 => \_gnd_net_\,
            in3 => \N__6217\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__6463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6213\,
            in2 => \_gnd_net_\,
            in3 => \N__6202\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__6463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6198\,
            in2 => \_gnd_net_\,
            in3 => \N__6187\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__6463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6183\,
            in2 => \_gnd_net_\,
            in3 => \N__6172\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__6463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6168\,
            in2 => \_gnd_net_\,
            in3 => \N__6151\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6147\,
            in2 => \_gnd_net_\,
            in3 => \N__6130\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6124\,
            in2 => \_gnd_net_\,
            in3 => \N__6127\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6428\,
            in2 => \N__6414\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_3_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_15_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6384\,
            in2 => \_gnd_net_\,
            in3 => \N__6373\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__6458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6369\,
            in2 => \_gnd_net_\,
            in3 => \N__6358\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__6458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_15_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6351\,
            in2 => \_gnd_net_\,
            in3 => \N__6340\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__6458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_15_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6337\,
            in3 => \N__6313\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6306\,
            in2 => \_gnd_net_\,
            in3 => \N__6283\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_15_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6279\,
            in2 => \_gnd_net_\,
            in3 => \N__6268\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__6458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_15_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6264\,
            in2 => \_gnd_net_\,
            in3 => \N__6253\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__6458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6618\,
            in2 => \_gnd_net_\,
            in3 => \N__6601\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_4_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6597\,
            in2 => \_gnd_net_\,
            in3 => \N__6586\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__6459\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6582\,
            in2 => \_gnd_net_\,
            in3 => \N__6565\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6561\,
            in2 => \_gnd_net_\,
            in3 => \N__6550\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__6459\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6546\,
            in2 => \_gnd_net_\,
            in3 => \N__6529\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6525\,
            in2 => \_gnd_net_\,
            in3 => \N__6502\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6498\,
            in2 => \_gnd_net_\,
            in3 => \N__6481\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6475\,
            in2 => \_gnd_net_\,
            in3 => \N__6478\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6459\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6969\,
            in2 => \N__7003\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_6_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6753\,
            in2 => \_gnd_net_\,
            in3 => \N__6655\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__6940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__6765\,
            in1 => \_gnd_net_\,
            in2 => \N__6637\,
            in3 => \N__6652\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \N__6940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6702\,
            in2 => \_gnd_net_\,
            in3 => \N__6649\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__6940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6766\,
            in1 => \N__6730\,
            in2 => \_gnd_net_\,
            in3 => \N__6646\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            clk => \N__6940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_6_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6873\,
            in2 => \_gnd_net_\,
            in3 => \N__6643\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\,
            clk => \N__6940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_7_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6891\,
            in2 => \_gnd_net_\,
            in3 => \N__6640\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6940\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6890\,
            in1 => \N__6872\,
            in2 => \_gnd_net_\,
            in3 => \N__6632\,
            lcout => \U409_CIA.N_104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_2_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6994\,
            in1 => \N__6700\,
            in2 => \_gnd_net_\,
            in3 => \N__6636\,
            lcout => OPEN,
            ltout => \U409_CIA.un1_CIA_CLK_COUNT_2_0_a4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_1_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6709\,
            in1 => \N__6892\,
            in2 => \N__6877\,
            in3 => \N__6874\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA_RNOZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6661\,
            in2 => \N__6859\,
            in3 => \N__6836\,
            lcout => \CLK_CIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_1_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__6701\,
            in1 => \_gnd_net_\,
            in2 => \N__6970\,
            in3 => \N__6995\,
            lcout => OPEN,
            ltout => \U409_CIA.un1_CIA_CLK_COUNT_3_0_a4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6675\,
            in1 => \N__6757\,
            in2 => \N__6820\,
            in3 => \N__6728\,
            lcout => OPEN,
            ltout => \U409_CIA.VMA_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__6817\,
            in1 => \N__6782\,
            in2 => \N__6799\,
            in3 => \N__6997\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6938\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6752\,
            in1 => \N__6727\,
            in2 => \_gnd_net_\,
            in3 => \N__6699\,
            lcout => OPEN,
            ltout => \U409_CIA.CIA_CLK_COUNT11_0_a4_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6968\,
            in1 => \N__6996\,
            in2 => \N__6769\,
            in3 => \N__6674\,
            lcout => \U409_CIA.CIA_CLK_COUNT11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNID3921_2_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6962\,
            in1 => \N__6751\,
            in2 => \_gnd_net_\,
            in3 => \N__6729\,
            lcout => \U409_CIA.CLK_CIA6_1\,
            ltout => \U409_CIA.CLK_CIA6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_0_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__7001\,
            in1 => \N__6703\,
            in2 => \N__6679\,
            in3 => \N__6676\,
            lcout => \U409_CIA.CLK_CIA6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__6964\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7002\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6939\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6963\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6939\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_iobuf_RNO_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6925\,
            lcout => \N_465_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jul 2 2025 17:00:31

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    CMA,
    DRA,
    DA,
    A,
    TBIn,
    RAMSPACEn,
    DBRn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    PRnW,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    BLSn,
    TCIn,
    WEn,
    REGENn,
    LLBEn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    output [10:0] CMA;
    input [9:0] DRA;
    output [2:0] DA;
    input [20:0] A;
    output TBIn;
    input RAMSPACEn;
    input DBRn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output PRnW;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    output BLSn;
    output TCIn;
    output WEn;
    output REGENn;
    output LLBEn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__13257;
    wire N__13256;
    wire N__13255;
    wire N__13248;
    wire N__13247;
    wire N__13246;
    wire N__13239;
    wire N__13238;
    wire N__13237;
    wire N__13230;
    wire N__13229;
    wire N__13228;
    wire N__13221;
    wire N__13220;
    wire N__13219;
    wire N__13212;
    wire N__13211;
    wire N__13210;
    wire N__13203;
    wire N__13202;
    wire N__13201;
    wire N__13194;
    wire N__13193;
    wire N__13192;
    wire N__13185;
    wire N__13184;
    wire N__13183;
    wire N__13176;
    wire N__13175;
    wire N__13174;
    wire N__13167;
    wire N__13166;
    wire N__13165;
    wire N__13158;
    wire N__13157;
    wire N__13156;
    wire N__13149;
    wire N__13148;
    wire N__13147;
    wire N__13140;
    wire N__13139;
    wire N__13138;
    wire N__13131;
    wire N__13130;
    wire N__13129;
    wire N__13122;
    wire N__13121;
    wire N__13120;
    wire N__13113;
    wire N__13112;
    wire N__13111;
    wire N__13104;
    wire N__13103;
    wire N__13102;
    wire N__13095;
    wire N__13094;
    wire N__13093;
    wire N__13086;
    wire N__13085;
    wire N__13084;
    wire N__13077;
    wire N__13076;
    wire N__13075;
    wire N__13068;
    wire N__13067;
    wire N__13066;
    wire N__13059;
    wire N__13058;
    wire N__13057;
    wire N__13050;
    wire N__13049;
    wire N__13048;
    wire N__13041;
    wire N__13040;
    wire N__13039;
    wire N__13032;
    wire N__13031;
    wire N__13030;
    wire N__13023;
    wire N__13022;
    wire N__13021;
    wire N__13014;
    wire N__13013;
    wire N__13012;
    wire N__13005;
    wire N__13004;
    wire N__13003;
    wire N__12996;
    wire N__12995;
    wire N__12994;
    wire N__12987;
    wire N__12986;
    wire N__12985;
    wire N__12978;
    wire N__12977;
    wire N__12976;
    wire N__12969;
    wire N__12968;
    wire N__12967;
    wire N__12960;
    wire N__12959;
    wire N__12958;
    wire N__12951;
    wire N__12950;
    wire N__12949;
    wire N__12942;
    wire N__12941;
    wire N__12940;
    wire N__12933;
    wire N__12932;
    wire N__12931;
    wire N__12924;
    wire N__12923;
    wire N__12922;
    wire N__12915;
    wire N__12914;
    wire N__12913;
    wire N__12906;
    wire N__12905;
    wire N__12904;
    wire N__12897;
    wire N__12896;
    wire N__12895;
    wire N__12888;
    wire N__12887;
    wire N__12886;
    wire N__12879;
    wire N__12878;
    wire N__12877;
    wire N__12870;
    wire N__12869;
    wire N__12868;
    wire N__12861;
    wire N__12860;
    wire N__12859;
    wire N__12852;
    wire N__12851;
    wire N__12850;
    wire N__12843;
    wire N__12842;
    wire N__12841;
    wire N__12834;
    wire N__12833;
    wire N__12832;
    wire N__12825;
    wire N__12824;
    wire N__12823;
    wire N__12816;
    wire N__12815;
    wire N__12814;
    wire N__12807;
    wire N__12806;
    wire N__12805;
    wire N__12798;
    wire N__12797;
    wire N__12796;
    wire N__12789;
    wire N__12788;
    wire N__12787;
    wire N__12780;
    wire N__12779;
    wire N__12778;
    wire N__12771;
    wire N__12770;
    wire N__12769;
    wire N__12762;
    wire N__12761;
    wire N__12760;
    wire N__12753;
    wire N__12752;
    wire N__12751;
    wire N__12744;
    wire N__12743;
    wire N__12742;
    wire N__12735;
    wire N__12734;
    wire N__12733;
    wire N__12726;
    wire N__12725;
    wire N__12724;
    wire N__12717;
    wire N__12716;
    wire N__12715;
    wire N__12708;
    wire N__12707;
    wire N__12706;
    wire N__12699;
    wire N__12698;
    wire N__12697;
    wire N__12690;
    wire N__12689;
    wire N__12688;
    wire N__12681;
    wire N__12680;
    wire N__12679;
    wire N__12672;
    wire N__12671;
    wire N__12670;
    wire N__12663;
    wire N__12662;
    wire N__12661;
    wire N__12654;
    wire N__12653;
    wire N__12652;
    wire N__12645;
    wire N__12644;
    wire N__12643;
    wire N__12636;
    wire N__12635;
    wire N__12634;
    wire N__12627;
    wire N__12626;
    wire N__12625;
    wire N__12618;
    wire N__12617;
    wire N__12616;
    wire N__12609;
    wire N__12608;
    wire N__12607;
    wire N__12600;
    wire N__12599;
    wire N__12598;
    wire N__12591;
    wire N__12590;
    wire N__12589;
    wire N__12582;
    wire N__12581;
    wire N__12580;
    wire N__12573;
    wire N__12572;
    wire N__12571;
    wire N__12564;
    wire N__12563;
    wire N__12562;
    wire N__12555;
    wire N__12554;
    wire N__12553;
    wire N__12546;
    wire N__12545;
    wire N__12544;
    wire N__12537;
    wire N__12536;
    wire N__12535;
    wire N__12528;
    wire N__12527;
    wire N__12526;
    wire N__12519;
    wire N__12518;
    wire N__12517;
    wire N__12510;
    wire N__12509;
    wire N__12508;
    wire N__12501;
    wire N__12500;
    wire N__12499;
    wire N__12492;
    wire N__12491;
    wire N__12490;
    wire N__12483;
    wire N__12482;
    wire N__12481;
    wire N__12474;
    wire N__12473;
    wire N__12472;
    wire N__12465;
    wire N__12464;
    wire N__12463;
    wire N__12456;
    wire N__12455;
    wire N__12454;
    wire N__12447;
    wire N__12446;
    wire N__12445;
    wire N__12438;
    wire N__12437;
    wire N__12436;
    wire N__12429;
    wire N__12428;
    wire N__12427;
    wire N__12420;
    wire N__12419;
    wire N__12418;
    wire N__12411;
    wire N__12410;
    wire N__12409;
    wire N__12402;
    wire N__12401;
    wire N__12400;
    wire N__12393;
    wire N__12392;
    wire N__12391;
    wire N__12374;
    wire N__12371;
    wire N__12368;
    wire N__12365;
    wire N__12362;
    wire N__12359;
    wire N__12358;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12350;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12332;
    wire N__12331;
    wire N__12330;
    wire N__12329;
    wire N__12326;
    wire N__12325;
    wire N__12324;
    wire N__12321;
    wire N__12320;
    wire N__12319;
    wire N__12318;
    wire N__12315;
    wire N__12314;
    wire N__12311;
    wire N__12308;
    wire N__12307;
    wire N__12306;
    wire N__12305;
    wire N__12304;
    wire N__12301;
    wire N__12298;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12286;
    wire N__12283;
    wire N__12278;
    wire N__12275;
    wire N__12268;
    wire N__12265;
    wire N__12262;
    wire N__12257;
    wire N__12252;
    wire N__12249;
    wire N__12246;
    wire N__12243;
    wire N__12232;
    wire N__12229;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12194;
    wire N__12191;
    wire N__12188;
    wire N__12185;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12175;
    wire N__12174;
    wire N__12173;
    wire N__12170;
    wire N__12167;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12155;
    wire N__12152;
    wire N__12149;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12121;
    wire N__12120;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12093;
    wire N__12090;
    wire N__12085;
    wire N__12082;
    wire N__12079;
    wire N__12076;
    wire N__12071;
    wire N__12070;
    wire N__12069;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12051;
    wire N__12046;
    wire N__12043;
    wire N__12040;
    wire N__12037;
    wire N__12034;
    wire N__12031;
    wire N__12026;
    wire N__12023;
    wire N__12020;
    wire N__12017;
    wire N__12014;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12006;
    wire N__12005;
    wire N__12000;
    wire N__11995;
    wire N__11992;
    wire N__11989;
    wire N__11986;
    wire N__11983;
    wire N__11980;
    wire N__11977;
    wire N__11974;
    wire N__11969;
    wire N__11966;
    wire N__11965;
    wire N__11964;
    wire N__11961;
    wire N__11958;
    wire N__11955;
    wire N__11948;
    wire N__11947;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11935;
    wire N__11932;
    wire N__11929;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11902;
    wire N__11899;
    wire N__11896;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11885;
    wire N__11880;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11868;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11837;
    wire N__11836;
    wire N__11835;
    wire N__11832;
    wire N__11831;
    wire N__11830;
    wire N__11829;
    wire N__11828;
    wire N__11827;
    wire N__11824;
    wire N__11823;
    wire N__11820;
    wire N__11819;
    wire N__11816;
    wire N__11813;
    wire N__11812;
    wire N__11811;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11801;
    wire N__11800;
    wire N__11799;
    wire N__11798;
    wire N__11795;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11765;
    wire N__11762;
    wire N__11761;
    wire N__11760;
    wire N__11759;
    wire N__11758;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11743;
    wire N__11738;
    wire N__11725;
    wire N__11720;
    wire N__11717;
    wire N__11712;
    wire N__11703;
    wire N__11700;
    wire N__11697;
    wire N__11694;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11668;
    wire N__11665;
    wire N__11660;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11647;
    wire N__11646;
    wire N__11645;
    wire N__11644;
    wire N__11643;
    wire N__11642;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11620;
    wire N__11619;
    wire N__11618;
    wire N__11617;
    wire N__11616;
    wire N__11615;
    wire N__11614;
    wire N__11613;
    wire N__11612;
    wire N__11611;
    wire N__11610;
    wire N__11609;
    wire N__11582;
    wire N__11579;
    wire N__11576;
    wire N__11575;
    wire N__11574;
    wire N__11573;
    wire N__11572;
    wire N__11571;
    wire N__11570;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11549;
    wire N__11546;
    wire N__11545;
    wire N__11544;
    wire N__11541;
    wire N__11540;
    wire N__11539;
    wire N__11538;
    wire N__11537;
    wire N__11536;
    wire N__11535;
    wire N__11534;
    wire N__11533;
    wire N__11532;
    wire N__11531;
    wire N__11530;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11522;
    wire N__11521;
    wire N__11520;
    wire N__11519;
    wire N__11518;
    wire N__11515;
    wire N__11514;
    wire N__11513;
    wire N__11512;
    wire N__11511;
    wire N__11510;
    wire N__11509;
    wire N__11508;
    wire N__11507;
    wire N__11506;
    wire N__11505;
    wire N__11502;
    wire N__11501;
    wire N__11500;
    wire N__11499;
    wire N__11496;
    wire N__11495;
    wire N__11494;
    wire N__11493;
    wire N__11492;
    wire N__11491;
    wire N__11490;
    wire N__11489;
    wire N__11488;
    wire N__11485;
    wire N__11484;
    wire N__11483;
    wire N__11482;
    wire N__11481;
    wire N__11480;
    wire N__11479;
    wire N__11478;
    wire N__11477;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11359;
    wire N__11358;
    wire N__11357;
    wire N__11356;
    wire N__11353;
    wire N__11352;
    wire N__11351;
    wire N__11350;
    wire N__11349;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11338;
    wire N__11335;
    wire N__11334;
    wire N__11333;
    wire N__11332;
    wire N__11325;
    wire N__11318;
    wire N__11317;
    wire N__11316;
    wire N__11313;
    wire N__11308;
    wire N__11305;
    wire N__11302;
    wire N__11301;
    wire N__11300;
    wire N__11295;
    wire N__11292;
    wire N__11291;
    wire N__11290;
    wire N__11285;
    wire N__11280;
    wire N__11271;
    wire N__11266;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11258;
    wire N__11253;
    wire N__11252;
    wire N__11251;
    wire N__11250;
    wire N__11249;
    wire N__11248;
    wire N__11247;
    wire N__11246;
    wire N__11245;
    wire N__11244;
    wire N__11243;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11231;
    wire N__11226;
    wire N__11223;
    wire N__11218;
    wire N__11209;
    wire N__11206;
    wire N__11197;
    wire N__11196;
    wire N__11195;
    wire N__11194;
    wire N__11193;
    wire N__11192;
    wire N__11187;
    wire N__11178;
    wire N__11175;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11144;
    wire N__11141;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11074;
    wire N__11071;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11056;
    wire N__11055;
    wire N__11054;
    wire N__11053;
    wire N__11052;
    wire N__11051;
    wire N__11050;
    wire N__11049;
    wire N__11048;
    wire N__11047;
    wire N__11046;
    wire N__11045;
    wire N__11044;
    wire N__11043;
    wire N__11042;
    wire N__11041;
    wire N__11040;
    wire N__11039;
    wire N__11038;
    wire N__11037;
    wire N__11036;
    wire N__11035;
    wire N__11034;
    wire N__11033;
    wire N__11032;
    wire N__11031;
    wire N__11030;
    wire N__11029;
    wire N__11026;
    wire N__11025;
    wire N__11024;
    wire N__11023;
    wire N__11022;
    wire N__11021;
    wire N__11020;
    wire N__11019;
    wire N__11018;
    wire N__11017;
    wire N__11016;
    wire N__11015;
    wire N__11014;
    wire N__11013;
    wire N__11012;
    wire N__11011;
    wire N__11010;
    wire N__11009;
    wire N__11008;
    wire N__11007;
    wire N__11006;
    wire N__11005;
    wire N__11004;
    wire N__11003;
    wire N__11002;
    wire N__11001;
    wire N__10892;
    wire N__10889;
    wire N__10888;
    wire N__10887;
    wire N__10884;
    wire N__10881;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10870;
    wire N__10867;
    wire N__10864;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10830;
    wire N__10827;
    wire N__10824;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10808;
    wire N__10807;
    wire N__10804;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10789;
    wire N__10788;
    wire N__10783;
    wire N__10780;
    wire N__10775;
    wire N__10772;
    wire N__10771;
    wire N__10768;
    wire N__10765;
    wire N__10764;
    wire N__10763;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10747;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10727;
    wire N__10724;
    wire N__10719;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10707;
    wire N__10704;
    wire N__10699;
    wire N__10694;
    wire N__10691;
    wire N__10690;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10679;
    wire N__10674;
    wire N__10671;
    wire N__10668;
    wire N__10667;
    wire N__10666;
    wire N__10663;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10644;
    wire N__10641;
    wire N__10638;
    wire N__10635;
    wire N__10632;
    wire N__10629;
    wire N__10626;
    wire N__10623;
    wire N__10616;
    wire N__10613;
    wire N__10612;
    wire N__10611;
    wire N__10610;
    wire N__10609;
    wire N__10606;
    wire N__10605;
    wire N__10602;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10598;
    wire N__10597;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10587;
    wire N__10586;
    wire N__10583;
    wire N__10576;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10562;
    wire N__10561;
    wire N__10560;
    wire N__10555;
    wire N__10554;
    wire N__10553;
    wire N__10552;
    wire N__10551;
    wire N__10550;
    wire N__10549;
    wire N__10548;
    wire N__10543;
    wire N__10542;
    wire N__10541;
    wire N__10534;
    wire N__10531;
    wire N__10528;
    wire N__10525;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10503;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10472;
    wire N__10469;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10422;
    wire N__10421;
    wire N__10416;
    wire N__10415;
    wire N__10412;
    wire N__10411;
    wire N__10408;
    wire N__10405;
    wire N__10400;
    wire N__10397;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10354;
    wire N__10353;
    wire N__10352;
    wire N__10349;
    wire N__10344;
    wire N__10341;
    wire N__10338;
    wire N__10333;
    wire N__10330;
    wire N__10327;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10313;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10305;
    wire N__10304;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10288;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10239;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10205;
    wire N__10202;
    wire N__10201;
    wire N__10198;
    wire N__10195;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10099;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10082;
    wire N__10081;
    wire N__10080;
    wire N__10079;
    wire N__10078;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10043;
    wire N__10042;
    wire N__10041;
    wire N__10040;
    wire N__10039;
    wire N__10038;
    wire N__10037;
    wire N__10034;
    wire N__10033;
    wire N__10032;
    wire N__10031;
    wire N__10030;
    wire N__10023;
    wire N__10016;
    wire N__10013;
    wire N__10006;
    wire N__10003;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9983;
    wire N__9980;
    wire N__9979;
    wire N__9978;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9967;
    wire N__9964;
    wire N__9963;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9942;
    wire N__9937;
    wire N__9934;
    wire N__9931;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9901;
    wire N__9898;
    wire N__9895;
    wire N__9892;
    wire N__9889;
    wire N__9884;
    wire N__9883;
    wire N__9882;
    wire N__9879;
    wire N__9878;
    wire N__9873;
    wire N__9870;
    wire N__9867;
    wire N__9864;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9844;
    wire N__9841;
    wire N__9838;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9805;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9788;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9766;
    wire N__9765;
    wire N__9762;
    wire N__9757;
    wire N__9756;
    wire N__9755;
    wire N__9754;
    wire N__9753;
    wire N__9752;
    wire N__9747;
    wire N__9744;
    wire N__9735;
    wire N__9730;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9710;
    wire N__9707;
    wire N__9706;
    wire N__9703;
    wire N__9702;
    wire N__9699;
    wire N__9696;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9684;
    wire N__9683;
    wire N__9682;
    wire N__9681;
    wire N__9680;
    wire N__9679;
    wire N__9678;
    wire N__9675;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9663;
    wire N__9654;
    wire N__9647;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9629;
    wire N__9626;
    wire N__9625;
    wire N__9624;
    wire N__9623;
    wire N__9622;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9614;
    wire N__9613;
    wire N__9612;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9585;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9571;
    wire N__9568;
    wire N__9563;
    wire N__9558;
    wire N__9555;
    wire N__9552;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9536;
    wire N__9533;
    wire N__9532;
    wire N__9529;
    wire N__9528;
    wire N__9525;
    wire N__9522;
    wire N__9521;
    wire N__9520;
    wire N__9519;
    wire N__9516;
    wire N__9515;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9503;
    wire N__9502;
    wire N__9499;
    wire N__9494;
    wire N__9491;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9475;
    wire N__9470;
    wire N__9467;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9451;
    wire N__9448;
    wire N__9445;
    wire N__9442;
    wire N__9439;
    wire N__9436;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9391;
    wire N__9390;
    wire N__9389;
    wire N__9388;
    wire N__9387;
    wire N__9386;
    wire N__9379;
    wire N__9376;
    wire N__9369;
    wire N__9368;
    wire N__9365;
    wire N__9360;
    wire N__9359;
    wire N__9356;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9329;
    wire N__9328;
    wire N__9327;
    wire N__9326;
    wire N__9325;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9297;
    wire N__9292;
    wire N__9289;
    wire N__9286;
    wire N__9283;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9250;
    wire N__9249;
    wire N__9246;
    wire N__9245;
    wire N__9244;
    wire N__9241;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9216;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9190;
    wire N__9179;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9165;
    wire N__9164;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9149;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9124;
    wire N__9123;
    wire N__9122;
    wire N__9121;
    wire N__9120;
    wire N__9119;
    wire N__9116;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9108;
    wire N__9105;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9085;
    wire N__9084;
    wire N__9083;
    wire N__9082;
    wire N__9081;
    wire N__9080;
    wire N__9079;
    wire N__9076;
    wire N__9075;
    wire N__9074;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9044;
    wire N__9039;
    wire N__9036;
    wire N__9035;
    wire N__9032;
    wire N__9027;
    wire N__9024;
    wire N__9021;
    wire N__9018;
    wire N__9015;
    wire N__9008;
    wire N__9003;
    wire N__9002;
    wire N__8999;
    wire N__8998;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8986;
    wire N__8983;
    wire N__8976;
    wire N__8969;
    wire N__8966;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8914;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8904;
    wire N__8897;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8889;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8864;
    wire N__8861;
    wire N__8860;
    wire N__8859;
    wire N__8858;
    wire N__8855;
    wire N__8850;
    wire N__8847;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8812;
    wire N__8811;
    wire N__8810;
    wire N__8805;
    wire N__8802;
    wire N__8799;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8668;
    wire N__8667;
    wire N__8666;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8640;
    wire N__8637;
    wire N__8634;
    wire N__8631;
    wire N__8628;
    wire N__8623;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8584;
    wire N__8581;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8379;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8367;
    wire N__8360;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8334;
    wire N__8333;
    wire N__8332;
    wire N__8331;
    wire N__8330;
    wire N__8329;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8300;
    wire N__8299;
    wire N__8294;
    wire N__8289;
    wire N__8286;
    wire N__8279;
    wire N__8276;
    wire N__8275;
    wire N__8274;
    wire N__8271;
    wire N__8266;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8251;
    wire N__8250;
    wire N__8245;
    wire N__8242;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8224;
    wire N__8221;
    wire N__8218;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8192;
    wire N__8189;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8165;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8126;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8116;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8066;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8029;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8014;
    wire N__8011;
    wire N__8008;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7909;
    wire N__7908;
    wire N__7907;
    wire N__7902;
    wire N__7897;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7865;
    wire N__7864;
    wire N__7861;
    wire N__7860;
    wire N__7855;
    wire N__7852;
    wire N__7847;
    wire N__7846;
    wire N__7845;
    wire N__7844;
    wire N__7841;
    wire N__7836;
    wire N__7833;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7819;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7798;
    wire N__7795;
    wire N__7792;
    wire N__7789;
    wire N__7784;
    wire N__7781;
    wire N__7778;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7753;
    wire N__7752;
    wire N__7751;
    wire N__7748;
    wire N__7745;
    wire N__7740;
    wire N__7733;
    wire N__7730;
    wire N__7727;
    wire N__7726;
    wire N__7721;
    wire N__7718;
    wire N__7715;
    wire N__7714;
    wire N__7711;
    wire N__7710;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7683;
    wire N__7678;
    wire N__7673;
    wire N__7670;
    wire N__7669;
    wire N__7666;
    wire N__7665;
    wire N__7662;
    wire N__7657;
    wire N__7652;
    wire N__7651;
    wire N__7648;
    wire N__7647;
    wire N__7644;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7632;
    wire N__7629;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7602;
    wire N__7601;
    wire N__7598;
    wire N__7593;
    wire N__7590;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7537;
    wire N__7532;
    wire N__7529;
    wire N__7528;
    wire N__7525;
    wire N__7522;
    wire N__7519;
    wire N__7516;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7502;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7474;
    wire N__7471;
    wire N__7468;
    wire N__7465;
    wire N__7462;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7424;
    wire N__7421;
    wire N__7418;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7408;
    wire N__7407;
    wire N__7406;
    wire N__7401;
    wire N__7398;
    wire N__7395;
    wire N__7388;
    wire N__7385;
    wire N__7382;
    wire N__7379;
    wire N__7376;
    wire N__7375;
    wire N__7374;
    wire N__7373;
    wire N__7370;
    wire N__7369;
    wire N__7368;
    wire N__7367;
    wire N__7364;
    wire N__7363;
    wire N__7362;
    wire N__7359;
    wire N__7356;
    wire N__7353;
    wire N__7350;
    wire N__7347;
    wire N__7344;
    wire N__7339;
    wire N__7338;
    wire N__7335;
    wire N__7334;
    wire N__7331;
    wire N__7328;
    wire N__7321;
    wire N__7320;
    wire N__7319;
    wire N__7318;
    wire N__7317;
    wire N__7316;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7302;
    wire N__7297;
    wire N__7296;
    wire N__7295;
    wire N__7294;
    wire N__7291;
    wire N__7288;
    wire N__7281;
    wire N__7278;
    wire N__7275;
    wire N__7268;
    wire N__7265;
    wire N__7258;
    wire N__7241;
    wire N__7240;
    wire N__7237;
    wire N__7236;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7226;
    wire N__7223;
    wire N__7222;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7214;
    wire N__7213;
    wire N__7212;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire N__7202;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7181;
    wire N__7178;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7148;
    wire N__7147;
    wire N__7146;
    wire N__7145;
    wire N__7144;
    wire N__7141;
    wire N__7140;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7132;
    wire N__7131;
    wire N__7128;
    wire N__7125;
    wire N__7122;
    wire N__7119;
    wire N__7116;
    wire N__7113;
    wire N__7112;
    wire N__7111;
    wire N__7110;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7098;
    wire N__7087;
    wire N__7080;
    wire N__7077;
    wire N__7064;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7051;
    wire N__7048;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7030;
    wire N__7027;
    wire N__7024;
    wire N__7023;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7001;
    wire N__6998;
    wire N__6997;
    wire N__6996;
    wire N__6995;
    wire N__6994;
    wire N__6991;
    wire N__6988;
    wire N__6985;
    wire N__6982;
    wire N__6979;
    wire N__6978;
    wire N__6977;
    wire N__6974;
    wire N__6971;
    wire N__6968;
    wire N__6965;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6949;
    wire N__6942;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6921;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6884;
    wire N__6881;
    wire N__6876;
    wire N__6873;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6820;
    wire N__6819;
    wire N__6818;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6800;
    wire N__6797;
    wire N__6796;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6775;
    wire N__6772;
    wire N__6769;
    wire N__6768;
    wire N__6767;
    wire N__6762;
    wire N__6761;
    wire N__6760;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6750;
    wire N__6745;
    wire N__6742;
    wire N__6731;
    wire N__6728;
    wire N__6727;
    wire N__6724;
    wire N__6723;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6697;
    wire N__6696;
    wire N__6693;
    wire N__6690;
    wire N__6687;
    wire N__6680;
    wire N__6677;
    wire N__6676;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6643;
    wire N__6642;
    wire N__6639;
    wire N__6636;
    wire N__6635;
    wire N__6634;
    wire N__6633;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6623;
    wire N__6622;
    wire N__6617;
    wire N__6614;
    wire N__6607;
    wire N__6602;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6584;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6563;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6551;
    wire N__6548;
    wire N__6547;
    wire N__6546;
    wire N__6543;
    wire N__6542;
    wire N__6541;
    wire N__6540;
    wire N__6539;
    wire N__6538;
    wire N__6537;
    wire N__6536;
    wire N__6535;
    wire N__6534;
    wire N__6533;
    wire N__6532;
    wire N__6531;
    wire N__6528;
    wire N__6527;
    wire N__6526;
    wire N__6525;
    wire N__6524;
    wire N__6523;
    wire N__6520;
    wire N__6519;
    wire N__6518;
    wire N__6517;
    wire N__6516;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6498;
    wire N__6495;
    wire N__6488;
    wire N__6479;
    wire N__6478;
    wire N__6477;
    wire N__6476;
    wire N__6471;
    wire N__6464;
    wire N__6461;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6439;
    wire N__6430;
    wire N__6429;
    wire N__6424;
    wire N__6421;
    wire N__6416;
    wire N__6411;
    wire N__6402;
    wire N__6399;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6377;
    wire N__6374;
    wire N__6371;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6302;
    wire N__6299;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6268;
    wire N__6265;
    wire N__6262;
    wire N__6257;
    wire N__6254;
    wire N__6251;
    wire N__6250;
    wire N__6249;
    wire N__6246;
    wire N__6243;
    wire N__6240;
    wire N__6237;
    wire N__6230;
    wire N__6227;
    wire N__6224;
    wire N__6221;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6209;
    wire N__6206;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6195;
    wire N__6194;
    wire N__6193;
    wire N__6192;
    wire N__6191;
    wire N__6190;
    wire N__6187;
    wire N__6184;
    wire N__6177;
    wire N__6170;
    wire N__6161;
    wire N__6158;
    wire N__6157;
    wire N__6154;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6133;
    wire N__6132;
    wire N__6131;
    wire N__6130;
    wire N__6129;
    wire N__6128;
    wire N__6127;
    wire N__6126;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6116;
    wire N__6111;
    wire N__6106;
    wire N__6099;
    wire N__6086;
    wire N__6085;
    wire N__6084;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6068;
    wire N__6065;
    wire N__6062;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6050;
    wire N__6047;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6035;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6008;
    wire N__6005;
    wire N__6002;
    wire N__5999;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5975;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5940;
    wire N__5935;
    wire N__5932;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5869;
    wire N__5866;
    wire N__5863;
    wire N__5858;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5846;
    wire N__5845;
    wire N__5842;
    wire N__5839;
    wire N__5836;
    wire N__5831;
    wire N__5830;
    wire N__5827;
    wire N__5824;
    wire N__5819;
    wire N__5816;
    wire N__5815;
    wire N__5812;
    wire N__5807;
    wire N__5806;
    wire N__5805;
    wire N__5802;
    wire N__5801;
    wire N__5800;
    wire N__5799;
    wire N__5798;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5788;
    wire N__5785;
    wire N__5782;
    wire N__5777;
    wire N__5774;
    wire N__5759;
    wire N__5756;
    wire N__5753;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5745;
    wire N__5744;
    wire N__5743;
    wire N__5738;
    wire N__5733;
    wire N__5730;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5707;
    wire N__5704;
    wire N__5703;
    wire N__5700;
    wire N__5699;
    wire N__5698;
    wire N__5697;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5679;
    wire N__5678;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5666;
    wire N__5661;
    wire N__5658;
    wire N__5653;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5628;
    wire N__5625;
    wire N__5622;
    wire N__5619;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5607;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5572;
    wire N__5571;
    wire N__5568;
    wire N__5563;
    wire N__5558;
    wire N__5555;
    wire N__5554;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5530;
    wire N__5527;
    wire N__5522;
    wire N__5519;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5500;
    wire N__5499;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5491;
    wire N__5482;
    wire N__5481;
    wire N__5480;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5459;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5407;
    wire N__5406;
    wire N__5405;
    wire N__5404;
    wire N__5403;
    wire N__5402;
    wire N__5399;
    wire N__5392;
    wire N__5385;
    wire N__5382;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5342;
    wire N__5339;
    wire N__5336;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5290;
    wire N__5289;
    wire N__5288;
    wire N__5285;
    wire N__5278;
    wire N__5273;
    wire N__5270;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5189;
    wire N__5188;
    wire N__5183;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5101;
    wire N__5098;
    wire N__5095;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5069;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5026;
    wire N__5023;
    wire N__5022;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4930;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4903;
    wire N__4900;
    wire N__4897;
    wire N__4894;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4879;
    wire N__4876;
    wire N__4873;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4849;
    wire N__4846;
    wire N__4843;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4727;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4672;
    wire N__4671;
    wire N__4670;
    wire N__4669;
    wire N__4668;
    wire N__4667;
    wire N__4666;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4642;
    wire N__4639;
    wire N__4636;
    wire N__4631;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4619;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4604;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4592;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4580;
    wire N__4579;
    wire N__4576;
    wire N__4573;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire DBRn_c_i_0;
    wire CLK80_PLL_i_i;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_6_7_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire A_c_6;
    wire A_c_2;
    wire A_c_3;
    wire A_c_4;
    wire A_c_7;
    wire A_c_8;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0 ;
    wire DBRn_c;
    wire VBENn_c;
    wire A_c_18;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_a2_1_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_165_i_i_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire \U712_CHIP_RAM.N_90_i_cascade_ ;
    wire \U712_CHIP_RAM.N_298_cascade_ ;
    wire \U712_CHIP_RAM.N_300_cascade_ ;
    wire \U712_CHIP_RAM.N_310 ;
    wire \U712_CHIP_RAM.N_310_cascade_ ;
    wire \U712_CHIP_RAM.N_313 ;
    wire \U712_CHIP_RAM.N_389 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_5 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_4 ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_ ;
    wire bfn_8_12_0_;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ;
    wire DBR_SYNC_i_1;
    wire DBR_SYNCZ0Z_0;
    wire A_c_5;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ;
    wire A_c_16;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a3_0_a2_0 ;
    wire N_178_i;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ;
    wire N_176_i;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ;
    wire A_c_12;
    wire \U712_CHIP_RAM.SDRAM_COUNTER19 ;
    wire \U712_CHIP_RAM.N_464_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0 ;
    wire \U712_CHIP_RAM.N_390 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0 ;
    wire bfn_9_8_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_90_i ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire N_188_i;
    wire \U712_CHIP_RAM.N_302 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ;
    wire \U712_CHIP_RAM.N_455 ;
    wire \U712_CHIP_RAM.N_417_cascade_ ;
    wire RAMSPACEn_c;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH5lto7_0 ;
    wire \U712_CHIP_RAM.REFRESH5lt7 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.N_419 ;
    wire \U712_BYTE_ENABLE.N_326 ;
    wire \U712_BYTE_ENABLE.N_323 ;
    wire \U712_BYTE_ENABLE.N_324 ;
    wire A_c_17;
    wire \U712_CHIP_RAM.N_463_cascade_ ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.N_385_cascade_ ;
    wire \U712_CHIP_RAM.N_384 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_461 ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0_a2_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0_a2_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_1_cascade_ ;
    wire \U712_CHIP_RAM.N_533_cascade_ ;
    wire \U712_CHIP_RAM.N_370 ;
    wire \U712_CHIP_RAM.N_391_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0 ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_295_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_1 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_546 ;
    wire \U712_CHIP_RAM.N_464 ;
    wire \U712_CHIP_RAM.N_465 ;
    wire \U712_CHIP_RAM.N_465_cascade_ ;
    wire A_c_20;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0 ;
    wire \U712_CHIP_RAM.DBENn_8_0_0 ;
    wire DBDIR_c;
    wire CLK40_PLL_i_i;
    wire N_167_i;
    wire CONSTANT_ONE_NET;
    wire A_c_11;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ;
    wire LATCH_CLK_c;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_a2_0_1 ;
    wire \U712_CHIP_RAM.N_533 ;
    wire \U712_CHIP_RAM.N_296_cascade_ ;
    wire \U712_CHIP_RAM.N_550 ;
    wire \U712_CHIP_RAM.N_463 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ;
    wire \U712_CHIP_RAM.N_442_cascade_ ;
    wire \U712_CHIP_RAM.N_441 ;
    wire \U712_CHIP_RAM.CPU_TACK_8_iv_i_a2_1 ;
    wire \U712_CHIP_RAM.N_295 ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_551 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ;
    wire \U712_CHIP_RAM.N_458 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_0_0_0_a2_1 ;
    wire \U712_CHIP_RAM.N_428 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_0_cascade_ ;
    wire \U712_CHIP_RAM.N_300 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_438 ;
    wire \U712_CHIP_RAM.N_469 ;
    wire \U712_CHIP_RAM.N_438_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_a2_1 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_a2_2 ;
    wire DBENn_c;
    wire DMA_CYCLEm;
    wire \U712_CYCLE_TERM.N_321 ;
    wire TACK_EN;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire A_c_13;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ;
    wire A_c_15;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire A_c_9;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ;
    wire A_c_10;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.N_305_cascade_ ;
    wire A_c_14;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0 ;
    wire \U712_BYTE_ENABLE.N_325 ;
    wire N_186_i;
    wire CPU_TACKm;
    wire \U712_CYCLE_TERM.N_450_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_STATEZ1Z_2 ;
    wire CLK40_PLL_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire TACK_OUTn;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire REG_TACK;
    wire \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_5 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_6 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_4 ;
    wire \U712_REG_SM.N_320_cascade_ ;
    wire RESETn_c_i;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.un1_CMA25_0_i ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.N_346 ;
    wire \U712_CHIP_RAM.N_352 ;
    wire CMA_c_5;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ;
    wire N_169_i;
    wire REGSPACEn_c;
    wire \U712_REG_SM.N_397_cascade_ ;
    wire TSn_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_3 ;
    wire \U712_REG_SM.N_548 ;
    wire \U712_REG_SM.N_319_cascade_ ;
    wire \U712_REG_SM.REG_CYCLE_5_iv_0_0_cascade_ ;
    wire \U712_REG_SM.N_409 ;
    wire REG_CYCLEm;
    wire \U712_REG_SM.STATE_COUNTsr_0 ;
    wire \U712_REG_SM.N_328 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_REG_SM.N_412_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_3 ;
    wire \U712_REG_SM.N_360_cascade_ ;
    wire \U712_REG_SM.N_320 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire \U712_REG_SM.START_RSTZ0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_7 ;
    wire \U712_REG_SM.N_319 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire \U712_REG_SM.N_318_cascade_ ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire BLSn_c;
    wire \U712_REG_SM.REGENn_e_1 ;
    wire N_326_i;
    wire N_325_i;
    wire N_323_i;
    wire A_c_1;
    wire SIZ_c_1;
    wire A_c_0;
    wire SIZ_c_0;
    wire N_324_i;
    wire WEn_c;
    wire \U712_CHIP_RAM.N_305 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.un1_CMA25_0_i_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire \U712_CHIP_RAM.CMA_5_i_0_9 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire CPU_CYCLEm;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_8 ;
    wire \U712_REG_SM.N_400 ;
    wire UDSn_c;
    wire \U712_REG_SM.WRITE_CYCLEZ0 ;
    wire PRnW_c;
    wire \U712_REG_SM.N_398 ;
    wire LDSn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire DRA_c_5;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire DRA_c_1;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_2 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_152 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire ASn_c;
    wire \U712_REG_SM.N_152_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire DRA_c_7;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_2;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_9;
    wire AGNUS_REV_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire RESETn_c;
    wire RAS1n_c;
    wire RAS0n_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire CLK80_PLL;
    wire RnW_c;
    wire DMA_WRITE_CYCLE;
    wire CASLn_c;
    wire CASUn_c;
    wire N_362;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__4445),
            .RESETB(N__6377),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__13257),
            .DIN(N__13256),
            .DOUT(N__13255),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__13257),
            .PADOUT(N__13256),
            .PADIN(N__13255),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7040),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__13248),
            .DIN(N__13247),
            .DOUT(N__13246),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__13248),
            .PADOUT(N__13247),
            .PADIN(N__13246),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__13239),
            .DIN(N__13238),
            .DOUT(N__13237),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__13239),
            .PADOUT(N__13238),
            .PADIN(N__13237),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10454),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__13230),
            .DIN(N__13229),
            .DOUT(N__13228),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__13230),
            .PADOUT(N__13229),
            .PADIN(N__13228),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12374),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__13221),
            .DIN(N__13220),
            .DOUT(N__13219),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__13221),
            .PADOUT(N__13220),
            .PADIN(N__13219),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__13212),
            .DIN(N__13211),
            .DOUT(N__13210),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__13212),
            .PADOUT(N__13211),
            .PADIN(N__13210),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__13203),
            .DIN(N__13202),
            .DOUT(N__13201),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__13203),
            .PADOUT(N__13202),
            .PADIN(N__13201),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__13194),
            .DIN(N__13193),
            .DOUT(N__13192),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__13194),
            .PADOUT(N__13193),
            .PADIN(N__13192),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__13185),
            .DIN(N__13184),
            .DOUT(N__13183),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__13185),
            .PADOUT(N__13184),
            .PADIN(N__13183),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__13176),
            .DIN(N__13175),
            .DOUT(N__13174),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__13176),
            .PADOUT(N__13175),
            .PADIN(N__13174),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__13167),
            .DIN(N__13166),
            .DOUT(N__13165),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__13167),
            .PADOUT(N__13166),
            .PADIN(N__13165),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__13158),
            .DIN(N__13157),
            .DOUT(N__13156),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__13158),
            .PADOUT(N__13157),
            .PADIN(N__13156),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8420),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__13149),
            .DIN(N__13148),
            .DOUT(N__13147),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__13149),
            .PADOUT(N__13148),
            .PADIN(N__13147),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8786),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__13140),
            .DIN(N__13139),
            .DOUT(N__13138),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__13140),
            .PADOUT(N__13139),
            .PADIN(N__13138),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__13131),
            .DIN(N__13130),
            .DOUT(N__13129),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__13131),
            .PADOUT(N__13130),
            .PADIN(N__13129),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__13122),
            .DIN(N__13121),
            .DOUT(N__13120),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__13122),
            .PADOUT(N__13121),
            .PADIN(N__13120),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__13113),
            .DIN(N__13112),
            .DOUT(N__13111),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__13113),
            .PADOUT(N__13112),
            .PADIN(N__13111),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4691),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__13104),
            .DIN(N__13103),
            .DOUT(N__13102),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__13104),
            .PADOUT(N__13103),
            .PADIN(N__13102),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__13095),
            .DIN(N__13094),
            .DOUT(N__13093),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__13095),
            .PADOUT(N__13094),
            .PADIN(N__13093),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__13086),
            .DIN(N__13085),
            .DOUT(N__13084),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__13086),
            .PADOUT(N__13085),
            .PADIN(N__13084),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8549),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__13077),
            .DIN(N__13076),
            .DOUT(N__13075),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__13077),
            .PADOUT(N__13076),
            .PADIN(N__13075),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__13068),
            .DIN(N__13067),
            .DOUT(N__13066),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__13068),
            .PADOUT(N__13067),
            .PADIN(N__13066),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12140),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__13059),
            .DIN(N__13058),
            .DOUT(N__13057),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__13059),
            .PADOUT(N__13058),
            .PADIN(N__13057),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__13050),
            .DIN(N__13049),
            .DOUT(N__13048),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__13050),
            .PADOUT(N__13049),
            .PADIN(N__13048),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9782),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__13041),
            .DIN(N__13040),
            .DOUT(N__13039),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__13041),
            .PADOUT(N__13040),
            .PADIN(N__13039),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6921),
            .DIN0(),
            .DOUT0(N__7647),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__13032),
            .DIN(N__13031),
            .DOUT(N__13030),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__13032),
            .PADOUT(N__13031),
            .PADIN(N__13030),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__13023),
            .DIN(N__13022),
            .DOUT(N__13021),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__13023),
            .PADOUT(N__13022),
            .PADIN(N__13021),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__13014),
            .DIN(N__13013),
            .DOUT(N__13012),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__13014),
            .PADOUT(N__13013),
            .PADIN(N__13012),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__13005),
            .DIN(N__13004),
            .DOUT(N__13003),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__13005),
            .PADOUT(N__13004),
            .PADIN(N__13003),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__12996),
            .DIN(N__12995),
            .DOUT(N__12994),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__12996),
            .PADOUT(N__12995),
            .PADIN(N__12994),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__12987),
            .DIN(N__12986),
            .DOUT(N__12985),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__12987),
            .PADOUT(N__12986),
            .PADIN(N__12985),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5924),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__12978),
            .DIN(N__12977),
            .DOUT(N__12976),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__12978),
            .PADOUT(N__12977),
            .PADIN(N__12976),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__12969),
            .DIN(N__12968),
            .DOUT(N__12967),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__12969),
            .PADOUT(N__12968),
            .PADIN(N__12967),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__12960),
            .DIN(N__12959),
            .DOUT(N__12958),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__12960),
            .PADOUT(N__12959),
            .PADIN(N__12958),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__12951),
            .DIN(N__12950),
            .DOUT(N__12949),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__12951),
            .PADOUT(N__12950),
            .PADIN(N__12949),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__12942),
            .DIN(N__12941),
            .DOUT(N__12940),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__12942),
            .PADOUT(N__12941),
            .PADIN(N__12940),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__12933),
            .DIN(N__12932),
            .DOUT(N__12931),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__12933),
            .PADOUT(N__12932),
            .PADIN(N__12931),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10388),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__12924),
            .DIN(N__12923),
            .DOUT(N__12922),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__12924),
            .PADOUT(N__12923),
            .PADIN(N__12922),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__12915),
            .DIN(N__12914),
            .DOUT(N__12913),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__12915),
            .PADOUT(N__12914),
            .PADIN(N__12913),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__12906),
            .DIN(N__12905),
            .DOUT(N__12904),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__12906),
            .PADOUT(N__12905),
            .PADIN(N__12904),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12218),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_0_iopad (
            .OE(N__12897),
            .DIN(N__12896),
            .DOUT(N__12895),
            .PACKAGEPIN(DA[0]));
    defparam DA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_0_preio (
            .PADOEN(N__12897),
            .PADOUT(N__12896),
            .PADIN(N__12895),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7532),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__12888),
            .DIN(N__12887),
            .DOUT(N__12886),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__12888),
            .PADOUT(N__12887),
            .PADIN(N__12886),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__12879),
            .DIN(N__12878),
            .DOUT(N__12877),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__12879),
            .PADOUT(N__12878),
            .PADIN(N__12877),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8531),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__12870),
            .DIN(N__12869),
            .DOUT(N__12868),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__12870),
            .PADOUT(N__12869),
            .PADIN(N__12868),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8447),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__12861),
            .DIN(N__12860),
            .DOUT(N__12859),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__12861),
            .PADOUT(N__12860),
            .PADIN(N__12859),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8840),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__12852),
            .DIN(N__12851),
            .DOUT(N__12850),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__12852),
            .PADOUT(N__12851),
            .PADIN(N__12850),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__12843),
            .DIN(N__12842),
            .DOUT(N__12841),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__12843),
            .PADOUT(N__12842),
            .PADIN(N__12841),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7769),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__12834),
            .DIN(N__12833),
            .DOUT(N__12832),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__12834),
            .PADOUT(N__12833),
            .PADIN(N__12832),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6928),
            .DIN0(),
            .DOUT0(N__7651),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__12825),
            .DIN(N__12824),
            .DOUT(N__12823),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__12825),
            .PADOUT(N__12824),
            .PADIN(N__12823),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9413),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__12816),
            .DIN(N__12815),
            .DOUT(N__12814),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__12816),
            .PADOUT(N__12815),
            .PADIN(N__12814),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6002),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__12807),
            .DIN(N__12806),
            .DOUT(N__12805),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__12807),
            .PADOUT(N__12806),
            .PADIN(N__12805),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4952),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__12798),
            .DIN(N__12797),
            .DOUT(N__12796),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__12798),
            .PADOUT(N__12797),
            .PADIN(N__12796),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__12789),
            .DIN(N__12788),
            .DOUT(N__12787),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__12789),
            .PADOUT(N__12788),
            .PADIN(N__12787),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_2_iopad (
            .OE(N__12780),
            .DIN(N__12779),
            .DOUT(N__12778),
            .PACKAGEPIN(DA[2]));
    defparam DA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_2_preio (
            .PADOEN(N__12780),
            .PADOUT(N__12779),
            .PADIN(N__12778),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6347),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__12771),
            .DIN(N__12770),
            .DOUT(N__12769),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__12771),
            .PADOUT(N__12770),
            .PADIN(N__12769),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__12762),
            .DIN(N__12761),
            .DOUT(N__12760),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__12762),
            .PADOUT(N__12761),
            .PADIN(N__12760),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__12753),
            .DIN(N__12752),
            .DOUT(N__12751),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__12753),
            .PADOUT(N__12752),
            .PADIN(N__12751),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7934),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__12744),
            .DIN(N__12743),
            .DOUT(N__12742),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__12744),
            .PADOUT(N__12743),
            .PADIN(N__12742),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9800),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__12735),
            .DIN(N__12734),
            .DOUT(N__12733),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__12735),
            .PADOUT(N__12734),
            .PADIN(N__12733),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__12726),
            .DIN(N__12725),
            .DOUT(N__12724),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__12726),
            .PADOUT(N__12725),
            .PADIN(N__12724),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5177),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__12717),
            .DIN(N__12716),
            .DOUT(N__12715),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__12717),
            .PADOUT(N__12716),
            .PADIN(N__12715),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6929),
            .DIN0(),
            .DOUT0(N__7652),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__12708),
            .DIN(N__12707),
            .DOUT(N__12706),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__12708),
            .PADOUT(N__12707),
            .PADIN(N__12706),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6860),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__12699),
            .DIN(N__12698),
            .DOUT(N__12697),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__12699),
            .PADOUT(N__12698),
            .PADIN(N__12697),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__12690),
            .DIN(N__12689),
            .DOUT(N__12688),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__12690),
            .PADOUT(N__12689),
            .PADIN(N__12688),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__12681),
            .DIN(N__12680),
            .DOUT(N__12679),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__12681),
            .PADOUT(N__12680),
            .PADIN(N__12679),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8480),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__12672),
            .DIN(N__12671),
            .DOUT(N__12670),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__12672),
            .PADOUT(N__12671),
            .PADIN(N__12670),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__12663),
            .DIN(N__12662),
            .DOUT(N__12661),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__12663),
            .PADOUT(N__12662),
            .PADIN(N__12661),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_1_iopad (
            .OE(N__12654),
            .DIN(N__12653),
            .DOUT(N__12652),
            .PACKAGEPIN(DA[1]));
    defparam DA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_1_preio (
            .PADOEN(N__12654),
            .PADOUT(N__12653),
            .PADIN(N__12652),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7493),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__12645),
            .DIN(N__12644),
            .DOUT(N__12643),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__12645),
            .PADOUT(N__12644),
            .PADIN(N__12643),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__12636),
            .DIN(N__12635),
            .DOUT(N__12634),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__12636),
            .PADOUT(N__12635),
            .PADIN(N__12634),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__12627),
            .DIN(N__12626),
            .DOUT(N__12625),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__12627),
            .PADOUT(N__12626),
            .PADIN(N__12625),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8177),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__12618),
            .DIN(N__12617),
            .DOUT(N__12616),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__12618),
            .PADOUT(N__12617),
            .PADIN(N__12616),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9914),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__12609),
            .DIN(N__12608),
            .DOUT(N__12607),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__12609),
            .PADOUT(N__12608),
            .PADIN(N__12607),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9431),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__12600),
            .DIN(N__12599),
            .DOUT(N__12598),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__12600),
            .PADOUT(N__12599),
            .PADIN(N__12598),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5885),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__12591),
            .DIN(N__12590),
            .DOUT(N__12589),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__12591),
            .PADOUT(N__12590),
            .PADIN(N__12589),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__12582),
            .DIN(N__12581),
            .DOUT(N__12580),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__12582),
            .PADOUT(N__12581),
            .PADIN(N__12580),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__12573),
            .DIN(N__12572),
            .DOUT(N__12571),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__12573),
            .PADOUT(N__12572),
            .PADIN(N__12571),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8507),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__12564),
            .DIN(N__12563),
            .DOUT(N__12562),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__12564),
            .PADOUT(N__12563),
            .PADIN(N__12562),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__12555),
            .DIN(N__12554),
            .DOUT(N__12553),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__12555),
            .PADOUT(N__12554),
            .PADIN(N__12553),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__12546),
            .DIN(N__12545),
            .DOUT(N__12544),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__12546),
            .PADOUT(N__12545),
            .PADIN(N__12544),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6287),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__12537),
            .DIN(N__12536),
            .DOUT(N__12535),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__12537),
            .PADOUT(N__12536),
            .PADIN(N__12535),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9827),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__12528),
            .DIN(N__12527),
            .DOUT(N__12526),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__12528),
            .PADOUT(N__12527),
            .PADIN(N__12526),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5975),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PRnW_obuf_iopad (
            .OE(N__12519),
            .DIN(N__12518),
            .DOUT(N__12517),
            .PACKAGEPIN(PRnW));
    defparam PRnW_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PRnW_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PRnW_obuf_preio (
            .PADOEN(N__12519),
            .PADOUT(N__12518),
            .PADIN(N__12517),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9857),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__12510),
            .DIN(N__12509),
            .DOUT(N__12508),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__12510),
            .PADOUT(N__12509),
            .PADIN(N__12508),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__12501),
            .DIN(N__12500),
            .DOUT(N__12499),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__12501),
            .PADOUT(N__12500),
            .PADIN(N__12499),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5974),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__12492),
            .DIN(N__12491),
            .DOUT(N__12490),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__12492),
            .PADOUT(N__12491),
            .PADIN(N__12490),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4484),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__12483),
            .DIN(N__12482),
            .DOUT(N__12481),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__12483),
            .PADOUT(N__12482),
            .PADIN(N__12481),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9272),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__12474),
            .DIN(N__12473),
            .DOUT(N__12472),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__12474),
            .PADOUT(N__12473),
            .PADIN(N__12472),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__12465),
            .DIN(N__12464),
            .DOUT(N__12463),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__12465),
            .PADOUT(N__12464),
            .PADIN(N__12463),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__12456),
            .DIN(N__12455),
            .DOUT(N__12454),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__12456),
            .PADOUT(N__12455),
            .PADIN(N__12454),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BLSn_obuf_iopad (
            .OE(N__12447),
            .DIN(N__12446),
            .DOUT(N__12445),
            .PACKAGEPIN(BLSn));
    defparam BLSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BLSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BLSn_obuf_preio (
            .PADOEN(N__12447),
            .PADOUT(N__12446),
            .PADIN(N__12445),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8830),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__12438),
            .DIN(N__12437),
            .DOUT(N__12436),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__12438),
            .PADOUT(N__12437),
            .PADIN(N__12436),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__12429),
            .DIN(N__12428),
            .DOUT(N__12427),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__12429),
            .PADOUT(N__12428),
            .PADIN(N__12427),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5949),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__12420),
            .DIN(N__12419),
            .DOUT(N__12418),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__12420),
            .PADOUT(N__12419),
            .PADIN(N__12418),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8111),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__12411),
            .DIN(N__12410),
            .DOUT(N__12409),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__12411),
            .PADOUT(N__12410),
            .PADIN(N__12409),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5372),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__12402),
            .DIN(N__12401),
            .DOUT(N__12400),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__12402),
            .PADOUT(N__12401),
            .PADIN(N__12400),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8750),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__12393),
            .DIN(N__12392),
            .DOUT(N__12391),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__12393),
            .PADOUT(N__12392),
            .PADIN(N__12391),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__3032 (
            .O(N__12374),
            .I(N__12371));
    LocalMux I__3031 (
            .O(N__12371),
            .I(N__12368));
    Span4Mux_s3_h I__3030 (
            .O(N__12368),
            .I(N__12365));
    Span4Mux_v I__3029 (
            .O(N__12365),
            .I(N__12362));
    Odrv4 I__3028 (
            .O(N__12362),
            .I(N_362));
    CascadeMux I__3027 (
            .O(N__12359),
            .I(N__12354));
    InMux I__3026 (
            .O(N__12358),
            .I(N__12351));
    InMux I__3025 (
            .O(N__12357),
            .I(N__12345));
    InMux I__3024 (
            .O(N__12354),
            .I(N__12345));
    LocalMux I__3023 (
            .O(N__12351),
            .I(N__12342));
    InMux I__3022 (
            .O(N__12350),
            .I(N__12339));
    LocalMux I__3021 (
            .O(N__12345),
            .I(\U712_REG_SM.N_152 ));
    Odrv4 I__3020 (
            .O(N__12342),
            .I(\U712_REG_SM.N_152 ));
    LocalMux I__3019 (
            .O(N__12339),
            .I(\U712_REG_SM.N_152 ));
    CascadeMux I__3018 (
            .O(N__12332),
            .I(N__12326));
    InMux I__3017 (
            .O(N__12331),
            .I(N__12321));
    InMux I__3016 (
            .O(N__12330),
            .I(N__12315));
    CascadeMux I__3015 (
            .O(N__12329),
            .I(N__12311));
    InMux I__3014 (
            .O(N__12326),
            .I(N__12308));
    CascadeMux I__3013 (
            .O(N__12325),
            .I(N__12301));
    CascadeMux I__3012 (
            .O(N__12324),
            .I(N__12298));
    LocalMux I__3011 (
            .O(N__12321),
            .I(N__12294));
    InMux I__3010 (
            .O(N__12320),
            .I(N__12291));
    InMux I__3009 (
            .O(N__12319),
            .I(N__12286));
    InMux I__3008 (
            .O(N__12318),
            .I(N__12286));
    LocalMux I__3007 (
            .O(N__12315),
            .I(N__12283));
    InMux I__3006 (
            .O(N__12314),
            .I(N__12278));
    InMux I__3005 (
            .O(N__12311),
            .I(N__12278));
    LocalMux I__3004 (
            .O(N__12308),
            .I(N__12275));
    InMux I__3003 (
            .O(N__12307),
            .I(N__12268));
    InMux I__3002 (
            .O(N__12306),
            .I(N__12268));
    InMux I__3001 (
            .O(N__12305),
            .I(N__12268));
    InMux I__3000 (
            .O(N__12304),
            .I(N__12265));
    InMux I__2999 (
            .O(N__12301),
            .I(N__12262));
    InMux I__2998 (
            .O(N__12298),
            .I(N__12257));
    InMux I__2997 (
            .O(N__12297),
            .I(N__12257));
    Span4Mux_v I__2996 (
            .O(N__12294),
            .I(N__12252));
    LocalMux I__2995 (
            .O(N__12291),
            .I(N__12252));
    LocalMux I__2994 (
            .O(N__12286),
            .I(N__12249));
    Span4Mux_v I__2993 (
            .O(N__12283),
            .I(N__12246));
    LocalMux I__2992 (
            .O(N__12278),
            .I(N__12243));
    Span4Mux_h I__2991 (
            .O(N__12275),
            .I(N__12232));
    LocalMux I__2990 (
            .O(N__12268),
            .I(N__12232));
    LocalMux I__2989 (
            .O(N__12265),
            .I(N__12232));
    LocalMux I__2988 (
            .O(N__12262),
            .I(N__12232));
    LocalMux I__2987 (
            .O(N__12257),
            .I(N__12232));
    Span4Mux_h I__2986 (
            .O(N__12252),
            .I(N__12229));
    Odrv4 I__2985 (
            .O(N__12249),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2984 (
            .O(N__12246),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2983 (
            .O(N__12243),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2982 (
            .O(N__12232),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2981 (
            .O(N__12229),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    IoInMux I__2980 (
            .O(N__12218),
            .I(N__12215));
    LocalMux I__2979 (
            .O(N__12215),
            .I(N__12212));
    Span4Mux_s3_v I__2978 (
            .O(N__12212),
            .I(N__12209));
    Span4Mux_v I__2977 (
            .O(N__12209),
            .I(N__12206));
    Span4Mux_v I__2976 (
            .O(N__12206),
            .I(N__12203));
    Sp12to4 I__2975 (
            .O(N__12203),
            .I(N__12200));
    Odrv12 I__2974 (
            .O(N__12200),
            .I(ASn_c));
    CEMux I__2973 (
            .O(N__12197),
            .I(N__12194));
    LocalMux I__2972 (
            .O(N__12194),
            .I(N__12191));
    Span4Mux_h I__2971 (
            .O(N__12191),
            .I(N__12188));
    Odrv4 I__2970 (
            .O(N__12188),
            .I(\U712_REG_SM.N_152_0 ));
    InMux I__2969 (
            .O(N__12185),
            .I(N__12181));
    InMux I__2968 (
            .O(N__12184),
            .I(N__12178));
    LocalMux I__2967 (
            .O(N__12181),
            .I(N__12175));
    LocalMux I__2966 (
            .O(N__12178),
            .I(N__12170));
    Span4Mux_h I__2965 (
            .O(N__12175),
            .I(N__12167));
    CascadeMux I__2964 (
            .O(N__12174),
            .I(N__12163));
    InMux I__2963 (
            .O(N__12173),
            .I(N__12160));
    Span4Mux_h I__2962 (
            .O(N__12170),
            .I(N__12155));
    Span4Mux_h I__2961 (
            .O(N__12167),
            .I(N__12155));
    InMux I__2960 (
            .O(N__12166),
            .I(N__12152));
    InMux I__2959 (
            .O(N__12163),
            .I(N__12149));
    LocalMux I__2958 (
            .O(N__12160),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__2957 (
            .O(N__12155),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__2956 (
            .O(N__12152),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__2955 (
            .O(N__12149),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__2954 (
            .O(N__12140),
            .I(N__12137));
    LocalMux I__2953 (
            .O(N__12137),
            .I(N__12134));
    Span4Mux_s1_v I__2952 (
            .O(N__12134),
            .I(N__12131));
    Span4Mux_v I__2951 (
            .O(N__12131),
            .I(N__12128));
    Span4Mux_v I__2950 (
            .O(N__12128),
            .I(N__12125));
    Odrv4 I__2949 (
            .O(N__12125),
            .I(CRCSn_c));
    InMux I__2948 (
            .O(N__12122),
            .I(N__12116));
    InMux I__2947 (
            .O(N__12121),
            .I(N__12113));
    InMux I__2946 (
            .O(N__12120),
            .I(N__12110));
    InMux I__2945 (
            .O(N__12119),
            .I(N__12107));
    LocalMux I__2944 (
            .O(N__12116),
            .I(N__12102));
    LocalMux I__2943 (
            .O(N__12113),
            .I(N__12102));
    LocalMux I__2942 (
            .O(N__12110),
            .I(N__12099));
    LocalMux I__2941 (
            .O(N__12107),
            .I(N__12096));
    Span4Mux_v I__2940 (
            .O(N__12102),
            .I(N__12093));
    Span4Mux_h I__2939 (
            .O(N__12099),
            .I(N__12090));
    Span12Mux_v I__2938 (
            .O(N__12096),
            .I(N__12085));
    Sp12to4 I__2937 (
            .O(N__12093),
            .I(N__12085));
    Span4Mux_v I__2936 (
            .O(N__12090),
            .I(N__12082));
    Span12Mux_h I__2935 (
            .O(N__12085),
            .I(N__12079));
    Span4Mux_h I__2934 (
            .O(N__12082),
            .I(N__12076));
    Odrv12 I__2933 (
            .O(N__12079),
            .I(DRA_c_7));
    Odrv4 I__2932 (
            .O(N__12076),
            .I(DRA_c_7));
    InMux I__2931 (
            .O(N__12071),
            .I(N__12065));
    InMux I__2930 (
            .O(N__12070),
            .I(N__12062));
    InMux I__2929 (
            .O(N__12069),
            .I(N__12059));
    InMux I__2928 (
            .O(N__12068),
            .I(N__12056));
    LocalMux I__2927 (
            .O(N__12065),
            .I(N__12051));
    LocalMux I__2926 (
            .O(N__12062),
            .I(N__12051));
    LocalMux I__2925 (
            .O(N__12059),
            .I(N__12046));
    LocalMux I__2924 (
            .O(N__12056),
            .I(N__12046));
    Span4Mux_v I__2923 (
            .O(N__12051),
            .I(N__12043));
    Span4Mux_v I__2922 (
            .O(N__12046),
            .I(N__12040));
    Sp12to4 I__2921 (
            .O(N__12043),
            .I(N__12037));
    Sp12to4 I__2920 (
            .O(N__12040),
            .I(N__12034));
    Span12Mux_h I__2919 (
            .O(N__12037),
            .I(N__12031));
    Odrv12 I__2918 (
            .O(N__12034),
            .I(DRA_c_8));
    Odrv12 I__2917 (
            .O(N__12031),
            .I(DRA_c_8));
    InMux I__2916 (
            .O(N__12026),
            .I(N__12023));
    LocalMux I__2915 (
            .O(N__12023),
            .I(N__12020));
    Span4Mux_h I__2914 (
            .O(N__12020),
            .I(N__12017));
    Odrv4 I__2913 (
            .O(N__12017),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2912 (
            .O(N__12014),
            .I(N__12010));
    InMux I__2911 (
            .O(N__12013),
            .I(N__12007));
    LocalMux I__2910 (
            .O(N__12010),
            .I(N__12000));
    LocalMux I__2909 (
            .O(N__12007),
            .I(N__12000));
    InMux I__2908 (
            .O(N__12006),
            .I(N__11995));
    InMux I__2907 (
            .O(N__12005),
            .I(N__11995));
    Span4Mux_v I__2906 (
            .O(N__12000),
            .I(N__11992));
    LocalMux I__2905 (
            .O(N__11995),
            .I(N__11989));
    Sp12to4 I__2904 (
            .O(N__11992),
            .I(N__11986));
    Span12Mux_v I__2903 (
            .O(N__11989),
            .I(N__11983));
    Span12Mux_h I__2902 (
            .O(N__11986),
            .I(N__11980));
    Span12Mux_h I__2901 (
            .O(N__11983),
            .I(N__11977));
    Span12Mux_v I__2900 (
            .O(N__11980),
            .I(N__11974));
    Odrv12 I__2899 (
            .O(N__11977),
            .I(DRA_c_2));
    Odrv12 I__2898 (
            .O(N__11974),
            .I(DRA_c_2));
    InMux I__2897 (
            .O(N__11969),
            .I(N__11966));
    LocalMux I__2896 (
            .O(N__11966),
            .I(N__11961));
    InMux I__2895 (
            .O(N__11965),
            .I(N__11958));
    InMux I__2894 (
            .O(N__11964),
            .I(N__11955));
    Span4Mux_h I__2893 (
            .O(N__11961),
            .I(N__11948));
    LocalMux I__2892 (
            .O(N__11958),
            .I(N__11948));
    LocalMux I__2891 (
            .O(N__11955),
            .I(N__11948));
    Span4Mux_v I__2890 (
            .O(N__11948),
            .I(N__11944));
    InMux I__2889 (
            .O(N__11947),
            .I(N__11941));
    Span4Mux_v I__2888 (
            .O(N__11944),
            .I(N__11938));
    LocalMux I__2887 (
            .O(N__11941),
            .I(N__11935));
    Span4Mux_h I__2886 (
            .O(N__11938),
            .I(N__11932));
    Sp12to4 I__2885 (
            .O(N__11935),
            .I(N__11929));
    Sp12to4 I__2884 (
            .O(N__11932),
            .I(N__11924));
    Span12Mux_v I__2883 (
            .O(N__11929),
            .I(N__11924));
    Odrv12 I__2882 (
            .O(N__11924),
            .I(DRA_c_3));
    InMux I__2881 (
            .O(N__11921),
            .I(N__11918));
    LocalMux I__2880 (
            .O(N__11918),
            .I(N__11915));
    Span4Mux_h I__2879 (
            .O(N__11915),
            .I(N__11912));
    Span4Mux_h I__2878 (
            .O(N__11912),
            .I(N__11909));
    Odrv4 I__2877 (
            .O(N__11909),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    CascadeMux I__2876 (
            .O(N__11906),
            .I(N__11903));
    InMux I__2875 (
            .O(N__11903),
            .I(N__11899));
    InMux I__2874 (
            .O(N__11902),
            .I(N__11896));
    LocalMux I__2873 (
            .O(N__11899),
            .I(N__11892));
    LocalMux I__2872 (
            .O(N__11896),
            .I(N__11889));
    InMux I__2871 (
            .O(N__11895),
            .I(N__11886));
    Span4Mux_h I__2870 (
            .O(N__11892),
            .I(N__11880));
    Span4Mux_v I__2869 (
            .O(N__11889),
            .I(N__11880));
    LocalMux I__2868 (
            .O(N__11886),
            .I(N__11877));
    InMux I__2867 (
            .O(N__11885),
            .I(N__11874));
    Span4Mux_v I__2866 (
            .O(N__11880),
            .I(N__11871));
    Span4Mux_h I__2865 (
            .O(N__11877),
            .I(N__11868));
    LocalMux I__2864 (
            .O(N__11874),
            .I(N__11865));
    Sp12to4 I__2863 (
            .O(N__11871),
            .I(N__11862));
    Span4Mux_v I__2862 (
            .O(N__11868),
            .I(N__11859));
    Span4Mux_v I__2861 (
            .O(N__11865),
            .I(N__11856));
    Span12Mux_h I__2860 (
            .O(N__11862),
            .I(N__11853));
    Sp12to4 I__2859 (
            .O(N__11859),
            .I(N__11848));
    Sp12to4 I__2858 (
            .O(N__11856),
            .I(N__11848));
    Span12Mux_v I__2857 (
            .O(N__11853),
            .I(N__11845));
    Span12Mux_v I__2856 (
            .O(N__11848),
            .I(N__11842));
    Odrv12 I__2855 (
            .O(N__11845),
            .I(DRA_c_9));
    Odrv12 I__2854 (
            .O(N__11842),
            .I(DRA_c_9));
    CascadeMux I__2853 (
            .O(N__11837),
            .I(N__11832));
    CascadeMux I__2852 (
            .O(N__11836),
            .I(N__11824));
    InMux I__2851 (
            .O(N__11835),
            .I(N__11820));
    InMux I__2850 (
            .O(N__11832),
            .I(N__11816));
    InMux I__2849 (
            .O(N__11831),
            .I(N__11813));
    InMux I__2848 (
            .O(N__11830),
            .I(N__11808));
    InMux I__2847 (
            .O(N__11829),
            .I(N__11805));
    InMux I__2846 (
            .O(N__11828),
            .I(N__11802));
    InMux I__2845 (
            .O(N__11827),
            .I(N__11795));
    InMux I__2844 (
            .O(N__11824),
            .I(N__11790));
    InMux I__2843 (
            .O(N__11823),
            .I(N__11790));
    LocalMux I__2842 (
            .O(N__11820),
            .I(N__11787));
    InMux I__2841 (
            .O(N__11819),
            .I(N__11784));
    LocalMux I__2840 (
            .O(N__11816),
            .I(N__11781));
    LocalMux I__2839 (
            .O(N__11813),
            .I(N__11778));
    InMux I__2838 (
            .O(N__11812),
            .I(N__11775));
    InMux I__2837 (
            .O(N__11811),
            .I(N__11772));
    LocalMux I__2836 (
            .O(N__11808),
            .I(N__11765));
    LocalMux I__2835 (
            .O(N__11805),
            .I(N__11765));
    LocalMux I__2834 (
            .O(N__11802),
            .I(N__11765));
    InMux I__2833 (
            .O(N__11801),
            .I(N__11762));
    InMux I__2832 (
            .O(N__11800),
            .I(N__11754));
    InMux I__2831 (
            .O(N__11799),
            .I(N__11751));
    InMux I__2830 (
            .O(N__11798),
            .I(N__11748));
    LocalMux I__2829 (
            .O(N__11795),
            .I(N__11743));
    LocalMux I__2828 (
            .O(N__11790),
            .I(N__11743));
    Span4Mux_v I__2827 (
            .O(N__11787),
            .I(N__11738));
    LocalMux I__2826 (
            .O(N__11784),
            .I(N__11738));
    Span4Mux_h I__2825 (
            .O(N__11781),
            .I(N__11725));
    Span4Mux_v I__2824 (
            .O(N__11778),
            .I(N__11725));
    LocalMux I__2823 (
            .O(N__11775),
            .I(N__11725));
    LocalMux I__2822 (
            .O(N__11772),
            .I(N__11725));
    Span4Mux_v I__2821 (
            .O(N__11765),
            .I(N__11725));
    LocalMux I__2820 (
            .O(N__11762),
            .I(N__11725));
    InMux I__2819 (
            .O(N__11761),
            .I(N__11720));
    InMux I__2818 (
            .O(N__11760),
            .I(N__11720));
    InMux I__2817 (
            .O(N__11759),
            .I(N__11717));
    InMux I__2816 (
            .O(N__11758),
            .I(N__11712));
    InMux I__2815 (
            .O(N__11757),
            .I(N__11712));
    LocalMux I__2814 (
            .O(N__11754),
            .I(N__11703));
    LocalMux I__2813 (
            .O(N__11751),
            .I(N__11703));
    LocalMux I__2812 (
            .O(N__11748),
            .I(N__11703));
    Span4Mux_v I__2811 (
            .O(N__11743),
            .I(N__11703));
    Span4Mux_v I__2810 (
            .O(N__11738),
            .I(N__11700));
    Span4Mux_h I__2809 (
            .O(N__11725),
            .I(N__11697));
    LocalMux I__2808 (
            .O(N__11720),
            .I(N__11694));
    LocalMux I__2807 (
            .O(N__11717),
            .I(N__11685));
    LocalMux I__2806 (
            .O(N__11712),
            .I(N__11685));
    Sp12to4 I__2805 (
            .O(N__11703),
            .I(N__11685));
    Sp12to4 I__2804 (
            .O(N__11700),
            .I(N__11685));
    Sp12to4 I__2803 (
            .O(N__11697),
            .I(N__11682));
    Span12Mux_v I__2802 (
            .O(N__11694),
            .I(N__11679));
    Span12Mux_h I__2801 (
            .O(N__11685),
            .I(N__11676));
    Span12Mux_v I__2800 (
            .O(N__11682),
            .I(N__11673));
    Span12Mux_h I__2799 (
            .O(N__11679),
            .I(N__11668));
    Span12Mux_v I__2798 (
            .O(N__11676),
            .I(N__11668));
    Span12Mux_h I__2797 (
            .O(N__11673),
            .I(N__11665));
    Odrv12 I__2796 (
            .O(N__11668),
            .I(AGNUS_REV_c));
    Odrv12 I__2795 (
            .O(N__11665),
            .I(AGNUS_REV_c));
    InMux I__2794 (
            .O(N__11660),
            .I(N__11657));
    LocalMux I__2793 (
            .O(N__11657),
            .I(N__11654));
    Span4Mux_h I__2792 (
            .O(N__11654),
            .I(N__11651));
    Odrv4 I__2791 (
            .O(N__11651),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    ClkMux I__2790 (
            .O(N__11648),
            .I(N__11627));
    ClkMux I__2789 (
            .O(N__11647),
            .I(N__11627));
    ClkMux I__2788 (
            .O(N__11646),
            .I(N__11627));
    ClkMux I__2787 (
            .O(N__11645),
            .I(N__11627));
    ClkMux I__2786 (
            .O(N__11644),
            .I(N__11627));
    ClkMux I__2785 (
            .O(N__11643),
            .I(N__11627));
    ClkMux I__2784 (
            .O(N__11642),
            .I(N__11627));
    GlobalMux I__2783 (
            .O(N__11627),
            .I(N__11624));
    gio2CtrlBuf I__2782 (
            .O(N__11624),
            .I(C3_c_g));
    CEMux I__2781 (
            .O(N__11621),
            .I(N__11582));
    CEMux I__2780 (
            .O(N__11620),
            .I(N__11582));
    CEMux I__2779 (
            .O(N__11619),
            .I(N__11582));
    CEMux I__2778 (
            .O(N__11618),
            .I(N__11582));
    CEMux I__2777 (
            .O(N__11617),
            .I(N__11582));
    CEMux I__2776 (
            .O(N__11616),
            .I(N__11582));
    CEMux I__2775 (
            .O(N__11615),
            .I(N__11582));
    CEMux I__2774 (
            .O(N__11614),
            .I(N__11582));
    CEMux I__2773 (
            .O(N__11613),
            .I(N__11582));
    CEMux I__2772 (
            .O(N__11612),
            .I(N__11582));
    CEMux I__2771 (
            .O(N__11611),
            .I(N__11582));
    CEMux I__2770 (
            .O(N__11610),
            .I(N__11582));
    CEMux I__2769 (
            .O(N__11609),
            .I(N__11582));
    GlobalMux I__2768 (
            .O(N__11582),
            .I(N__11579));
    gio2CtrlBuf I__2767 (
            .O(N__11579),
            .I(DBRn_c_i_0_g));
    InMux I__2766 (
            .O(N__11576),
            .I(N__11566));
    InMux I__2765 (
            .O(N__11575),
            .I(N__11563));
    InMux I__2764 (
            .O(N__11574),
            .I(N__11558));
    InMux I__2763 (
            .O(N__11573),
            .I(N__11558));
    InMux I__2762 (
            .O(N__11572),
            .I(N__11555));
    InMux I__2761 (
            .O(N__11571),
            .I(N__11552));
    InMux I__2760 (
            .O(N__11570),
            .I(N__11549));
    InMux I__2759 (
            .O(N__11569),
            .I(N__11546));
    LocalMux I__2758 (
            .O(N__11566),
            .I(N__11541));
    LocalMux I__2757 (
            .O(N__11563),
            .I(N__11526));
    LocalMux I__2756 (
            .O(N__11558),
            .I(N__11523));
    LocalMux I__2755 (
            .O(N__11555),
            .I(N__11515));
    LocalMux I__2754 (
            .O(N__11552),
            .I(N__11502));
    LocalMux I__2753 (
            .O(N__11549),
            .I(N__11496));
    LocalMux I__2752 (
            .O(N__11546),
            .I(N__11485));
    SRMux I__2751 (
            .O(N__11545),
            .I(N__11366));
    SRMux I__2750 (
            .O(N__11544),
            .I(N__11366));
    Glb2LocalMux I__2749 (
            .O(N__11541),
            .I(N__11366));
    SRMux I__2748 (
            .O(N__11540),
            .I(N__11366));
    SRMux I__2747 (
            .O(N__11539),
            .I(N__11366));
    SRMux I__2746 (
            .O(N__11538),
            .I(N__11366));
    SRMux I__2745 (
            .O(N__11537),
            .I(N__11366));
    SRMux I__2744 (
            .O(N__11536),
            .I(N__11366));
    SRMux I__2743 (
            .O(N__11535),
            .I(N__11366));
    SRMux I__2742 (
            .O(N__11534),
            .I(N__11366));
    SRMux I__2741 (
            .O(N__11533),
            .I(N__11366));
    SRMux I__2740 (
            .O(N__11532),
            .I(N__11366));
    SRMux I__2739 (
            .O(N__11531),
            .I(N__11366));
    SRMux I__2738 (
            .O(N__11530),
            .I(N__11366));
    SRMux I__2737 (
            .O(N__11529),
            .I(N__11366));
    Glb2LocalMux I__2736 (
            .O(N__11526),
            .I(N__11366));
    Glb2LocalMux I__2735 (
            .O(N__11523),
            .I(N__11366));
    SRMux I__2734 (
            .O(N__11522),
            .I(N__11366));
    SRMux I__2733 (
            .O(N__11521),
            .I(N__11366));
    SRMux I__2732 (
            .O(N__11520),
            .I(N__11366));
    SRMux I__2731 (
            .O(N__11519),
            .I(N__11366));
    SRMux I__2730 (
            .O(N__11518),
            .I(N__11366));
    Glb2LocalMux I__2729 (
            .O(N__11515),
            .I(N__11366));
    SRMux I__2728 (
            .O(N__11514),
            .I(N__11366));
    SRMux I__2727 (
            .O(N__11513),
            .I(N__11366));
    SRMux I__2726 (
            .O(N__11512),
            .I(N__11366));
    SRMux I__2725 (
            .O(N__11511),
            .I(N__11366));
    SRMux I__2724 (
            .O(N__11510),
            .I(N__11366));
    SRMux I__2723 (
            .O(N__11509),
            .I(N__11366));
    SRMux I__2722 (
            .O(N__11508),
            .I(N__11366));
    SRMux I__2721 (
            .O(N__11507),
            .I(N__11366));
    SRMux I__2720 (
            .O(N__11506),
            .I(N__11366));
    SRMux I__2719 (
            .O(N__11505),
            .I(N__11366));
    Glb2LocalMux I__2718 (
            .O(N__11502),
            .I(N__11366));
    SRMux I__2717 (
            .O(N__11501),
            .I(N__11366));
    SRMux I__2716 (
            .O(N__11500),
            .I(N__11366));
    SRMux I__2715 (
            .O(N__11499),
            .I(N__11366));
    Glb2LocalMux I__2714 (
            .O(N__11496),
            .I(N__11366));
    SRMux I__2713 (
            .O(N__11495),
            .I(N__11366));
    SRMux I__2712 (
            .O(N__11494),
            .I(N__11366));
    SRMux I__2711 (
            .O(N__11493),
            .I(N__11366));
    SRMux I__2710 (
            .O(N__11492),
            .I(N__11366));
    SRMux I__2709 (
            .O(N__11491),
            .I(N__11366));
    SRMux I__2708 (
            .O(N__11490),
            .I(N__11366));
    SRMux I__2707 (
            .O(N__11489),
            .I(N__11366));
    SRMux I__2706 (
            .O(N__11488),
            .I(N__11366));
    Glb2LocalMux I__2705 (
            .O(N__11485),
            .I(N__11366));
    SRMux I__2704 (
            .O(N__11484),
            .I(N__11366));
    SRMux I__2703 (
            .O(N__11483),
            .I(N__11366));
    SRMux I__2702 (
            .O(N__11482),
            .I(N__11366));
    SRMux I__2701 (
            .O(N__11481),
            .I(N__11366));
    SRMux I__2700 (
            .O(N__11480),
            .I(N__11366));
    SRMux I__2699 (
            .O(N__11479),
            .I(N__11366));
    SRMux I__2698 (
            .O(N__11478),
            .I(N__11366));
    SRMux I__2697 (
            .O(N__11477),
            .I(N__11366));
    GlobalMux I__2696 (
            .O(N__11366),
            .I(N__11363));
    gio2CtrlBuf I__2695 (
            .O(N__11363),
            .I(RESETn_c_i_g));
    CascadeMux I__2694 (
            .O(N__11360),
            .I(N__11353));
    InMux I__2693 (
            .O(N__11359),
            .I(N__11345));
    InMux I__2692 (
            .O(N__11358),
            .I(N__11342));
    InMux I__2691 (
            .O(N__11357),
            .I(N__11339));
    CascadeMux I__2690 (
            .O(N__11356),
            .I(N__11335));
    InMux I__2689 (
            .O(N__11353),
            .I(N__11325));
    InMux I__2688 (
            .O(N__11352),
            .I(N__11325));
    InMux I__2687 (
            .O(N__11351),
            .I(N__11325));
    InMux I__2686 (
            .O(N__11350),
            .I(N__11318));
    InMux I__2685 (
            .O(N__11349),
            .I(N__11318));
    InMux I__2684 (
            .O(N__11348),
            .I(N__11318));
    LocalMux I__2683 (
            .O(N__11345),
            .I(N__11313));
    LocalMux I__2682 (
            .O(N__11342),
            .I(N__11308));
    LocalMux I__2681 (
            .O(N__11339),
            .I(N__11308));
    InMux I__2680 (
            .O(N__11338),
            .I(N__11305));
    InMux I__2679 (
            .O(N__11335),
            .I(N__11302));
    InMux I__2678 (
            .O(N__11334),
            .I(N__11295));
    InMux I__2677 (
            .O(N__11333),
            .I(N__11295));
    InMux I__2676 (
            .O(N__11332),
            .I(N__11292));
    LocalMux I__2675 (
            .O(N__11325),
            .I(N__11285));
    LocalMux I__2674 (
            .O(N__11318),
            .I(N__11285));
    InMux I__2673 (
            .O(N__11317),
            .I(N__11280));
    InMux I__2672 (
            .O(N__11316),
            .I(N__11280));
    Span4Mux_v I__2671 (
            .O(N__11313),
            .I(N__11271));
    Span4Mux_v I__2670 (
            .O(N__11308),
            .I(N__11271));
    LocalMux I__2669 (
            .O(N__11305),
            .I(N__11271));
    LocalMux I__2668 (
            .O(N__11302),
            .I(N__11271));
    InMux I__2667 (
            .O(N__11301),
            .I(N__11266));
    InMux I__2666 (
            .O(N__11300),
            .I(N__11266));
    LocalMux I__2665 (
            .O(N__11295),
            .I(N__11258));
    LocalMux I__2664 (
            .O(N__11292),
            .I(N__11258));
    InMux I__2663 (
            .O(N__11291),
            .I(N__11253));
    InMux I__2662 (
            .O(N__11290),
            .I(N__11253));
    Span4Mux_v I__2661 (
            .O(N__11285),
            .I(N__11239));
    LocalMux I__2660 (
            .O(N__11280),
            .I(N__11236));
    Span4Mux_h I__2659 (
            .O(N__11271),
            .I(N__11231));
    LocalMux I__2658 (
            .O(N__11266),
            .I(N__11231));
    InMux I__2657 (
            .O(N__11265),
            .I(N__11226));
    InMux I__2656 (
            .O(N__11264),
            .I(N__11226));
    InMux I__2655 (
            .O(N__11263),
            .I(N__11223));
    Span4Mux_v I__2654 (
            .O(N__11258),
            .I(N__11218));
    LocalMux I__2653 (
            .O(N__11253),
            .I(N__11218));
    InMux I__2652 (
            .O(N__11252),
            .I(N__11209));
    InMux I__2651 (
            .O(N__11251),
            .I(N__11209));
    InMux I__2650 (
            .O(N__11250),
            .I(N__11209));
    InMux I__2649 (
            .O(N__11249),
            .I(N__11209));
    InMux I__2648 (
            .O(N__11248),
            .I(N__11206));
    InMux I__2647 (
            .O(N__11247),
            .I(N__11197));
    InMux I__2646 (
            .O(N__11246),
            .I(N__11197));
    InMux I__2645 (
            .O(N__11245),
            .I(N__11197));
    InMux I__2644 (
            .O(N__11244),
            .I(N__11197));
    InMux I__2643 (
            .O(N__11243),
            .I(N__11187));
    InMux I__2642 (
            .O(N__11242),
            .I(N__11187));
    Span4Mux_h I__2641 (
            .O(N__11239),
            .I(N__11178));
    Span4Mux_v I__2640 (
            .O(N__11236),
            .I(N__11178));
    Span4Mux_v I__2639 (
            .O(N__11231),
            .I(N__11178));
    LocalMux I__2638 (
            .O(N__11226),
            .I(N__11178));
    LocalMux I__2637 (
            .O(N__11223),
            .I(N__11175));
    Sp12to4 I__2636 (
            .O(N__11218),
            .I(N__11170));
    LocalMux I__2635 (
            .O(N__11209),
            .I(N__11170));
    LocalMux I__2634 (
            .O(N__11206),
            .I(N__11167));
    LocalMux I__2633 (
            .O(N__11197),
            .I(N__11164));
    InMux I__2632 (
            .O(N__11196),
            .I(N__11155));
    InMux I__2631 (
            .O(N__11195),
            .I(N__11155));
    InMux I__2630 (
            .O(N__11194),
            .I(N__11155));
    InMux I__2629 (
            .O(N__11193),
            .I(N__11155));
    InMux I__2628 (
            .O(N__11192),
            .I(N__11152));
    LocalMux I__2627 (
            .O(N__11187),
            .I(N__11149));
    Span4Mux_h I__2626 (
            .O(N__11178),
            .I(N__11144));
    Span4Mux_v I__2625 (
            .O(N__11175),
            .I(N__11144));
    Span12Mux_v I__2624 (
            .O(N__11170),
            .I(N__11141));
    Span12Mux_v I__2623 (
            .O(N__11167),
            .I(N__11132));
    Span12Mux_v I__2622 (
            .O(N__11164),
            .I(N__11132));
    LocalMux I__2621 (
            .O(N__11155),
            .I(N__11132));
    LocalMux I__2620 (
            .O(N__11152),
            .I(N__11132));
    Span12Mux_v I__2619 (
            .O(N__11149),
            .I(N__11129));
    Span4Mux_h I__2618 (
            .O(N__11144),
            .I(N__11126));
    Span12Mux_h I__2617 (
            .O(N__11141),
            .I(N__11123));
    Span12Mux_h I__2616 (
            .O(N__11132),
            .I(N__11120));
    Span12Mux_h I__2615 (
            .O(N__11129),
            .I(N__11117));
    Span4Mux_h I__2614 (
            .O(N__11126),
            .I(N__11114));
    Odrv12 I__2613 (
            .O(N__11123),
            .I(RESETn_c));
    Odrv12 I__2612 (
            .O(N__11120),
            .I(RESETn_c));
    Odrv12 I__2611 (
            .O(N__11117),
            .I(RESETn_c));
    Odrv4 I__2610 (
            .O(N__11114),
            .I(RESETn_c));
    InMux I__2609 (
            .O(N__11105),
            .I(N__11102));
    LocalMux I__2608 (
            .O(N__11102),
            .I(N__11099));
    Span12Mux_h I__2607 (
            .O(N__11099),
            .I(N__11096));
    Odrv12 I__2606 (
            .O(N__11096),
            .I(RAS1n_c));
    InMux I__2605 (
            .O(N__11093),
            .I(N__11090));
    LocalMux I__2604 (
            .O(N__11090),
            .I(N__11086));
    InMux I__2603 (
            .O(N__11089),
            .I(N__11083));
    Sp12to4 I__2602 (
            .O(N__11086),
            .I(N__11080));
    LocalMux I__2601 (
            .O(N__11083),
            .I(N__11077));
    Span12Mux_v I__2600 (
            .O(N__11080),
            .I(N__11074));
    Span12Mux_h I__2599 (
            .O(N__11077),
            .I(N__11071));
    Odrv12 I__2598 (
            .O(N__11074),
            .I(RAS0n_c));
    Odrv12 I__2597 (
            .O(N__11071),
            .I(RAS0n_c));
    InMux I__2596 (
            .O(N__11066),
            .I(N__11063));
    LocalMux I__2595 (
            .O(N__11063),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2594 (
            .O(N__11060),
            .I(N__11057));
    LocalMux I__2593 (
            .O(N__11057),
            .I(N__11026));
    ClkMux I__2592 (
            .O(N__11056),
            .I(N__10892));
    ClkMux I__2591 (
            .O(N__11055),
            .I(N__10892));
    ClkMux I__2590 (
            .O(N__11054),
            .I(N__10892));
    ClkMux I__2589 (
            .O(N__11053),
            .I(N__10892));
    ClkMux I__2588 (
            .O(N__11052),
            .I(N__10892));
    ClkMux I__2587 (
            .O(N__11051),
            .I(N__10892));
    ClkMux I__2586 (
            .O(N__11050),
            .I(N__10892));
    ClkMux I__2585 (
            .O(N__11049),
            .I(N__10892));
    ClkMux I__2584 (
            .O(N__11048),
            .I(N__10892));
    ClkMux I__2583 (
            .O(N__11047),
            .I(N__10892));
    ClkMux I__2582 (
            .O(N__11046),
            .I(N__10892));
    ClkMux I__2581 (
            .O(N__11045),
            .I(N__10892));
    ClkMux I__2580 (
            .O(N__11044),
            .I(N__10892));
    ClkMux I__2579 (
            .O(N__11043),
            .I(N__10892));
    ClkMux I__2578 (
            .O(N__11042),
            .I(N__10892));
    ClkMux I__2577 (
            .O(N__11041),
            .I(N__10892));
    ClkMux I__2576 (
            .O(N__11040),
            .I(N__10892));
    ClkMux I__2575 (
            .O(N__11039),
            .I(N__10892));
    ClkMux I__2574 (
            .O(N__11038),
            .I(N__10892));
    ClkMux I__2573 (
            .O(N__11037),
            .I(N__10892));
    ClkMux I__2572 (
            .O(N__11036),
            .I(N__10892));
    ClkMux I__2571 (
            .O(N__11035),
            .I(N__10892));
    ClkMux I__2570 (
            .O(N__11034),
            .I(N__10892));
    ClkMux I__2569 (
            .O(N__11033),
            .I(N__10892));
    ClkMux I__2568 (
            .O(N__11032),
            .I(N__10892));
    ClkMux I__2567 (
            .O(N__11031),
            .I(N__10892));
    ClkMux I__2566 (
            .O(N__11030),
            .I(N__10892));
    ClkMux I__2565 (
            .O(N__11029),
            .I(N__10892));
    Glb2LocalMux I__2564 (
            .O(N__11026),
            .I(N__10892));
    ClkMux I__2563 (
            .O(N__11025),
            .I(N__10892));
    ClkMux I__2562 (
            .O(N__11024),
            .I(N__10892));
    ClkMux I__2561 (
            .O(N__11023),
            .I(N__10892));
    ClkMux I__2560 (
            .O(N__11022),
            .I(N__10892));
    ClkMux I__2559 (
            .O(N__11021),
            .I(N__10892));
    ClkMux I__2558 (
            .O(N__11020),
            .I(N__10892));
    ClkMux I__2557 (
            .O(N__11019),
            .I(N__10892));
    ClkMux I__2556 (
            .O(N__11018),
            .I(N__10892));
    ClkMux I__2555 (
            .O(N__11017),
            .I(N__10892));
    ClkMux I__2554 (
            .O(N__11016),
            .I(N__10892));
    ClkMux I__2553 (
            .O(N__11015),
            .I(N__10892));
    ClkMux I__2552 (
            .O(N__11014),
            .I(N__10892));
    ClkMux I__2551 (
            .O(N__11013),
            .I(N__10892));
    ClkMux I__2550 (
            .O(N__11012),
            .I(N__10892));
    ClkMux I__2549 (
            .O(N__11011),
            .I(N__10892));
    ClkMux I__2548 (
            .O(N__11010),
            .I(N__10892));
    ClkMux I__2547 (
            .O(N__11009),
            .I(N__10892));
    ClkMux I__2546 (
            .O(N__11008),
            .I(N__10892));
    ClkMux I__2545 (
            .O(N__11007),
            .I(N__10892));
    ClkMux I__2544 (
            .O(N__11006),
            .I(N__10892));
    ClkMux I__2543 (
            .O(N__11005),
            .I(N__10892));
    ClkMux I__2542 (
            .O(N__11004),
            .I(N__10892));
    ClkMux I__2541 (
            .O(N__11003),
            .I(N__10892));
    ClkMux I__2540 (
            .O(N__11002),
            .I(N__10892));
    ClkMux I__2539 (
            .O(N__11001),
            .I(N__10892));
    GlobalMux I__2538 (
            .O(N__10892),
            .I(CLK80_PLL));
    InMux I__2537 (
            .O(N__10889),
            .I(N__10884));
    CascadeMux I__2536 (
            .O(N__10888),
            .I(N__10881));
    InMux I__2535 (
            .O(N__10887),
            .I(N__10877));
    LocalMux I__2534 (
            .O(N__10884),
            .I(N__10874));
    InMux I__2533 (
            .O(N__10881),
            .I(N__10871));
    InMux I__2532 (
            .O(N__10880),
            .I(N__10867));
    LocalMux I__2531 (
            .O(N__10877),
            .I(N__10864));
    Span4Mux_h I__2530 (
            .O(N__10874),
            .I(N__10859));
    LocalMux I__2529 (
            .O(N__10871),
            .I(N__10859));
    InMux I__2528 (
            .O(N__10870),
            .I(N__10856));
    LocalMux I__2527 (
            .O(N__10867),
            .I(N__10853));
    Span4Mux_v I__2526 (
            .O(N__10864),
            .I(N__10850));
    Span4Mux_v I__2525 (
            .O(N__10859),
            .I(N__10845));
    LocalMux I__2524 (
            .O(N__10856),
            .I(N__10845));
    Span4Mux_v I__2523 (
            .O(N__10853),
            .I(N__10842));
    Span4Mux_v I__2522 (
            .O(N__10850),
            .I(N__10839));
    Span4Mux_h I__2521 (
            .O(N__10845),
            .I(N__10836));
    Sp12to4 I__2520 (
            .O(N__10842),
            .I(N__10833));
    Sp12to4 I__2519 (
            .O(N__10839),
            .I(N__10830));
    Sp12to4 I__2518 (
            .O(N__10836),
            .I(N__10827));
    Span12Mux_h I__2517 (
            .O(N__10833),
            .I(N__10824));
    Span12Mux_h I__2516 (
            .O(N__10830),
            .I(N__10819));
    Span12Mux_v I__2515 (
            .O(N__10827),
            .I(N__10819));
    Span12Mux_v I__2514 (
            .O(N__10824),
            .I(N__10816));
    Span12Mux_h I__2513 (
            .O(N__10819),
            .I(N__10813));
    Odrv12 I__2512 (
            .O(N__10816),
            .I(RnW_c));
    Odrv12 I__2511 (
            .O(N__10813),
            .I(RnW_c));
    InMux I__2510 (
            .O(N__10808),
            .I(N__10804));
    InMux I__2509 (
            .O(N__10807),
            .I(N__10801));
    LocalMux I__2508 (
            .O(N__10804),
            .I(N__10798));
    LocalMux I__2507 (
            .O(N__10801),
            .I(N__10795));
    Span12Mux_s8_h I__2506 (
            .O(N__10798),
            .I(N__10792));
    Span12Mux_h I__2505 (
            .O(N__10795),
            .I(N__10789));
    Span12Mux_v I__2504 (
            .O(N__10792),
            .I(N__10783));
    Span12Mux_v I__2503 (
            .O(N__10789),
            .I(N__10783));
    InMux I__2502 (
            .O(N__10788),
            .I(N__10780));
    Odrv12 I__2501 (
            .O(N__10783),
            .I(DMA_WRITE_CYCLE));
    LocalMux I__2500 (
            .O(N__10780),
            .I(DMA_WRITE_CYCLE));
    CascadeMux I__2499 (
            .O(N__10775),
            .I(N__10772));
    InMux I__2498 (
            .O(N__10772),
            .I(N__10768));
    CascadeMux I__2497 (
            .O(N__10771),
            .I(N__10765));
    LocalMux I__2496 (
            .O(N__10768),
            .I(N__10759));
    InMux I__2495 (
            .O(N__10765),
            .I(N__10756));
    InMux I__2494 (
            .O(N__10764),
            .I(N__10753));
    CascadeMux I__2493 (
            .O(N__10763),
            .I(N__10750));
    InMux I__2492 (
            .O(N__10762),
            .I(N__10747));
    Span4Mux_v I__2491 (
            .O(N__10759),
            .I(N__10740));
    LocalMux I__2490 (
            .O(N__10756),
            .I(N__10740));
    LocalMux I__2489 (
            .O(N__10753),
            .I(N__10740));
    InMux I__2488 (
            .O(N__10750),
            .I(N__10737));
    LocalMux I__2487 (
            .O(N__10747),
            .I(N__10734));
    Span4Mux_v I__2486 (
            .O(N__10740),
            .I(N__10731));
    LocalMux I__2485 (
            .O(N__10737),
            .I(N__10728));
    Span4Mux_v I__2484 (
            .O(N__10734),
            .I(N__10724));
    Span4Mux_h I__2483 (
            .O(N__10731),
            .I(N__10719));
    Span4Mux_v I__2482 (
            .O(N__10728),
            .I(N__10719));
    CascadeMux I__2481 (
            .O(N__10727),
            .I(N__10716));
    Span4Mux_v I__2480 (
            .O(N__10724),
            .I(N__10713));
    Sp12to4 I__2479 (
            .O(N__10719),
            .I(N__10710));
    InMux I__2478 (
            .O(N__10716),
            .I(N__10707));
    Sp12to4 I__2477 (
            .O(N__10713),
            .I(N__10704));
    Span12Mux_h I__2476 (
            .O(N__10710),
            .I(N__10699));
    LocalMux I__2475 (
            .O(N__10707),
            .I(N__10699));
    Span12Mux_h I__2474 (
            .O(N__10704),
            .I(N__10694));
    Span12Mux_v I__2473 (
            .O(N__10699),
            .I(N__10694));
    Odrv12 I__2472 (
            .O(N__10694),
            .I(CASLn_c));
    InMux I__2471 (
            .O(N__10691),
            .I(N__10686));
    InMux I__2470 (
            .O(N__10690),
            .I(N__10683));
    InMux I__2469 (
            .O(N__10689),
            .I(N__10680));
    LocalMux I__2468 (
            .O(N__10686),
            .I(N__10674));
    LocalMux I__2467 (
            .O(N__10683),
            .I(N__10674));
    LocalMux I__2466 (
            .O(N__10680),
            .I(N__10671));
    InMux I__2465 (
            .O(N__10679),
            .I(N__10668));
    Span4Mux_v I__2464 (
            .O(N__10674),
            .I(N__10663));
    Span4Mux_v I__2463 (
            .O(N__10671),
            .I(N__10658));
    LocalMux I__2462 (
            .O(N__10668),
            .I(N__10658));
    InMux I__2461 (
            .O(N__10667),
            .I(N__10655));
    InMux I__2460 (
            .O(N__10666),
            .I(N__10652));
    Sp12to4 I__2459 (
            .O(N__10663),
            .I(N__10649));
    Sp12to4 I__2458 (
            .O(N__10658),
            .I(N__10644));
    LocalMux I__2457 (
            .O(N__10655),
            .I(N__10644));
    LocalMux I__2456 (
            .O(N__10652),
            .I(N__10641));
    Span12Mux_h I__2455 (
            .O(N__10649),
            .I(N__10638));
    Span12Mux_v I__2454 (
            .O(N__10644),
            .I(N__10635));
    Span4Mux_h I__2453 (
            .O(N__10641),
            .I(N__10632));
    Span12Mux_v I__2452 (
            .O(N__10638),
            .I(N__10629));
    Span12Mux_h I__2451 (
            .O(N__10635),
            .I(N__10626));
    Span4Mux_v I__2450 (
            .O(N__10632),
            .I(N__10623));
    Odrv12 I__2449 (
            .O(N__10629),
            .I(CASUn_c));
    Odrv12 I__2448 (
            .O(N__10626),
            .I(CASUn_c));
    Odrv4 I__2447 (
            .O(N__10623),
            .I(CASUn_c));
    CascadeMux I__2446 (
            .O(N__10616),
            .I(N__10613));
    InMux I__2445 (
            .O(N__10613),
            .I(N__10606));
    CascadeMux I__2444 (
            .O(N__10612),
            .I(N__10602));
    InMux I__2443 (
            .O(N__10611),
            .I(N__10594));
    InMux I__2442 (
            .O(N__10610),
            .I(N__10591));
    InMux I__2441 (
            .O(N__10609),
            .I(N__10588));
    LocalMux I__2440 (
            .O(N__10606),
            .I(N__10583));
    InMux I__2439 (
            .O(N__10605),
            .I(N__10576));
    InMux I__2438 (
            .O(N__10602),
            .I(N__10576));
    InMux I__2437 (
            .O(N__10601),
            .I(N__10576));
    InMux I__2436 (
            .O(N__10600),
            .I(N__10569));
    InMux I__2435 (
            .O(N__10599),
            .I(N__10569));
    InMux I__2434 (
            .O(N__10598),
            .I(N__10569));
    CascadeMux I__2433 (
            .O(N__10597),
            .I(N__10566));
    LocalMux I__2432 (
            .O(N__10594),
            .I(N__10563));
    LocalMux I__2431 (
            .O(N__10591),
            .I(N__10555));
    LocalMux I__2430 (
            .O(N__10588),
            .I(N__10555));
    InMux I__2429 (
            .O(N__10587),
            .I(N__10543));
    InMux I__2428 (
            .O(N__10586),
            .I(N__10543));
    Span4Mux_v I__2427 (
            .O(N__10583),
            .I(N__10534));
    LocalMux I__2426 (
            .O(N__10576),
            .I(N__10534));
    LocalMux I__2425 (
            .O(N__10569),
            .I(N__10534));
    InMux I__2424 (
            .O(N__10566),
            .I(N__10531));
    Span4Mux_v I__2423 (
            .O(N__10563),
            .I(N__10528));
    InMux I__2422 (
            .O(N__10562),
            .I(N__10525));
    InMux I__2421 (
            .O(N__10561),
            .I(N__10520));
    InMux I__2420 (
            .O(N__10560),
            .I(N__10520));
    Span4Mux_v I__2419 (
            .O(N__10555),
            .I(N__10517));
    InMux I__2418 (
            .O(N__10554),
            .I(N__10514));
    InMux I__2417 (
            .O(N__10553),
            .I(N__10503));
    InMux I__2416 (
            .O(N__10552),
            .I(N__10503));
    InMux I__2415 (
            .O(N__10551),
            .I(N__10503));
    InMux I__2414 (
            .O(N__10550),
            .I(N__10503));
    InMux I__2413 (
            .O(N__10549),
            .I(N__10503));
    InMux I__2412 (
            .O(N__10548),
            .I(N__10499));
    LocalMux I__2411 (
            .O(N__10543),
            .I(N__10496));
    InMux I__2410 (
            .O(N__10542),
            .I(N__10493));
    InMux I__2409 (
            .O(N__10541),
            .I(N__10490));
    Span4Mux_h I__2408 (
            .O(N__10534),
            .I(N__10487));
    LocalMux I__2407 (
            .O(N__10531),
            .I(N__10472));
    Sp12to4 I__2406 (
            .O(N__10528),
            .I(N__10472));
    LocalMux I__2405 (
            .O(N__10525),
            .I(N__10472));
    LocalMux I__2404 (
            .O(N__10520),
            .I(N__10472));
    Sp12to4 I__2403 (
            .O(N__10517),
            .I(N__10472));
    LocalMux I__2402 (
            .O(N__10514),
            .I(N__10472));
    LocalMux I__2401 (
            .O(N__10503),
            .I(N__10472));
    InMux I__2400 (
            .O(N__10502),
            .I(N__10469));
    LocalMux I__2399 (
            .O(N__10499),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2398 (
            .O(N__10496),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2397 (
            .O(N__10493),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2396 (
            .O(N__10490),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2395 (
            .O(N__10487),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__2394 (
            .O(N__10472),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2393 (
            .O(N__10469),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__2392 (
            .O(N__10454),
            .I(N__10451));
    LocalMux I__2391 (
            .O(N__10451),
            .I(N__10448));
    Span4Mux_s3_v I__2390 (
            .O(N__10448),
            .I(N__10445));
    Span4Mux_v I__2389 (
            .O(N__10445),
            .I(N__10442));
    Sp12to4 I__2388 (
            .O(N__10442),
            .I(N__10439));
    Span12Mux_h I__2387 (
            .O(N__10439),
            .I(N__10436));
    Odrv12 I__2386 (
            .O(N__10436),
            .I(CASn_c));
    InMux I__2385 (
            .O(N__10433),
            .I(N__10430));
    LocalMux I__2384 (
            .O(N__10430),
            .I(N__10426));
    InMux I__2383 (
            .O(N__10429),
            .I(N__10423));
    Span4Mux_v I__2382 (
            .O(N__10426),
            .I(N__10416));
    LocalMux I__2381 (
            .O(N__10423),
            .I(N__10416));
    CascadeMux I__2380 (
            .O(N__10422),
            .I(N__10412));
    InMux I__2379 (
            .O(N__10421),
            .I(N__10408));
    Span4Mux_h I__2378 (
            .O(N__10416),
            .I(N__10405));
    InMux I__2377 (
            .O(N__10415),
            .I(N__10400));
    InMux I__2376 (
            .O(N__10412),
            .I(N__10400));
    InMux I__2375 (
            .O(N__10411),
            .I(N__10397));
    LocalMux I__2374 (
            .O(N__10408),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2373 (
            .O(N__10405),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__2372 (
            .O(N__10400),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__2371 (
            .O(N__10397),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__2370 (
            .O(N__10388),
            .I(N__10385));
    LocalMux I__2369 (
            .O(N__10385),
            .I(N__10382));
    Span4Mux_s3_v I__2368 (
            .O(N__10382),
            .I(N__10379));
    Span4Mux_v I__2367 (
            .O(N__10379),
            .I(N__10376));
    Span4Mux_h I__2366 (
            .O(N__10376),
            .I(N__10373));
    Odrv4 I__2365 (
            .O(N__10373),
            .I(RASn_c));
    CascadeMux I__2364 (
            .O(N__10370),
            .I(N__10367));
    InMux I__2363 (
            .O(N__10367),
            .I(N__10364));
    LocalMux I__2362 (
            .O(N__10364),
            .I(N__10361));
    Span4Mux_h I__2361 (
            .O(N__10361),
            .I(N__10358));
    Odrv4 I__2360 (
            .O(N__10358),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2359 (
            .O(N__10355),
            .I(N__10349));
    InMux I__2358 (
            .O(N__10354),
            .I(N__10344));
    InMux I__2357 (
            .O(N__10353),
            .I(N__10344));
    InMux I__2356 (
            .O(N__10352),
            .I(N__10341));
    LocalMux I__2355 (
            .O(N__10349),
            .I(N__10338));
    LocalMux I__2354 (
            .O(N__10344),
            .I(N__10333));
    LocalMux I__2353 (
            .O(N__10341),
            .I(N__10333));
    Span4Mux_v I__2352 (
            .O(N__10338),
            .I(N__10330));
    Span12Mux_v I__2351 (
            .O(N__10333),
            .I(N__10327));
    Span4Mux_v I__2350 (
            .O(N__10330),
            .I(N__10324));
    Span12Mux_h I__2349 (
            .O(N__10327),
            .I(N__10321));
    Sp12to4 I__2348 (
            .O(N__10324),
            .I(N__10318));
    Odrv12 I__2347 (
            .O(N__10321),
            .I(DRA_c_5));
    Odrv12 I__2346 (
            .O(N__10318),
            .I(DRA_c_5));
    InMux I__2345 (
            .O(N__10313),
            .I(N__10309));
    InMux I__2344 (
            .O(N__10312),
            .I(N__10306));
    LocalMux I__2343 (
            .O(N__10309),
            .I(N__10299));
    LocalMux I__2342 (
            .O(N__10306),
            .I(N__10299));
    InMux I__2341 (
            .O(N__10305),
            .I(N__10296));
    InMux I__2340 (
            .O(N__10304),
            .I(N__10293));
    Span4Mux_h I__2339 (
            .O(N__10299),
            .I(N__10288));
    LocalMux I__2338 (
            .O(N__10296),
            .I(N__10288));
    LocalMux I__2337 (
            .O(N__10293),
            .I(N__10283));
    Sp12to4 I__2336 (
            .O(N__10288),
            .I(N__10283));
    Span12Mux_v I__2335 (
            .O(N__10283),
            .I(N__10280));
    Span12Mux_h I__2334 (
            .O(N__10280),
            .I(N__10277));
    Odrv12 I__2333 (
            .O(N__10277),
            .I(DRA_c_4));
    InMux I__2332 (
            .O(N__10274),
            .I(N__10271));
    LocalMux I__2331 (
            .O(N__10271),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__2330 (
            .O(N__10268),
            .I(N__10264));
    InMux I__2329 (
            .O(N__10267),
            .I(N__10261));
    LocalMux I__2328 (
            .O(N__10264),
            .I(N__10256));
    LocalMux I__2327 (
            .O(N__10261),
            .I(N__10256));
    Span4Mux_h I__2326 (
            .O(N__10256),
            .I(N__10253));
    Odrv4 I__2325 (
            .O(N__10253),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2324 (
            .O(N__10250),
            .I(N__10246));
    InMux I__2323 (
            .O(N__10249),
            .I(N__10243));
    LocalMux I__2322 (
            .O(N__10246),
            .I(N__10240));
    LocalMux I__2321 (
            .O(N__10243),
            .I(N__10235));
    Span4Mux_v I__2320 (
            .O(N__10240),
            .I(N__10232));
    InMux I__2319 (
            .O(N__10239),
            .I(N__10229));
    InMux I__2318 (
            .O(N__10238),
            .I(N__10226));
    Sp12to4 I__2317 (
            .O(N__10235),
            .I(N__10223));
    Sp12to4 I__2316 (
            .O(N__10232),
            .I(N__10216));
    LocalMux I__2315 (
            .O(N__10229),
            .I(N__10216));
    LocalMux I__2314 (
            .O(N__10226),
            .I(N__10216));
    Span12Mux_v I__2313 (
            .O(N__10223),
            .I(N__10213));
    Span12Mux_h I__2312 (
            .O(N__10216),
            .I(N__10210));
    Span12Mux_h I__2311 (
            .O(N__10213),
            .I(N__10205));
    Span12Mux_v I__2310 (
            .O(N__10210),
            .I(N__10205));
    Odrv12 I__2309 (
            .O(N__10205),
            .I(DRA_c_1));
    InMux I__2308 (
            .O(N__10202),
            .I(N__10198));
    InMux I__2307 (
            .O(N__10201),
            .I(N__10195));
    LocalMux I__2306 (
            .O(N__10198),
            .I(N__10190));
    LocalMux I__2305 (
            .O(N__10195),
            .I(N__10190));
    Sp12to4 I__2304 (
            .O(N__10190),
            .I(N__10187));
    Span12Mux_v I__2303 (
            .O(N__10187),
            .I(N__10184));
    Span12Mux_h I__2302 (
            .O(N__10184),
            .I(N__10181));
    Odrv12 I__2301 (
            .O(N__10181),
            .I(DRA_c_0));
    InMux I__2300 (
            .O(N__10178),
            .I(N__10175));
    LocalMux I__2299 (
            .O(N__10175),
            .I(N__10172));
    Span4Mux_h I__2298 (
            .O(N__10172),
            .I(N__10169));
    Odrv4 I__2297 (
            .O(N__10169),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__2296 (
            .O(N__10166),
            .I(N__10163));
    LocalMux I__2295 (
            .O(N__10163),
            .I(N__10160));
    Odrv12 I__2294 (
            .O(N__10160),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ));
    InMux I__2293 (
            .O(N__10157),
            .I(N__10154));
    LocalMux I__2292 (
            .O(N__10154),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__2291 (
            .O(N__10151),
            .I(N__10148));
    LocalMux I__2290 (
            .O(N__10148),
            .I(N__10145));
    Span4Mux_h I__2289 (
            .O(N__10145),
            .I(N__10142));
    Odrv4 I__2288 (
            .O(N__10142),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2287 (
            .O(N__10139),
            .I(N__10136));
    LocalMux I__2286 (
            .O(N__10136),
            .I(N__10133));
    Span4Mux_h I__2285 (
            .O(N__10133),
            .I(N__10130));
    Odrv4 I__2284 (
            .O(N__10130),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2283 (
            .O(N__10127),
            .I(N__10124));
    LocalMux I__2282 (
            .O(N__10124),
            .I(N__10121));
    Span4Mux_h I__2281 (
            .O(N__10121),
            .I(N__10118));
    Odrv4 I__2280 (
            .O(N__10118),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    CascadeMux I__2279 (
            .O(N__10115),
            .I(N__10112));
    InMux I__2278 (
            .O(N__10112),
            .I(N__10109));
    LocalMux I__2277 (
            .O(N__10109),
            .I(N__10106));
    Span4Mux_v I__2276 (
            .O(N__10106),
            .I(N__10103));
    Odrv4 I__2275 (
            .O(N__10103),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2274 (
            .O(N__10100),
            .I(N__10095));
    InMux I__2273 (
            .O(N__10099),
            .I(N__10092));
    InMux I__2272 (
            .O(N__10098),
            .I(N__10089));
    LocalMux I__2271 (
            .O(N__10095),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    LocalMux I__2270 (
            .O(N__10092),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    LocalMux I__2269 (
            .O(N__10089),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    CascadeMux I__2268 (
            .O(N__10082),
            .I(N__10075));
    CascadeMux I__2267 (
            .O(N__10081),
            .I(N__10072));
    InMux I__2266 (
            .O(N__10080),
            .I(N__10069));
    InMux I__2265 (
            .O(N__10079),
            .I(N__10066));
    InMux I__2264 (
            .O(N__10078),
            .I(N__10063));
    InMux I__2263 (
            .O(N__10075),
            .I(N__10060));
    InMux I__2262 (
            .O(N__10072),
            .I(N__10057));
    LocalMux I__2261 (
            .O(N__10069),
            .I(N__10054));
    LocalMux I__2260 (
            .O(N__10066),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__2259 (
            .O(N__10063),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__2258 (
            .O(N__10060),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__2257 (
            .O(N__10057),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    Odrv4 I__2256 (
            .O(N__10054),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    CascadeMux I__2255 (
            .O(N__10043),
            .I(N__10034));
    InMux I__2254 (
            .O(N__10042),
            .I(N__10023));
    InMux I__2253 (
            .O(N__10041),
            .I(N__10023));
    InMux I__2252 (
            .O(N__10040),
            .I(N__10023));
    InMux I__2251 (
            .O(N__10039),
            .I(N__10016));
    InMux I__2250 (
            .O(N__10038),
            .I(N__10016));
    InMux I__2249 (
            .O(N__10037),
            .I(N__10016));
    InMux I__2248 (
            .O(N__10034),
            .I(N__10013));
    InMux I__2247 (
            .O(N__10033),
            .I(N__10006));
    InMux I__2246 (
            .O(N__10032),
            .I(N__10006));
    InMux I__2245 (
            .O(N__10031),
            .I(N__10006));
    InMux I__2244 (
            .O(N__10030),
            .I(N__10003));
    LocalMux I__2243 (
            .O(N__10023),
            .I(N__10000));
    LocalMux I__2242 (
            .O(N__10016),
            .I(N__9997));
    LocalMux I__2241 (
            .O(N__10013),
            .I(N__9994));
    LocalMux I__2240 (
            .O(N__10006),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__2239 (
            .O(N__10003),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__2238 (
            .O(N__10000),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__2237 (
            .O(N__9997),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__2236 (
            .O(N__9994),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__2235 (
            .O(N__9983),
            .I(N__9980));
    LocalMux I__2234 (
            .O(N__9980),
            .I(N__9974));
    CascadeMux I__2233 (
            .O(N__9979),
            .I(N__9971));
    InMux I__2232 (
            .O(N__9978),
            .I(N__9968));
    CascadeMux I__2231 (
            .O(N__9977),
            .I(N__9964));
    Span4Mux_v I__2230 (
            .O(N__9974),
            .I(N__9959));
    InMux I__2229 (
            .O(N__9971),
            .I(N__9956));
    LocalMux I__2228 (
            .O(N__9968),
            .I(N__9953));
    InMux I__2227 (
            .O(N__9967),
            .I(N__9950));
    InMux I__2226 (
            .O(N__9964),
            .I(N__9947));
    InMux I__2225 (
            .O(N__9963),
            .I(N__9942));
    InMux I__2224 (
            .O(N__9962),
            .I(N__9942));
    Span4Mux_h I__2223 (
            .O(N__9959),
            .I(N__9937));
    LocalMux I__2222 (
            .O(N__9956),
            .I(N__9937));
    Span4Mux_h I__2221 (
            .O(N__9953),
            .I(N__9934));
    LocalMux I__2220 (
            .O(N__9950),
            .I(N__9931));
    LocalMux I__2219 (
            .O(N__9947),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    LocalMux I__2218 (
            .O(N__9942),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    Odrv4 I__2217 (
            .O(N__9937),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    Odrv4 I__2216 (
            .O(N__9934),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    Odrv4 I__2215 (
            .O(N__9931),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    InMux I__2214 (
            .O(N__9920),
            .I(N__9917));
    LocalMux I__2213 (
            .O(N__9917),
            .I(\U712_REG_SM.N_400 ));
    IoInMux I__2212 (
            .O(N__9914),
            .I(N__9911));
    LocalMux I__2211 (
            .O(N__9911),
            .I(N__9908));
    Span4Mux_s2_v I__2210 (
            .O(N__9908),
            .I(N__9905));
    Span4Mux_h I__2209 (
            .O(N__9905),
            .I(N__9902));
    Span4Mux_h I__2208 (
            .O(N__9902),
            .I(N__9898));
    CascadeMux I__2207 (
            .O(N__9901),
            .I(N__9895));
    Sp12to4 I__2206 (
            .O(N__9898),
            .I(N__9892));
    InMux I__2205 (
            .O(N__9895),
            .I(N__9889));
    Odrv12 I__2204 (
            .O(N__9892),
            .I(UDSn_c));
    LocalMux I__2203 (
            .O(N__9889),
            .I(UDSn_c));
    InMux I__2202 (
            .O(N__9884),
            .I(N__9879));
    InMux I__2201 (
            .O(N__9883),
            .I(N__9873));
    InMux I__2200 (
            .O(N__9882),
            .I(N__9873));
    LocalMux I__2199 (
            .O(N__9879),
            .I(N__9870));
    InMux I__2198 (
            .O(N__9878),
            .I(N__9867));
    LocalMux I__2197 (
            .O(N__9873),
            .I(N__9864));
    Odrv4 I__2196 (
            .O(N__9870),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    LocalMux I__2195 (
            .O(N__9867),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    Odrv4 I__2194 (
            .O(N__9864),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    IoInMux I__2193 (
            .O(N__9857),
            .I(N__9854));
    LocalMux I__2192 (
            .O(N__9854),
            .I(N__9851));
    IoSpan4Mux I__2191 (
            .O(N__9851),
            .I(N__9848));
    Sp12to4 I__2190 (
            .O(N__9848),
            .I(N__9845));
    Span12Mux_v I__2189 (
            .O(N__9845),
            .I(N__9841));
    InMux I__2188 (
            .O(N__9844),
            .I(N__9838));
    Odrv12 I__2187 (
            .O(N__9841),
            .I(PRnW_c));
    LocalMux I__2186 (
            .O(N__9838),
            .I(PRnW_c));
    InMux I__2185 (
            .O(N__9833),
            .I(N__9830));
    LocalMux I__2184 (
            .O(N__9830),
            .I(\U712_REG_SM.N_398 ));
    IoInMux I__2183 (
            .O(N__9827),
            .I(N__9824));
    LocalMux I__2182 (
            .O(N__9824),
            .I(N__9821));
    Span4Mux_s3_v I__2181 (
            .O(N__9821),
            .I(N__9818));
    Sp12to4 I__2180 (
            .O(N__9818),
            .I(N__9814));
    CascadeMux I__2179 (
            .O(N__9817),
            .I(N__9811));
    Span12Mux_h I__2178 (
            .O(N__9814),
            .I(N__9808));
    InMux I__2177 (
            .O(N__9811),
            .I(N__9805));
    Odrv12 I__2176 (
            .O(N__9808),
            .I(LDSn_c));
    LocalMux I__2175 (
            .O(N__9805),
            .I(LDSn_c));
    IoInMux I__2174 (
            .O(N__9800),
            .I(N__9797));
    LocalMux I__2173 (
            .O(N__9797),
            .I(N__9794));
    IoSpan4Mux I__2172 (
            .O(N__9794),
            .I(N__9791));
    Span4Mux_s2_v I__2171 (
            .O(N__9791),
            .I(N__9788));
    Span4Mux_v I__2170 (
            .O(N__9788),
            .I(N__9785));
    Odrv4 I__2169 (
            .O(N__9785),
            .I(N_325_i));
    IoInMux I__2168 (
            .O(N__9782),
            .I(N__9779));
    LocalMux I__2167 (
            .O(N__9779),
            .I(N__9776));
    Span4Mux_s2_v I__2166 (
            .O(N__9776),
            .I(N__9773));
    Span4Mux_v I__2165 (
            .O(N__9773),
            .I(N__9770));
    Odrv4 I__2164 (
            .O(N__9770),
            .I(N_323_i));
    InMux I__2163 (
            .O(N__9767),
            .I(N__9762));
    InMux I__2162 (
            .O(N__9766),
            .I(N__9757));
    InMux I__2161 (
            .O(N__9765),
            .I(N__9757));
    LocalMux I__2160 (
            .O(N__9762),
            .I(N__9747));
    LocalMux I__2159 (
            .O(N__9757),
            .I(N__9747));
    InMux I__2158 (
            .O(N__9756),
            .I(N__9744));
    InMux I__2157 (
            .O(N__9755),
            .I(N__9735));
    InMux I__2156 (
            .O(N__9754),
            .I(N__9735));
    InMux I__2155 (
            .O(N__9753),
            .I(N__9735));
    InMux I__2154 (
            .O(N__9752),
            .I(N__9735));
    Span4Mux_h I__2153 (
            .O(N__9747),
            .I(N__9730));
    LocalMux I__2152 (
            .O(N__9744),
            .I(N__9730));
    LocalMux I__2151 (
            .O(N__9735),
            .I(N__9727));
    Span4Mux_v I__2150 (
            .O(N__9730),
            .I(N__9724));
    Span4Mux_v I__2149 (
            .O(N__9727),
            .I(N__9721));
    Span4Mux_v I__2148 (
            .O(N__9724),
            .I(N__9718));
    Sp12to4 I__2147 (
            .O(N__9721),
            .I(N__9715));
    Sp12to4 I__2146 (
            .O(N__9718),
            .I(N__9710));
    Span12Mux_h I__2145 (
            .O(N__9715),
            .I(N__9710));
    Odrv12 I__2144 (
            .O(N__9710),
            .I(A_c_1));
    CascadeMux I__2143 (
            .O(N__9707),
            .I(N__9703));
    CascadeMux I__2142 (
            .O(N__9706),
            .I(N__9699));
    InMux I__2141 (
            .O(N__9703),
            .I(N__9696));
    InMux I__2140 (
            .O(N__9702),
            .I(N__9691));
    InMux I__2139 (
            .O(N__9699),
            .I(N__9691));
    LocalMux I__2138 (
            .O(N__9696),
            .I(N__9688));
    LocalMux I__2137 (
            .O(N__9691),
            .I(N__9685));
    Span4Mux_v I__2136 (
            .O(N__9688),
            .I(N__9675));
    Span4Mux_v I__2135 (
            .O(N__9685),
            .I(N__9672));
    InMux I__2134 (
            .O(N__9684),
            .I(N__9669));
    InMux I__2133 (
            .O(N__9683),
            .I(N__9666));
    InMux I__2132 (
            .O(N__9682),
            .I(N__9663));
    InMux I__2131 (
            .O(N__9681),
            .I(N__9654));
    InMux I__2130 (
            .O(N__9680),
            .I(N__9654));
    InMux I__2129 (
            .O(N__9679),
            .I(N__9654));
    InMux I__2128 (
            .O(N__9678),
            .I(N__9654));
    Sp12to4 I__2127 (
            .O(N__9675),
            .I(N__9647));
    Sp12to4 I__2126 (
            .O(N__9672),
            .I(N__9647));
    LocalMux I__2125 (
            .O(N__9669),
            .I(N__9647));
    LocalMux I__2124 (
            .O(N__9666),
            .I(N__9640));
    LocalMux I__2123 (
            .O(N__9663),
            .I(N__9640));
    LocalMux I__2122 (
            .O(N__9654),
            .I(N__9640));
    Span12Mux_h I__2121 (
            .O(N__9647),
            .I(N__9637));
    Span12Mux_v I__2120 (
            .O(N__9640),
            .I(N__9634));
    Span12Mux_v I__2119 (
            .O(N__9637),
            .I(N__9629));
    Span12Mux_h I__2118 (
            .O(N__9634),
            .I(N__9629));
    Odrv12 I__2117 (
            .O(N__9629),
            .I(SIZ_c_1));
    CascadeMux I__2116 (
            .O(N__9626),
            .I(N__9618));
    CascadeMux I__2115 (
            .O(N__9625),
            .I(N__9615));
    InMux I__2114 (
            .O(N__9624),
            .I(N__9608));
    CascadeMux I__2113 (
            .O(N__9623),
            .I(N__9605));
    InMux I__2112 (
            .O(N__9622),
            .I(N__9596));
    InMux I__2111 (
            .O(N__9621),
            .I(N__9596));
    InMux I__2110 (
            .O(N__9618),
            .I(N__9596));
    InMux I__2109 (
            .O(N__9615),
            .I(N__9596));
    InMux I__2108 (
            .O(N__9614),
            .I(N__9593));
    InMux I__2107 (
            .O(N__9613),
            .I(N__9590));
    InMux I__2106 (
            .O(N__9612),
            .I(N__9585));
    InMux I__2105 (
            .O(N__9611),
            .I(N__9585));
    LocalMux I__2104 (
            .O(N__9608),
            .I(N__9582));
    InMux I__2103 (
            .O(N__9605),
            .I(N__9579));
    LocalMux I__2102 (
            .O(N__9596),
            .I(N__9576));
    LocalMux I__2101 (
            .O(N__9593),
            .I(N__9571));
    LocalMux I__2100 (
            .O(N__9590),
            .I(N__9571));
    LocalMux I__2099 (
            .O(N__9585),
            .I(N__9568));
    Span4Mux_v I__2098 (
            .O(N__9582),
            .I(N__9563));
    LocalMux I__2097 (
            .O(N__9579),
            .I(N__9563));
    Span4Mux_v I__2096 (
            .O(N__9576),
            .I(N__9558));
    Span4Mux_v I__2095 (
            .O(N__9571),
            .I(N__9558));
    Span4Mux_v I__2094 (
            .O(N__9568),
            .I(N__9555));
    Span4Mux_h I__2093 (
            .O(N__9563),
            .I(N__9552));
    Sp12to4 I__2092 (
            .O(N__9558),
            .I(N__9549));
    Span4Mux_v I__2091 (
            .O(N__9555),
            .I(N__9546));
    Span4Mux_v I__2090 (
            .O(N__9552),
            .I(N__9543));
    Span12Mux_h I__2089 (
            .O(N__9549),
            .I(N__9536));
    Sp12to4 I__2088 (
            .O(N__9546),
            .I(N__9536));
    Sp12to4 I__2087 (
            .O(N__9543),
            .I(N__9536));
    Odrv12 I__2086 (
            .O(N__9536),
            .I(A_c_0));
    CascadeMux I__2085 (
            .O(N__9533),
            .I(N__9529));
    InMux I__2084 (
            .O(N__9532),
            .I(N__9525));
    InMux I__2083 (
            .O(N__9529),
            .I(N__9522));
    CascadeMux I__2082 (
            .O(N__9528),
            .I(N__9516));
    LocalMux I__2081 (
            .O(N__9525),
            .I(N__9510));
    LocalMux I__2080 (
            .O(N__9522),
            .I(N__9510));
    CascadeMux I__2079 (
            .O(N__9521),
            .I(N__9507));
    CascadeMux I__2078 (
            .O(N__9520),
            .I(N__9504));
    InMux I__2077 (
            .O(N__9519),
            .I(N__9499));
    InMux I__2076 (
            .O(N__9516),
            .I(N__9494));
    InMux I__2075 (
            .O(N__9515),
            .I(N__9494));
    Span4Mux_v I__2074 (
            .O(N__9510),
            .I(N__9491));
    InMux I__2073 (
            .O(N__9507),
            .I(N__9482));
    InMux I__2072 (
            .O(N__9504),
            .I(N__9482));
    InMux I__2071 (
            .O(N__9503),
            .I(N__9482));
    InMux I__2070 (
            .O(N__9502),
            .I(N__9482));
    LocalMux I__2069 (
            .O(N__9499),
            .I(N__9479));
    LocalMux I__2068 (
            .O(N__9494),
            .I(N__9476));
    Span4Mux_v I__2067 (
            .O(N__9491),
            .I(N__9470));
    LocalMux I__2066 (
            .O(N__9482),
            .I(N__9470));
    Span4Mux_v I__2065 (
            .O(N__9479),
            .I(N__9467));
    Span4Mux_v I__2064 (
            .O(N__9476),
            .I(N__9464));
    InMux I__2063 (
            .O(N__9475),
            .I(N__9461));
    Span4Mux_h I__2062 (
            .O(N__9470),
            .I(N__9458));
    Sp12to4 I__2061 (
            .O(N__9467),
            .I(N__9451));
    Sp12to4 I__2060 (
            .O(N__9464),
            .I(N__9451));
    LocalMux I__2059 (
            .O(N__9461),
            .I(N__9451));
    Span4Mux_v I__2058 (
            .O(N__9458),
            .I(N__9448));
    Span12Mux_h I__2057 (
            .O(N__9451),
            .I(N__9445));
    Span4Mux_h I__2056 (
            .O(N__9448),
            .I(N__9442));
    Span12Mux_v I__2055 (
            .O(N__9445),
            .I(N__9439));
    Sp12to4 I__2054 (
            .O(N__9442),
            .I(N__9436));
    Odrv12 I__2053 (
            .O(N__9439),
            .I(SIZ_c_0));
    Odrv12 I__2052 (
            .O(N__9436),
            .I(SIZ_c_0));
    IoInMux I__2051 (
            .O(N__9431),
            .I(N__9428));
    LocalMux I__2050 (
            .O(N__9428),
            .I(N__9425));
    Span4Mux_s2_v I__2049 (
            .O(N__9425),
            .I(N__9422));
    Span4Mux_h I__2048 (
            .O(N__9422),
            .I(N__9419));
    Span4Mux_v I__2047 (
            .O(N__9419),
            .I(N__9416));
    Odrv4 I__2046 (
            .O(N__9416),
            .I(N_324_i));
    IoInMux I__2045 (
            .O(N__9413),
            .I(N__9410));
    LocalMux I__2044 (
            .O(N__9410),
            .I(N__9407));
    Span4Mux_s2_h I__2043 (
            .O(N__9407),
            .I(N__9404));
    Span4Mux_v I__2042 (
            .O(N__9404),
            .I(N__9401));
    Sp12to4 I__2041 (
            .O(N__9401),
            .I(N__9398));
    Span12Mux_h I__2040 (
            .O(N__9398),
            .I(N__9395));
    Odrv12 I__2039 (
            .O(N__9395),
            .I(WEn_c));
    InMux I__2038 (
            .O(N__9392),
            .I(N__9379));
    InMux I__2037 (
            .O(N__9391),
            .I(N__9379));
    InMux I__2036 (
            .O(N__9390),
            .I(N__9379));
    InMux I__2035 (
            .O(N__9389),
            .I(N__9376));
    InMux I__2034 (
            .O(N__9388),
            .I(N__9369));
    InMux I__2033 (
            .O(N__9387),
            .I(N__9369));
    InMux I__2032 (
            .O(N__9386),
            .I(N__9369));
    LocalMux I__2031 (
            .O(N__9379),
            .I(N__9365));
    LocalMux I__2030 (
            .O(N__9376),
            .I(N__9360));
    LocalMux I__2029 (
            .O(N__9369),
            .I(N__9360));
    InMux I__2028 (
            .O(N__9368),
            .I(N__9356));
    Span4Mux_h I__2027 (
            .O(N__9365),
            .I(N__9352));
    Span4Mux_h I__2026 (
            .O(N__9360),
            .I(N__9349));
    InMux I__2025 (
            .O(N__9359),
            .I(N__9346));
    LocalMux I__2024 (
            .O(N__9356),
            .I(N__9343));
    InMux I__2023 (
            .O(N__9355),
            .I(N__9340));
    Odrv4 I__2022 (
            .O(N__9352),
            .I(\U712_CHIP_RAM.N_305 ));
    Odrv4 I__2021 (
            .O(N__9349),
            .I(\U712_CHIP_RAM.N_305 ));
    LocalMux I__2020 (
            .O(N__9346),
            .I(\U712_CHIP_RAM.N_305 ));
    Odrv4 I__2019 (
            .O(N__9343),
            .I(\U712_CHIP_RAM.N_305 ));
    LocalMux I__2018 (
            .O(N__9340),
            .I(\U712_CHIP_RAM.N_305 ));
    CascadeMux I__2017 (
            .O(N__9329),
            .I(N__9321));
    CascadeMux I__2016 (
            .O(N__9328),
            .I(N__9318));
    CascadeMux I__2015 (
            .O(N__9327),
            .I(N__9315));
    CascadeMux I__2014 (
            .O(N__9326),
            .I(N__9312));
    CascadeMux I__2013 (
            .O(N__9325),
            .I(N__9308));
    CascadeMux I__2012 (
            .O(N__9324),
            .I(N__9305));
    InMux I__2011 (
            .O(N__9321),
            .I(N__9302));
    InMux I__2010 (
            .O(N__9318),
            .I(N__9297));
    InMux I__2009 (
            .O(N__9315),
            .I(N__9297));
    InMux I__2008 (
            .O(N__9312),
            .I(N__9292));
    InMux I__2007 (
            .O(N__9311),
            .I(N__9292));
    InMux I__2006 (
            .O(N__9308),
            .I(N__9289));
    InMux I__2005 (
            .O(N__9305),
            .I(N__9286));
    LocalMux I__2004 (
            .O(N__9302),
            .I(N__9283));
    LocalMux I__2003 (
            .O(N__9297),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__2002 (
            .O(N__9292),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__2001 (
            .O(N__9289),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__2000 (
            .O(N__9286),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    Odrv4 I__1999 (
            .O(N__9283),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    IoInMux I__1998 (
            .O(N__9272),
            .I(N__9269));
    LocalMux I__1997 (
            .O(N__9269),
            .I(N__9266));
    IoSpan4Mux I__1996 (
            .O(N__9266),
            .I(N__9263));
    Sp12to4 I__1995 (
            .O(N__9263),
            .I(N__9260));
    Span12Mux_s1_h I__1994 (
            .O(N__9260),
            .I(N__9257));
    Span12Mux_h I__1993 (
            .O(N__9257),
            .I(N__9254));
    Odrv12 I__1992 (
            .O(N__9254),
            .I(CMA_c_3));
    CEMux I__1991 (
            .O(N__9251),
            .I(N__9246));
    CEMux I__1990 (
            .O(N__9250),
            .I(N__9241));
    CEMux I__1989 (
            .O(N__9249),
            .I(N__9237));
    LocalMux I__1988 (
            .O(N__9246),
            .I(N__9234));
    CEMux I__1987 (
            .O(N__9245),
            .I(N__9230));
    CEMux I__1986 (
            .O(N__9244),
            .I(N__9227));
    LocalMux I__1985 (
            .O(N__9241),
            .I(N__9224));
    CEMux I__1984 (
            .O(N__9240),
            .I(N__9221));
    LocalMux I__1983 (
            .O(N__9237),
            .I(N__9216));
    Span4Mux_v I__1982 (
            .O(N__9234),
            .I(N__9216));
    CEMux I__1981 (
            .O(N__9233),
            .I(N__9213));
    LocalMux I__1980 (
            .O(N__9230),
            .I(N__9210));
    LocalMux I__1979 (
            .O(N__9227),
            .I(N__9207));
    Span4Mux_v I__1978 (
            .O(N__9224),
            .I(N__9204));
    LocalMux I__1977 (
            .O(N__9221),
            .I(N__9199));
    Span4Mux_h I__1976 (
            .O(N__9216),
            .I(N__9199));
    LocalMux I__1975 (
            .O(N__9213),
            .I(N__9196));
    Sp12to4 I__1974 (
            .O(N__9210),
            .I(N__9193));
    Span4Mux_h I__1973 (
            .O(N__9207),
            .I(N__9190));
    Odrv4 I__1972 (
            .O(N__9204),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv4 I__1971 (
            .O(N__9199),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv4 I__1970 (
            .O(N__9196),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv12 I__1969 (
            .O(N__9193),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv4 I__1968 (
            .O(N__9190),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    InMux I__1967 (
            .O(N__9179),
            .I(N__9175));
    InMux I__1966 (
            .O(N__9178),
            .I(N__9172));
    LocalMux I__1965 (
            .O(N__9175),
            .I(N__9169));
    LocalMux I__1964 (
            .O(N__9172),
            .I(N__9166));
    Span4Mux_h I__1963 (
            .O(N__9169),
            .I(N__9160));
    Span4Mux_h I__1962 (
            .O(N__9166),
            .I(N__9157));
    InMux I__1961 (
            .O(N__9165),
            .I(N__9154));
    InMux I__1960 (
            .O(N__9164),
            .I(N__9149));
    InMux I__1959 (
            .O(N__9163),
            .I(N__9149));
    Odrv4 I__1958 (
            .O(N__9160),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1957 (
            .O(N__9157),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1956 (
            .O(N__9154),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1955 (
            .O(N__9149),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    InMux I__1954 (
            .O(N__9140),
            .I(N__9137));
    LocalMux I__1953 (
            .O(N__9137),
            .I(\U712_CHIP_RAM.CMA_5_i_0_9 ));
    InMux I__1952 (
            .O(N__9134),
            .I(N__9131));
    LocalMux I__1951 (
            .O(N__9131),
            .I(N__9128));
    Odrv12 I__1950 (
            .O(N__9128),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    CascadeMux I__1949 (
            .O(N__9125),
            .I(N__9116));
    CascadeMux I__1948 (
            .O(N__9124),
            .I(N__9112));
    CascadeMux I__1947 (
            .O(N__9123),
            .I(N__9109));
    InMux I__1946 (
            .O(N__9122),
            .I(N__9105));
    InMux I__1945 (
            .O(N__9121),
            .I(N__9098));
    InMux I__1944 (
            .O(N__9120),
            .I(N__9098));
    InMux I__1943 (
            .O(N__9119),
            .I(N__9098));
    InMux I__1942 (
            .O(N__9116),
            .I(N__9095));
    InMux I__1941 (
            .O(N__9115),
            .I(N__9092));
    InMux I__1940 (
            .O(N__9112),
            .I(N__9089));
    InMux I__1939 (
            .O(N__9109),
            .I(N__9086));
    InMux I__1938 (
            .O(N__9108),
            .I(N__9076));
    LocalMux I__1937 (
            .O(N__9105),
            .I(N__9070));
    LocalMux I__1936 (
            .O(N__9098),
            .I(N__9067));
    LocalMux I__1935 (
            .O(N__9095),
            .I(N__9058));
    LocalMux I__1934 (
            .O(N__9092),
            .I(N__9058));
    LocalMux I__1933 (
            .O(N__9089),
            .I(N__9058));
    LocalMux I__1932 (
            .O(N__9086),
            .I(N__9058));
    InMux I__1931 (
            .O(N__9085),
            .I(N__9055));
    InMux I__1930 (
            .O(N__9084),
            .I(N__9052));
    InMux I__1929 (
            .O(N__9083),
            .I(N__9049));
    InMux I__1928 (
            .O(N__9082),
            .I(N__9044));
    InMux I__1927 (
            .O(N__9081),
            .I(N__9044));
    InMux I__1926 (
            .O(N__9080),
            .I(N__9039));
    InMux I__1925 (
            .O(N__9079),
            .I(N__9039));
    LocalMux I__1924 (
            .O(N__9076),
            .I(N__9036));
    InMux I__1923 (
            .O(N__9075),
            .I(N__9032));
    InMux I__1922 (
            .O(N__9074),
            .I(N__9027));
    InMux I__1921 (
            .O(N__9073),
            .I(N__9027));
    Span4Mux_h I__1920 (
            .O(N__9070),
            .I(N__9024));
    Span4Mux_h I__1919 (
            .O(N__9067),
            .I(N__9021));
    Span4Mux_h I__1918 (
            .O(N__9058),
            .I(N__9018));
    LocalMux I__1917 (
            .O(N__9055),
            .I(N__9015));
    LocalMux I__1916 (
            .O(N__9052),
            .I(N__9008));
    LocalMux I__1915 (
            .O(N__9049),
            .I(N__9008));
    LocalMux I__1914 (
            .O(N__9044),
            .I(N__9008));
    LocalMux I__1913 (
            .O(N__9039),
            .I(N__9003));
    Span4Mux_v I__1912 (
            .O(N__9036),
            .I(N__9003));
    CascadeMux I__1911 (
            .O(N__9035),
            .I(N__8999));
    LocalMux I__1910 (
            .O(N__9032),
            .I(N__8994));
    LocalMux I__1909 (
            .O(N__9027),
            .I(N__8991));
    Span4Mux_h I__1908 (
            .O(N__9024),
            .I(N__8986));
    Span4Mux_h I__1907 (
            .O(N__9021),
            .I(N__8986));
    Span4Mux_h I__1906 (
            .O(N__9018),
            .I(N__8983));
    Span4Mux_v I__1905 (
            .O(N__9015),
            .I(N__8976));
    Span4Mux_v I__1904 (
            .O(N__9008),
            .I(N__8976));
    Span4Mux_h I__1903 (
            .O(N__9003),
            .I(N__8976));
    InMux I__1902 (
            .O(N__9002),
            .I(N__8969));
    InMux I__1901 (
            .O(N__8999),
            .I(N__8969));
    InMux I__1900 (
            .O(N__8998),
            .I(N__8969));
    InMux I__1899 (
            .O(N__8997),
            .I(N__8966));
    Odrv4 I__1898 (
            .O(N__8994),
            .I(CPU_CYCLEm));
    Odrv4 I__1897 (
            .O(N__8991),
            .I(CPU_CYCLEm));
    Odrv4 I__1896 (
            .O(N__8986),
            .I(CPU_CYCLEm));
    Odrv4 I__1895 (
            .O(N__8983),
            .I(CPU_CYCLEm));
    Odrv4 I__1894 (
            .O(N__8976),
            .I(CPU_CYCLEm));
    LocalMux I__1893 (
            .O(N__8969),
            .I(CPU_CYCLEm));
    LocalMux I__1892 (
            .O(N__8966),
            .I(CPU_CYCLEm));
    InMux I__1891 (
            .O(N__8951),
            .I(N__8948));
    LocalMux I__1890 (
            .O(N__8948),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    InMux I__1889 (
            .O(N__8945),
            .I(N__8942));
    LocalMux I__1888 (
            .O(N__8942),
            .I(N__8939));
    Odrv4 I__1887 (
            .O(N__8939),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__1886 (
            .O(N__8936),
            .I(N__8932));
    InMux I__1885 (
            .O(N__8935),
            .I(N__8929));
    LocalMux I__1884 (
            .O(N__8932),
            .I(\U712_REG_SM.START_RSTZ0 ));
    LocalMux I__1883 (
            .O(N__8929),
            .I(\U712_REG_SM.START_RSTZ0 ));
    InMux I__1882 (
            .O(N__8924),
            .I(N__8921));
    LocalMux I__1881 (
            .O(N__8921),
            .I(N__8918));
    Odrv12 I__1880 (
            .O(N__8918),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_7 ));
    InMux I__1879 (
            .O(N__8915),
            .I(N__8910));
    InMux I__1878 (
            .O(N__8914),
            .I(N__8907));
    InMux I__1877 (
            .O(N__8913),
            .I(N__8904));
    LocalMux I__1876 (
            .O(N__8910),
            .I(\U712_REG_SM.N_319 ));
    LocalMux I__1875 (
            .O(N__8907),
            .I(\U712_REG_SM.N_319 ));
    LocalMux I__1874 (
            .O(N__8904),
            .I(\U712_REG_SM.N_319 ));
    InMux I__1873 (
            .O(N__8897),
            .I(N__8893));
    InMux I__1872 (
            .O(N__8896),
            .I(N__8890));
    LocalMux I__1871 (
            .O(N__8893),
            .I(N__8885));
    LocalMux I__1870 (
            .O(N__8890),
            .I(N__8882));
    InMux I__1869 (
            .O(N__8889),
            .I(N__8879));
    InMux I__1868 (
            .O(N__8888),
            .I(N__8876));
    Span4Mux_h I__1867 (
            .O(N__8885),
            .I(N__8873));
    Odrv4 I__1866 (
            .O(N__8882),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__1865 (
            .O(N__8879),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__1864 (
            .O(N__8876),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    Odrv4 I__1863 (
            .O(N__8873),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    CascadeMux I__1862 (
            .O(N__8864),
            .I(\U712_REG_SM.N_318_cascade_ ));
    InMux I__1861 (
            .O(N__8861),
            .I(N__8855));
    InMux I__1860 (
            .O(N__8860),
            .I(N__8850));
    InMux I__1859 (
            .O(N__8859),
            .I(N__8850));
    InMux I__1858 (
            .O(N__8858),
            .I(N__8847));
    LocalMux I__1857 (
            .O(N__8855),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1856 (
            .O(N__8850),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1855 (
            .O(N__8847),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    IoInMux I__1854 (
            .O(N__8840),
            .I(N__8837));
    LocalMux I__1853 (
            .O(N__8837),
            .I(N__8834));
    Span4Mux_s0_v I__1852 (
            .O(N__8834),
            .I(N__8831));
    Span4Mux_v I__1851 (
            .O(N__8831),
            .I(N__8827));
    IoInMux I__1850 (
            .O(N__8830),
            .I(N__8824));
    Span4Mux_v I__1849 (
            .O(N__8827),
            .I(N__8821));
    LocalMux I__1848 (
            .O(N__8824),
            .I(N__8818));
    Sp12to4 I__1847 (
            .O(N__8821),
            .I(N__8815));
    Span12Mux_s8_v I__1846 (
            .O(N__8818),
            .I(N__8812));
    Span12Mux_h I__1845 (
            .O(N__8815),
            .I(N__8805));
    Span12Mux_h I__1844 (
            .O(N__8812),
            .I(N__8805));
    InMux I__1843 (
            .O(N__8811),
            .I(N__8802));
    InMux I__1842 (
            .O(N__8810),
            .I(N__8799));
    Odrv12 I__1841 (
            .O(N__8805),
            .I(BLSn_c));
    LocalMux I__1840 (
            .O(N__8802),
            .I(BLSn_c));
    LocalMux I__1839 (
            .O(N__8799),
            .I(BLSn_c));
    InMux I__1838 (
            .O(N__8792),
            .I(N__8789));
    LocalMux I__1837 (
            .O(N__8789),
            .I(\U712_REG_SM.REGENn_e_1 ));
    IoInMux I__1836 (
            .O(N__8786),
            .I(N__8783));
    LocalMux I__1835 (
            .O(N__8783),
            .I(N__8780));
    Span4Mux_s0_v I__1834 (
            .O(N__8780),
            .I(N__8777));
    Span4Mux_v I__1833 (
            .O(N__8777),
            .I(N__8774));
    Odrv4 I__1832 (
            .O(N__8774),
            .I(N_326_i));
    InMux I__1831 (
            .O(N__8771),
            .I(N__8768));
    LocalMux I__1830 (
            .O(N__8768),
            .I(N__8765));
    Span4Mux_v I__1829 (
            .O(N__8765),
            .I(N__8762));
    Span4Mux_v I__1828 (
            .O(N__8762),
            .I(N__8759));
    Sp12to4 I__1827 (
            .O(N__8759),
            .I(N__8756));
    Span12Mux_h I__1826 (
            .O(N__8756),
            .I(N__8753));
    Odrv12 I__1825 (
            .O(N__8753),
            .I(A_c_19));
    IoInMux I__1824 (
            .O(N__8750),
            .I(N__8747));
    LocalMux I__1823 (
            .O(N__8747),
            .I(N__8744));
    IoSpan4Mux I__1822 (
            .O(N__8744),
            .I(N__8741));
    Span4Mux_s0_h I__1821 (
            .O(N__8741),
            .I(N__8738));
    Sp12to4 I__1820 (
            .O(N__8738),
            .I(N__8735));
    Span12Mux_h I__1819 (
            .O(N__8735),
            .I(N__8732));
    Odrv12 I__1818 (
            .O(N__8732),
            .I(CMA_c_9));
    InMux I__1817 (
            .O(N__8729),
            .I(N__8726));
    LocalMux I__1816 (
            .O(N__8726),
            .I(N__8723));
    Odrv4 I__1815 (
            .O(N__8723),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__1814 (
            .O(N__8720),
            .I(N__8717));
    LocalMux I__1813 (
            .O(N__8717),
            .I(N__8714));
    Odrv4 I__1812 (
            .O(N__8714),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1811 (
            .O(N__8711),
            .I(N__8708));
    LocalMux I__1810 (
            .O(N__8708),
            .I(N__8705));
    Odrv12 I__1809 (
            .O(N__8705),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__1808 (
            .O(N__8702),
            .I(N__8699));
    LocalMux I__1807 (
            .O(N__8699),
            .I(N__8696));
    Span4Mux_h I__1806 (
            .O(N__8696),
            .I(N__8693));
    Odrv4 I__1805 (
            .O(N__8693),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1804 (
            .O(N__8690),
            .I(N__8687));
    LocalMux I__1803 (
            .O(N__8687),
            .I(N__8684));
    Odrv4 I__1802 (
            .O(N__8684),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1801 (
            .O(N__8681),
            .I(N__8678));
    LocalMux I__1800 (
            .O(N__8678),
            .I(N__8675));
    Span4Mux_h I__1799 (
            .O(N__8675),
            .I(N__8672));
    Odrv4 I__1798 (
            .O(N__8672),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__1797 (
            .O(N__8669),
            .I(N__8661));
    InMux I__1796 (
            .O(N__8668),
            .I(N__8661));
    InMux I__1795 (
            .O(N__8667),
            .I(N__8658));
    InMux I__1794 (
            .O(N__8666),
            .I(N__8655));
    LocalMux I__1793 (
            .O(N__8661),
            .I(N__8652));
    LocalMux I__1792 (
            .O(N__8658),
            .I(N__8649));
    LocalMux I__1791 (
            .O(N__8655),
            .I(N__8646));
    Span4Mux_h I__1790 (
            .O(N__8652),
            .I(N__8643));
    Span4Mux_h I__1789 (
            .O(N__8649),
            .I(N__8640));
    Span12Mux_v I__1788 (
            .O(N__8646),
            .I(N__8637));
    Sp12to4 I__1787 (
            .O(N__8643),
            .I(N__8634));
    Span4Mux_v I__1786 (
            .O(N__8640),
            .I(N__8631));
    Span12Mux_h I__1785 (
            .O(N__8637),
            .I(N__8628));
    Span12Mux_v I__1784 (
            .O(N__8634),
            .I(N__8623));
    Sp12to4 I__1783 (
            .O(N__8631),
            .I(N__8623));
    Odrv12 I__1782 (
            .O(N__8628),
            .I(DRA_c_6));
    Odrv12 I__1781 (
            .O(N__8623),
            .I(DRA_c_6));
    InMux I__1780 (
            .O(N__8618),
            .I(N__8615));
    LocalMux I__1779 (
            .O(N__8615),
            .I(N__8612));
    Span4Mux_h I__1778 (
            .O(N__8612),
            .I(N__8609));
    Span4Mux_v I__1777 (
            .O(N__8609),
            .I(N__8606));
    Odrv4 I__1776 (
            .O(N__8606),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__1775 (
            .O(N__8603),
            .I(N__8599));
    IoInMux I__1774 (
            .O(N__8602),
            .I(N__8596));
    LocalMux I__1773 (
            .O(N__8599),
            .I(N__8593));
    LocalMux I__1772 (
            .O(N__8596),
            .I(N__8590));
    Span4Mux_v I__1771 (
            .O(N__8593),
            .I(N__8587));
    IoSpan4Mux I__1770 (
            .O(N__8590),
            .I(N__8584));
    Sp12to4 I__1769 (
            .O(N__8587),
            .I(N__8581));
    IoSpan4Mux I__1768 (
            .O(N__8584),
            .I(N__8578));
    Span12Mux_h I__1767 (
            .O(N__8581),
            .I(N__8575));
    IoSpan4Mux I__1766 (
            .O(N__8578),
            .I(N__8572));
    Odrv12 I__1765 (
            .O(N__8575),
            .I(C1_c));
    Odrv4 I__1764 (
            .O(N__8572),
            .I(C1_c));
    InMux I__1763 (
            .O(N__8567),
            .I(N__8564));
    LocalMux I__1762 (
            .O(N__8564),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__1761 (
            .O(N__8561),
            .I(N__8558));
    LocalMux I__1760 (
            .O(N__8558),
            .I(N__8555));
    Span4Mux_v I__1759 (
            .O(N__8555),
            .I(N__8552));
    Odrv4 I__1758 (
            .O(N__8552),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__1757 (
            .O(N__8549),
            .I(N__8546));
    LocalMux I__1756 (
            .O(N__8546),
            .I(N__8543));
    Span4Mux_s1_v I__1755 (
            .O(N__8543),
            .I(N__8540));
    Span4Mux_v I__1754 (
            .O(N__8540),
            .I(N__8537));
    Span4Mux_v I__1753 (
            .O(N__8537),
            .I(N__8534));
    Odrv4 I__1752 (
            .O(N__8534),
            .I(CMA_c_0));
    IoInMux I__1751 (
            .O(N__8531),
            .I(N__8528));
    LocalMux I__1750 (
            .O(N__8528),
            .I(N__8525));
    Span4Mux_s0_v I__1749 (
            .O(N__8525),
            .I(N__8522));
    Sp12to4 I__1748 (
            .O(N__8522),
            .I(N__8519));
    Span12Mux_h I__1747 (
            .O(N__8519),
            .I(N__8516));
    Odrv12 I__1746 (
            .O(N__8516),
            .I(CMA_c_10));
    InMux I__1745 (
            .O(N__8513),
            .I(N__8510));
    LocalMux I__1744 (
            .O(N__8510),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__1743 (
            .O(N__8507),
            .I(N__8504));
    LocalMux I__1742 (
            .O(N__8504),
            .I(N__8501));
    IoSpan4Mux I__1741 (
            .O(N__8501),
            .I(N__8498));
    IoSpan4Mux I__1740 (
            .O(N__8498),
            .I(N__8495));
    Span4Mux_s3_h I__1739 (
            .O(N__8495),
            .I(N__8492));
    Sp12to4 I__1738 (
            .O(N__8492),
            .I(N__8489));
    Odrv12 I__1737 (
            .O(N__8489),
            .I(CMA_c_6));
    InMux I__1736 (
            .O(N__8486),
            .I(N__8483));
    LocalMux I__1735 (
            .O(N__8483),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ));
    IoInMux I__1734 (
            .O(N__8480),
            .I(N__8477));
    LocalMux I__1733 (
            .O(N__8477),
            .I(N__8474));
    IoSpan4Mux I__1732 (
            .O(N__8474),
            .I(N__8471));
    Span4Mux_s2_h I__1731 (
            .O(N__8471),
            .I(N__8468));
    Span4Mux_v I__1730 (
            .O(N__8468),
            .I(N__8465));
    Span4Mux_h I__1729 (
            .O(N__8465),
            .I(N__8462));
    Span4Mux_h I__1728 (
            .O(N__8462),
            .I(N__8459));
    Odrv4 I__1727 (
            .O(N__8459),
            .I(CMA_c_8));
    InMux I__1726 (
            .O(N__8456),
            .I(N__8453));
    LocalMux I__1725 (
            .O(N__8453),
            .I(N__8450));
    Odrv4 I__1724 (
            .O(N__8450),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__1723 (
            .O(N__8447),
            .I(N__8444));
    LocalMux I__1722 (
            .O(N__8444),
            .I(N__8441));
    Span4Mux_s2_h I__1721 (
            .O(N__8441),
            .I(N__8438));
    Sp12to4 I__1720 (
            .O(N__8438),
            .I(N__8435));
    Span12Mux_s11_v I__1719 (
            .O(N__8435),
            .I(N__8432));
    Span12Mux_h I__1718 (
            .O(N__8432),
            .I(N__8429));
    Odrv12 I__1717 (
            .O(N__8429),
            .I(CMA_c_4));
    InMux I__1716 (
            .O(N__8426),
            .I(N__8423));
    LocalMux I__1715 (
            .O(N__8423),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1714 (
            .O(N__8420),
            .I(N__8417));
    LocalMux I__1713 (
            .O(N__8417),
            .I(N__8414));
    Span4Mux_s2_h I__1712 (
            .O(N__8414),
            .I(N__8411));
    Sp12to4 I__1711 (
            .O(N__8411),
            .I(N__8408));
    Span12Mux_s10_v I__1710 (
            .O(N__8408),
            .I(N__8405));
    Odrv12 I__1709 (
            .O(N__8405),
            .I(CMA_c_7));
    CascadeMux I__1708 (
            .O(N__8402),
            .I(\U712_REG_SM.REG_CYCLE_5_iv_0_0_cascade_ ));
    InMux I__1707 (
            .O(N__8399),
            .I(N__8396));
    LocalMux I__1706 (
            .O(N__8396),
            .I(\U712_REG_SM.N_409 ));
    InMux I__1705 (
            .O(N__8393),
            .I(N__8390));
    LocalMux I__1704 (
            .O(N__8390),
            .I(N__8387));
    Span4Mux_v I__1703 (
            .O(N__8387),
            .I(N__8383));
    InMux I__1702 (
            .O(N__8386),
            .I(N__8380));
    Span4Mux_h I__1701 (
            .O(N__8383),
            .I(N__8375));
    LocalMux I__1700 (
            .O(N__8380),
            .I(N__8372));
    InMux I__1699 (
            .O(N__8379),
            .I(N__8367));
    InMux I__1698 (
            .O(N__8378),
            .I(N__8367));
    Odrv4 I__1697 (
            .O(N__8375),
            .I(REG_CYCLEm));
    Odrv4 I__1696 (
            .O(N__8372),
            .I(REG_CYCLEm));
    LocalMux I__1695 (
            .O(N__8367),
            .I(REG_CYCLEm));
    InMux I__1694 (
            .O(N__8360),
            .I(N__8357));
    LocalMux I__1693 (
            .O(N__8357),
            .I(\U712_REG_SM.STATE_COUNTsr_0 ));
    CascadeMux I__1692 (
            .O(N__8354),
            .I(N__8351));
    InMux I__1691 (
            .O(N__8351),
            .I(N__8348));
    LocalMux I__1690 (
            .O(N__8348),
            .I(\U712_REG_SM.N_328 ));
    CascadeMux I__1689 (
            .O(N__8345),
            .I(N__8341));
    CascadeMux I__1688 (
            .O(N__8344),
            .I(N__8338));
    InMux I__1687 (
            .O(N__8341),
            .I(N__8335));
    InMux I__1686 (
            .O(N__8338),
            .I(N__8326));
    LocalMux I__1685 (
            .O(N__8335),
            .I(N__8323));
    InMux I__1684 (
            .O(N__8334),
            .I(N__8320));
    InMux I__1683 (
            .O(N__8333),
            .I(N__8311));
    InMux I__1682 (
            .O(N__8332),
            .I(N__8311));
    InMux I__1681 (
            .O(N__8331),
            .I(N__8311));
    InMux I__1680 (
            .O(N__8330),
            .I(N__8311));
    InMux I__1679 (
            .O(N__8329),
            .I(N__8308));
    LocalMux I__1678 (
            .O(N__8326),
            .I(N__8305));
    Span4Mux_h I__1677 (
            .O(N__8323),
            .I(N__8300));
    LocalMux I__1676 (
            .O(N__8320),
            .I(N__8300));
    LocalMux I__1675 (
            .O(N__8311),
            .I(N__8294));
    LocalMux I__1674 (
            .O(N__8308),
            .I(N__8294));
    Span4Mux_v I__1673 (
            .O(N__8305),
            .I(N__8289));
    Span4Mux_h I__1672 (
            .O(N__8300),
            .I(N__8289));
    InMux I__1671 (
            .O(N__8299),
            .I(N__8286));
    Odrv4 I__1670 (
            .O(N__8294),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1669 (
            .O(N__8289),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1668 (
            .O(N__8286),
            .I(DBR_SYNCZ0Z_1));
    CascadeMux I__1667 (
            .O(N__8279),
            .I(\U712_REG_SM.N_412_cascade_ ));
    InMux I__1666 (
            .O(N__8276),
            .I(N__8271));
    InMux I__1665 (
            .O(N__8275),
            .I(N__8266));
    InMux I__1664 (
            .O(N__8274),
            .I(N__8266));
    LocalMux I__1663 (
            .O(N__8271),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_3 ));
    LocalMux I__1662 (
            .O(N__8266),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_3 ));
    CascadeMux I__1661 (
            .O(N__8261),
            .I(\U712_REG_SM.N_360_cascade_ ));
    InMux I__1660 (
            .O(N__8258),
            .I(N__8255));
    LocalMux I__1659 (
            .O(N__8255),
            .I(\U712_REG_SM.N_320 ));
    InMux I__1658 (
            .O(N__8252),
            .I(N__8245));
    InMux I__1657 (
            .O(N__8251),
            .I(N__8245));
    InMux I__1656 (
            .O(N__8250),
            .I(N__8242));
    LocalMux I__1655 (
            .O(N__8245),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__1654 (
            .O(N__8242),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    IoInMux I__1653 (
            .O(N__8237),
            .I(N__8234));
    LocalMux I__1652 (
            .O(N__8234),
            .I(N__8231));
    IoSpan4Mux I__1651 (
            .O(N__8231),
            .I(N__8228));
    Span4Mux_s3_h I__1650 (
            .O(N__8228),
            .I(N__8225));
    Span4Mux_v I__1649 (
            .O(N__8225),
            .I(N__8221));
    InMux I__1648 (
            .O(N__8224),
            .I(N__8218));
    Span4Mux_h I__1647 (
            .O(N__8221),
            .I(N__8215));
    LocalMux I__1646 (
            .O(N__8218),
            .I(N__8212));
    Sp12to4 I__1645 (
            .O(N__8215),
            .I(N__8209));
    Span4Mux_v I__1644 (
            .O(N__8212),
            .I(N__8206));
    Span12Mux_h I__1643 (
            .O(N__8209),
            .I(N__8201));
    Sp12to4 I__1642 (
            .O(N__8206),
            .I(N__8201));
    Span12Mux_h I__1641 (
            .O(N__8201),
            .I(N__8198));
    Odrv12 I__1640 (
            .O(N__8198),
            .I(C3_c));
    InMux I__1639 (
            .O(N__8195),
            .I(N__8192));
    LocalMux I__1638 (
            .O(N__8192),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__1637 (
            .O(N__8189),
            .I(N__8186));
    LocalMux I__1636 (
            .O(N__8186),
            .I(\U712_CHIP_RAM.N_346 ));
    InMux I__1635 (
            .O(N__8183),
            .I(N__8180));
    LocalMux I__1634 (
            .O(N__8180),
            .I(\U712_CHIP_RAM.N_352 ));
    IoInMux I__1633 (
            .O(N__8177),
            .I(N__8174));
    LocalMux I__1632 (
            .O(N__8174),
            .I(N__8171));
    IoSpan4Mux I__1631 (
            .O(N__8171),
            .I(N__8168));
    Sp12to4 I__1630 (
            .O(N__8168),
            .I(N__8165));
    Span12Mux_s7_h I__1629 (
            .O(N__8165),
            .I(N__8162));
    Span12Mux_v I__1628 (
            .O(N__8162),
            .I(N__8159));
    Odrv12 I__1627 (
            .O(N__8159),
            .I(CMA_c_5));
    InMux I__1626 (
            .O(N__8156),
            .I(N__8152));
    InMux I__1625 (
            .O(N__8155),
            .I(N__8149));
    LocalMux I__1624 (
            .O(N__8152),
            .I(N__8146));
    LocalMux I__1623 (
            .O(N__8149),
            .I(N__8143));
    Span4Mux_h I__1622 (
            .O(N__8146),
            .I(N__8140));
    Span4Mux_v I__1621 (
            .O(N__8143),
            .I(N__8137));
    Span4Mux_v I__1620 (
            .O(N__8140),
            .I(N__8134));
    Span4Mux_h I__1619 (
            .O(N__8137),
            .I(N__8131));
    Odrv4 I__1618 (
            .O(N__8134),
            .I(DBRn_c_i));
    Odrv4 I__1617 (
            .O(N__8131),
            .I(DBRn_c_i));
    InMux I__1616 (
            .O(N__8126),
            .I(N__8122));
    InMux I__1615 (
            .O(N__8125),
            .I(N__8119));
    LocalMux I__1614 (
            .O(N__8122),
            .I(N__8116));
    LocalMux I__1613 (
            .O(N__8119),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    Odrv4 I__1612 (
            .O(N__8116),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    IoInMux I__1611 (
            .O(N__8111),
            .I(N__8108));
    LocalMux I__1610 (
            .O(N__8108),
            .I(N__8105));
    Span4Mux_s0_v I__1609 (
            .O(N__8105),
            .I(N__8102));
    Span4Mux_v I__1608 (
            .O(N__8102),
            .I(N__8099));
    Span4Mux_v I__1607 (
            .O(N__8099),
            .I(N__8096));
    Sp12to4 I__1606 (
            .O(N__8096),
            .I(N__8093));
    Span12Mux_h I__1605 (
            .O(N__8093),
            .I(N__8090));
    Odrv12 I__1604 (
            .O(N__8090),
            .I(N_169_i));
    InMux I__1603 (
            .O(N__8087),
            .I(N__8084));
    LocalMux I__1602 (
            .O(N__8084),
            .I(N__8081));
    Span4Mux_v I__1601 (
            .O(N__8081),
            .I(N__8078));
    Span4Mux_v I__1600 (
            .O(N__8078),
            .I(N__8075));
    Span4Mux_v I__1599 (
            .O(N__8075),
            .I(N__8072));
    Sp12to4 I__1598 (
            .O(N__8072),
            .I(N__8069));
    Span12Mux_h I__1597 (
            .O(N__8069),
            .I(N__8066));
    Odrv12 I__1596 (
            .O(N__8066),
            .I(REGSPACEn_c));
    CascadeMux I__1595 (
            .O(N__8063),
            .I(\U712_REG_SM.N_397_cascade_ ));
    InMux I__1594 (
            .O(N__8060),
            .I(N__8057));
    LocalMux I__1593 (
            .O(N__8057),
            .I(N__8054));
    Span4Mux_v I__1592 (
            .O(N__8054),
            .I(N__8050));
    InMux I__1591 (
            .O(N__8053),
            .I(N__8047));
    Sp12to4 I__1590 (
            .O(N__8050),
            .I(N__8044));
    LocalMux I__1589 (
            .O(N__8047),
            .I(N__8041));
    Span12Mux_h I__1588 (
            .O(N__8044),
            .I(N__8038));
    Span12Mux_h I__1587 (
            .O(N__8041),
            .I(N__8035));
    Span12Mux_v I__1586 (
            .O(N__8038),
            .I(N__8032));
    Span12Mux_v I__1585 (
            .O(N__8035),
            .I(N__8029));
    Odrv12 I__1584 (
            .O(N__8032),
            .I(TSn_c));
    Odrv12 I__1583 (
            .O(N__8029),
            .I(TSn_c));
    InMux I__1582 (
            .O(N__8024),
            .I(N__8021));
    LocalMux I__1581 (
            .O(N__8021),
            .I(N__8018));
    Odrv12 I__1580 (
            .O(N__8018),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ));
    InMux I__1579 (
            .O(N__8015),
            .I(N__8011));
    InMux I__1578 (
            .O(N__8014),
            .I(N__8008));
    LocalMux I__1577 (
            .O(N__8011),
            .I(\U712_REG_SM.N_548 ));
    LocalMux I__1576 (
            .O(N__8008),
            .I(\U712_REG_SM.N_548 ));
    CascadeMux I__1575 (
            .O(N__8003),
            .I(\U712_REG_SM.N_319_cascade_ ));
    CascadeMux I__1574 (
            .O(N__8000),
            .I(\U712_REG_SM.N_320_cascade_ ));
    IoInMux I__1573 (
            .O(N__7997),
            .I(N__7994));
    LocalMux I__1572 (
            .O(N__7994),
            .I(N__7991));
    Span12Mux_s1_v I__1571 (
            .O(N__7991),
            .I(N__7988));
    Odrv12 I__1570 (
            .O(N__7988),
            .I(RESETn_c_i));
    InMux I__1569 (
            .O(N__7985),
            .I(N__7982));
    LocalMux I__1568 (
            .O(N__7982),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    CascadeMux I__1567 (
            .O(N__7979),
            .I(N__7976));
    InMux I__1566 (
            .O(N__7976),
            .I(N__7973));
    LocalMux I__1565 (
            .O(N__7973),
            .I(N__7970));
    Span4Mux_h I__1564 (
            .O(N__7970),
            .I(N__7967));
    Odrv4 I__1563 (
            .O(N__7967),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__1562 (
            .O(N__7964),
            .I(N__7961));
    LocalMux I__1561 (
            .O(N__7961),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i ));
    InMux I__1560 (
            .O(N__7958),
            .I(N__7955));
    LocalMux I__1559 (
            .O(N__7955),
            .I(N__7952));
    Odrv4 I__1558 (
            .O(N__7952),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8 ));
    InMux I__1557 (
            .O(N__7949),
            .I(N__7946));
    LocalMux I__1556 (
            .O(N__7946),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ));
    CascadeMux I__1555 (
            .O(N__7943),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ));
    InMux I__1554 (
            .O(N__7940),
            .I(N__7937));
    LocalMux I__1553 (
            .O(N__7937),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    IoInMux I__1552 (
            .O(N__7934),
            .I(N__7931));
    LocalMux I__1551 (
            .O(N__7931),
            .I(N__7928));
    Span4Mux_s3_v I__1550 (
            .O(N__7928),
            .I(N__7925));
    Span4Mux_v I__1549 (
            .O(N__7925),
            .I(N__7922));
    Span4Mux_v I__1548 (
            .O(N__7922),
            .I(N__7919));
    Odrv4 I__1547 (
            .O(N__7919),
            .I(CMA_c_1));
    InMux I__1546 (
            .O(N__7916),
            .I(N__7913));
    LocalMux I__1545 (
            .O(N__7913),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    InMux I__1544 (
            .O(N__7910),
            .I(N__7902));
    InMux I__1543 (
            .O(N__7909),
            .I(N__7902));
    InMux I__1542 (
            .O(N__7908),
            .I(N__7897));
    InMux I__1541 (
            .O(N__7907),
            .I(N__7897));
    LocalMux I__1540 (
            .O(N__7902),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1539 (
            .O(N__7897),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__1538 (
            .O(N__7892),
            .I(N__7889));
    LocalMux I__1537 (
            .O(N__7889),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ));
    CascadeMux I__1536 (
            .O(N__7886),
            .I(N__7883));
    InMux I__1535 (
            .O(N__7883),
            .I(N__7880));
    LocalMux I__1534 (
            .O(N__7880),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    InMux I__1533 (
            .O(N__7877),
            .I(N__7873));
    InMux I__1532 (
            .O(N__7876),
            .I(N__7870));
    LocalMux I__1531 (
            .O(N__7873),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__1530 (
            .O(N__7870),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__1529 (
            .O(N__7865),
            .I(N__7861));
    InMux I__1528 (
            .O(N__7864),
            .I(N__7855));
    InMux I__1527 (
            .O(N__7861),
            .I(N__7855));
    InMux I__1526 (
            .O(N__7860),
            .I(N__7852));
    LocalMux I__1525 (
            .O(N__7855),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__1524 (
            .O(N__7852),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__1523 (
            .O(N__7847),
            .I(N__7841));
    InMux I__1522 (
            .O(N__7846),
            .I(N__7836));
    InMux I__1521 (
            .O(N__7845),
            .I(N__7836));
    InMux I__1520 (
            .O(N__7844),
            .I(N__7833));
    LocalMux I__1519 (
            .O(N__7841),
            .I(REG_TACK));
    LocalMux I__1518 (
            .O(N__7836),
            .I(REG_TACK));
    LocalMux I__1517 (
            .O(N__7833),
            .I(REG_TACK));
    InMux I__1516 (
            .O(N__7826),
            .I(N__7823));
    LocalMux I__1515 (
            .O(N__7823),
            .I(\U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1 ));
    InMux I__1514 (
            .O(N__7820),
            .I(N__7814));
    InMux I__1513 (
            .O(N__7819),
            .I(N__7814));
    LocalMux I__1512 (
            .O(N__7814),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_5 ));
    InMux I__1511 (
            .O(N__7811),
            .I(N__7808));
    LocalMux I__1510 (
            .O(N__7808),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_6 ));
    InMux I__1509 (
            .O(N__7805),
            .I(N__7802));
    LocalMux I__1508 (
            .O(N__7802),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_4 ));
    InMux I__1507 (
            .O(N__7799),
            .I(N__7795));
    InMux I__1506 (
            .O(N__7798),
            .I(N__7792));
    LocalMux I__1505 (
            .O(N__7795),
            .I(N__7789));
    LocalMux I__1504 (
            .O(N__7792),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0 ));
    Odrv12 I__1503 (
            .O(N__7789),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0 ));
    CascadeMux I__1502 (
            .O(N__7784),
            .I(N__7781));
    InMux I__1501 (
            .O(N__7781),
            .I(N__7778));
    LocalMux I__1500 (
            .O(N__7778),
            .I(N__7775));
    Span4Mux_v I__1499 (
            .O(N__7775),
            .I(N__7772));
    Odrv4 I__1498 (
            .O(N__7772),
            .I(\U712_BYTE_ENABLE.N_325 ));
    IoInMux I__1497 (
            .O(N__7769),
            .I(N__7766));
    LocalMux I__1496 (
            .O(N__7766),
            .I(N__7763));
    Span12Mux_s10_h I__1495 (
            .O(N__7763),
            .I(N__7760));
    Span12Mux_v I__1494 (
            .O(N__7760),
            .I(N__7757));
    Odrv12 I__1493 (
            .O(N__7757),
            .I(N_186_i));
    InMux I__1492 (
            .O(N__7754),
            .I(N__7748));
    InMux I__1491 (
            .O(N__7753),
            .I(N__7745));
    InMux I__1490 (
            .O(N__7752),
            .I(N__7740));
    InMux I__1489 (
            .O(N__7751),
            .I(N__7740));
    LocalMux I__1488 (
            .O(N__7748),
            .I(CPU_TACKm));
    LocalMux I__1487 (
            .O(N__7745),
            .I(CPU_TACKm));
    LocalMux I__1486 (
            .O(N__7740),
            .I(CPU_TACKm));
    CascadeMux I__1485 (
            .O(N__7733),
            .I(\U712_CYCLE_TERM.N_450_cascade_ ));
    CascadeMux I__1484 (
            .O(N__7730),
            .I(N__7727));
    InMux I__1483 (
            .O(N__7727),
            .I(N__7721));
    InMux I__1482 (
            .O(N__7726),
            .I(N__7721));
    LocalMux I__1481 (
            .O(N__7721),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    InMux I__1480 (
            .O(N__7718),
            .I(N__7715));
    LocalMux I__1479 (
            .O(N__7715),
            .I(N__7711));
    CascadeMux I__1478 (
            .O(N__7714),
            .I(N__7706));
    Span4Mux_v I__1477 (
            .O(N__7711),
            .I(N__7703));
    InMux I__1476 (
            .O(N__7710),
            .I(N__7698));
    InMux I__1475 (
            .O(N__7709),
            .I(N__7698));
    InMux I__1474 (
            .O(N__7706),
            .I(N__7695));
    Span4Mux_v I__1473 (
            .O(N__7703),
            .I(N__7692));
    LocalMux I__1472 (
            .O(N__7698),
            .I(N__7689));
    LocalMux I__1471 (
            .O(N__7695),
            .I(N__7686));
    Sp12to4 I__1470 (
            .O(N__7692),
            .I(N__7683));
    Sp12to4 I__1469 (
            .O(N__7689),
            .I(N__7678));
    Sp12to4 I__1468 (
            .O(N__7686),
            .I(N__7678));
    Span12Mux_h I__1467 (
            .O(N__7683),
            .I(N__7673));
    Span12Mux_v I__1466 (
            .O(N__7678),
            .I(N__7673));
    Odrv12 I__1465 (
            .O(N__7673),
            .I(CLK40_PLL_i));
    CascadeMux I__1464 (
            .O(N__7670),
            .I(N__7666));
    InMux I__1463 (
            .O(N__7669),
            .I(N__7662));
    InMux I__1462 (
            .O(N__7666),
            .I(N__7657));
    InMux I__1461 (
            .O(N__7665),
            .I(N__7657));
    LocalMux I__1460 (
            .O(N__7662),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__1459 (
            .O(N__7657),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    IoInMux I__1458 (
            .O(N__7652),
            .I(N__7648));
    IoInMux I__1457 (
            .O(N__7651),
            .I(N__7644));
    LocalMux I__1456 (
            .O(N__7648),
            .I(N__7641));
    IoInMux I__1455 (
            .O(N__7647),
            .I(N__7638));
    LocalMux I__1454 (
            .O(N__7644),
            .I(N__7635));
    IoSpan4Mux I__1453 (
            .O(N__7641),
            .I(N__7632));
    LocalMux I__1452 (
            .O(N__7638),
            .I(N__7629));
    Span4Mux_s3_v I__1451 (
            .O(N__7635),
            .I(N__7626));
    Span4Mux_s3_h I__1450 (
            .O(N__7632),
            .I(N__7623));
    Span4Mux_s0_v I__1449 (
            .O(N__7629),
            .I(N__7620));
    Sp12to4 I__1448 (
            .O(N__7626),
            .I(N__7617));
    Sp12to4 I__1447 (
            .O(N__7623),
            .I(N__7614));
    Sp12to4 I__1446 (
            .O(N__7620),
            .I(N__7611));
    Span12Mux_s9_h I__1445 (
            .O(N__7617),
            .I(N__7608));
    Span12Mux_v I__1444 (
            .O(N__7614),
            .I(N__7605));
    Span12Mux_h I__1443 (
            .O(N__7611),
            .I(N__7602));
    Span12Mux_v I__1442 (
            .O(N__7608),
            .I(N__7598));
    Span12Mux_h I__1441 (
            .O(N__7605),
            .I(N__7593));
    Span12Mux_v I__1440 (
            .O(N__7602),
            .I(N__7593));
    InMux I__1439 (
            .O(N__7601),
            .I(N__7590));
    Odrv12 I__1438 (
            .O(N__7598),
            .I(TACK_OUTn));
    Odrv12 I__1437 (
            .O(N__7593),
            .I(TACK_OUTn));
    LocalMux I__1436 (
            .O(N__7590),
            .I(TACK_OUTn));
    InMux I__1435 (
            .O(N__7583),
            .I(N__7580));
    LocalMux I__1434 (
            .O(N__7580),
            .I(N__7577));
    Span12Mux_v I__1433 (
            .O(N__7577),
            .I(N__7574));
    Span12Mux_h I__1432 (
            .O(N__7574),
            .I(N__7571));
    Odrv12 I__1431 (
            .O(N__7571),
            .I(A_c_15));
    InMux I__1430 (
            .O(N__7568),
            .I(N__7565));
    LocalMux I__1429 (
            .O(N__7565),
            .I(N__7562));
    Span4Mux_h I__1428 (
            .O(N__7562),
            .I(N__7559));
    Span4Mux_h I__1427 (
            .O(N__7559),
            .I(N__7556));
    Odrv4 I__1426 (
            .O(N__7556),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ));
    SRMux I__1425 (
            .O(N__7553),
            .I(N__7550));
    LocalMux I__1424 (
            .O(N__7550),
            .I(N__7547));
    Span4Mux_h I__1423 (
            .O(N__7547),
            .I(N__7543));
    InMux I__1422 (
            .O(N__7546),
            .I(N__7540));
    Span4Mux_h I__1421 (
            .O(N__7543),
            .I(N__7537));
    LocalMux I__1420 (
            .O(N__7540),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    Odrv4 I__1419 (
            .O(N__7537),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    IoInMux I__1418 (
            .O(N__7532),
            .I(N__7529));
    LocalMux I__1417 (
            .O(N__7529),
            .I(N__7525));
    InMux I__1416 (
            .O(N__7528),
            .I(N__7522));
    Span12Mux_s4_v I__1415 (
            .O(N__7525),
            .I(N__7519));
    LocalMux I__1414 (
            .O(N__7522),
            .I(N__7516));
    Span12Mux_v I__1413 (
            .O(N__7519),
            .I(N__7511));
    Span12Mux_v I__1412 (
            .O(N__7516),
            .I(N__7511));
    Span12Mux_h I__1411 (
            .O(N__7511),
            .I(N__7508));
    Odrv12 I__1410 (
            .O(N__7508),
            .I(A_c_9));
    InMux I__1409 (
            .O(N__7505),
            .I(N__7502));
    LocalMux I__1408 (
            .O(N__7502),
            .I(N__7499));
    Odrv12 I__1407 (
            .O(N__7499),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ));
    CascadeMux I__1406 (
            .O(N__7496),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ));
    IoInMux I__1405 (
            .O(N__7493),
            .I(N__7490));
    LocalMux I__1404 (
            .O(N__7490),
            .I(N__7487));
    IoSpan4Mux I__1403 (
            .O(N__7487),
            .I(N__7484));
    IoSpan4Mux I__1402 (
            .O(N__7484),
            .I(N__7481));
    IoSpan4Mux I__1401 (
            .O(N__7481),
            .I(N__7478));
    Span4Mux_s2_v I__1400 (
            .O(N__7478),
            .I(N__7475));
    Sp12to4 I__1399 (
            .O(N__7475),
            .I(N__7471));
    InMux I__1398 (
            .O(N__7474),
            .I(N__7468));
    Span12Mux_s8_v I__1397 (
            .O(N__7471),
            .I(N__7465));
    LocalMux I__1396 (
            .O(N__7468),
            .I(N__7462));
    Span12Mux_v I__1395 (
            .O(N__7465),
            .I(N__7457));
    Span12Mux_h I__1394 (
            .O(N__7462),
            .I(N__7457));
    Odrv12 I__1393 (
            .O(N__7457),
            .I(A_c_10));
    InMux I__1392 (
            .O(N__7454),
            .I(N__7451));
    LocalMux I__1391 (
            .O(N__7451),
            .I(N__7448));
    Odrv12 I__1390 (
            .O(N__7448),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ));
    CascadeMux I__1389 (
            .O(N__7445),
            .I(\U712_CHIP_RAM.N_305_cascade_ ));
    InMux I__1388 (
            .O(N__7442),
            .I(N__7439));
    LocalMux I__1387 (
            .O(N__7439),
            .I(N__7436));
    Span4Mux_v I__1386 (
            .O(N__7436),
            .I(N__7433));
    Span4Mux_v I__1385 (
            .O(N__7433),
            .I(N__7430));
    Sp12to4 I__1384 (
            .O(N__7430),
            .I(N__7427));
    Span12Mux_h I__1383 (
            .O(N__7427),
            .I(N__7424));
    Odrv12 I__1382 (
            .O(N__7424),
            .I(A_c_14));
    InMux I__1381 (
            .O(N__7421),
            .I(N__7418));
    LocalMux I__1380 (
            .O(N__7418),
            .I(N__7415));
    Span12Mux_v I__1379 (
            .O(N__7415),
            .I(N__7412));
    Odrv12 I__1378 (
            .O(N__7412),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ));
    InMux I__1377 (
            .O(N__7409),
            .I(N__7401));
    InMux I__1376 (
            .O(N__7408),
            .I(N__7401));
    InMux I__1375 (
            .O(N__7407),
            .I(N__7398));
    InMux I__1374 (
            .O(N__7406),
            .I(N__7395));
    LocalMux I__1373 (
            .O(N__7401),
            .I(\U712_CHIP_RAM.N_469 ));
    LocalMux I__1372 (
            .O(N__7398),
            .I(\U712_CHIP_RAM.N_469 ));
    LocalMux I__1371 (
            .O(N__7395),
            .I(\U712_CHIP_RAM.N_469 ));
    CascadeMux I__1370 (
            .O(N__7388),
            .I(\U712_CHIP_RAM.N_438_cascade_ ));
    InMux I__1369 (
            .O(N__7385),
            .I(N__7382));
    LocalMux I__1368 (
            .O(N__7382),
            .I(N__7379));
    Odrv4 I__1367 (
            .O(N__7379),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ));
    CascadeMux I__1366 (
            .O(N__7376),
            .I(N__7370));
    CascadeMux I__1365 (
            .O(N__7375),
            .I(N__7364));
    InMux I__1364 (
            .O(N__7374),
            .I(N__7359));
    InMux I__1363 (
            .O(N__7373),
            .I(N__7356));
    InMux I__1362 (
            .O(N__7370),
            .I(N__7353));
    InMux I__1361 (
            .O(N__7369),
            .I(N__7350));
    InMux I__1360 (
            .O(N__7368),
            .I(N__7347));
    InMux I__1359 (
            .O(N__7367),
            .I(N__7344));
    InMux I__1358 (
            .O(N__7364),
            .I(N__7339));
    InMux I__1357 (
            .O(N__7363),
            .I(N__7339));
    CascadeMux I__1356 (
            .O(N__7362),
            .I(N__7335));
    LocalMux I__1355 (
            .O(N__7359),
            .I(N__7331));
    LocalMux I__1354 (
            .O(N__7356),
            .I(N__7328));
    LocalMux I__1353 (
            .O(N__7353),
            .I(N__7321));
    LocalMux I__1352 (
            .O(N__7350),
            .I(N__7321));
    LocalMux I__1351 (
            .O(N__7347),
            .I(N__7321));
    LocalMux I__1350 (
            .O(N__7344),
            .I(N__7311));
    LocalMux I__1349 (
            .O(N__7339),
            .I(N__7311));
    InMux I__1348 (
            .O(N__7338),
            .I(N__7308));
    InMux I__1347 (
            .O(N__7335),
            .I(N__7305));
    InMux I__1346 (
            .O(N__7334),
            .I(N__7302));
    Span4Mux_h I__1345 (
            .O(N__7331),
            .I(N__7297));
    Span4Mux_h I__1344 (
            .O(N__7328),
            .I(N__7297));
    Span4Mux_h I__1343 (
            .O(N__7321),
            .I(N__7291));
    InMux I__1342 (
            .O(N__7320),
            .I(N__7288));
    InMux I__1341 (
            .O(N__7319),
            .I(N__7281));
    InMux I__1340 (
            .O(N__7318),
            .I(N__7281));
    InMux I__1339 (
            .O(N__7317),
            .I(N__7281));
    InMux I__1338 (
            .O(N__7316),
            .I(N__7278));
    Span4Mux_h I__1337 (
            .O(N__7311),
            .I(N__7275));
    LocalMux I__1336 (
            .O(N__7308),
            .I(N__7268));
    LocalMux I__1335 (
            .O(N__7305),
            .I(N__7268));
    LocalMux I__1334 (
            .O(N__7302),
            .I(N__7268));
    Sp12to4 I__1333 (
            .O(N__7297),
            .I(N__7265));
    InMux I__1332 (
            .O(N__7296),
            .I(N__7258));
    InMux I__1331 (
            .O(N__7295),
            .I(N__7258));
    InMux I__1330 (
            .O(N__7294),
            .I(N__7258));
    Odrv4 I__1329 (
            .O(N__7291),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1328 (
            .O(N__7288),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1327 (
            .O(N__7281),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1326 (
            .O(N__7278),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1325 (
            .O(N__7275),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1324 (
            .O(N__7268),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv12 I__1323 (
            .O(N__7265),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1322 (
            .O(N__7258),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__1321 (
            .O(N__7241),
            .I(N__7237));
    CascadeMux I__1320 (
            .O(N__7240),
            .I(N__7233));
    InMux I__1319 (
            .O(N__7237),
            .I(N__7230));
    InMux I__1318 (
            .O(N__7236),
            .I(N__7227));
    InMux I__1317 (
            .O(N__7233),
            .I(N__7223));
    LocalMux I__1316 (
            .O(N__7230),
            .I(N__7218));
    LocalMux I__1315 (
            .O(N__7227),
            .I(N__7215));
    InMux I__1314 (
            .O(N__7226),
            .I(N__7208));
    LocalMux I__1313 (
            .O(N__7223),
            .I(N__7205));
    CascadeMux I__1312 (
            .O(N__7222),
            .I(N__7202));
    InMux I__1311 (
            .O(N__7221),
            .I(N__7198));
    Span4Mux_v I__1310 (
            .O(N__7218),
            .I(N__7195));
    Span4Mux_h I__1309 (
            .O(N__7215),
            .I(N__7192));
    InMux I__1308 (
            .O(N__7214),
            .I(N__7189));
    InMux I__1307 (
            .O(N__7213),
            .I(N__7186));
    InMux I__1306 (
            .O(N__7212),
            .I(N__7181));
    InMux I__1305 (
            .O(N__7211),
            .I(N__7181));
    LocalMux I__1304 (
            .O(N__7208),
            .I(N__7178));
    Span4Mux_v I__1303 (
            .O(N__7205),
            .I(N__7175));
    InMux I__1302 (
            .O(N__7202),
            .I(N__7172));
    InMux I__1301 (
            .O(N__7201),
            .I(N__7169));
    LocalMux I__1300 (
            .O(N__7198),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1299 (
            .O(N__7195),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1298 (
            .O(N__7192),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1297 (
            .O(N__7189),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1296 (
            .O(N__7186),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1295 (
            .O(N__7181),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1294 (
            .O(N__7178),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1293 (
            .O(N__7175),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1292 (
            .O(N__7172),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1291 (
            .O(N__7169),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__1290 (
            .O(N__7148),
            .I(N__7141));
    CascadeMux I__1289 (
            .O(N__7147),
            .I(N__7136));
    InMux I__1288 (
            .O(N__7146),
            .I(N__7133));
    CascadeMux I__1287 (
            .O(N__7145),
            .I(N__7128));
    InMux I__1286 (
            .O(N__7144),
            .I(N__7125));
    LocalMux I__1285 (
            .O(N__7141),
            .I(N__7122));
    InMux I__1284 (
            .O(N__7140),
            .I(N__7119));
    InMux I__1283 (
            .O(N__7139),
            .I(N__7116));
    InMux I__1282 (
            .O(N__7136),
            .I(N__7113));
    LocalMux I__1281 (
            .O(N__7133),
            .I(N__7106));
    InMux I__1280 (
            .O(N__7132),
            .I(N__7103));
    InMux I__1279 (
            .O(N__7131),
            .I(N__7098));
    InMux I__1278 (
            .O(N__7128),
            .I(N__7098));
    LocalMux I__1277 (
            .O(N__7125),
            .I(N__7087));
    Span4Mux_v I__1276 (
            .O(N__7122),
            .I(N__7087));
    LocalMux I__1275 (
            .O(N__7119),
            .I(N__7087));
    LocalMux I__1274 (
            .O(N__7116),
            .I(N__7087));
    LocalMux I__1273 (
            .O(N__7113),
            .I(N__7087));
    InMux I__1272 (
            .O(N__7112),
            .I(N__7080));
    InMux I__1271 (
            .O(N__7111),
            .I(N__7080));
    InMux I__1270 (
            .O(N__7110),
            .I(N__7080));
    InMux I__1269 (
            .O(N__7109),
            .I(N__7077));
    Odrv4 I__1268 (
            .O(N__7106),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1267 (
            .O(N__7103),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1266 (
            .O(N__7098),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1265 (
            .O(N__7087),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1264 (
            .O(N__7080),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1263 (
            .O(N__7077),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1262 (
            .O(N__7064),
            .I(N__7061));
    LocalMux I__1261 (
            .O(N__7061),
            .I(N__7058));
    Span4Mux_h I__1260 (
            .O(N__7058),
            .I(N__7055));
    Odrv4 I__1259 (
            .O(N__7055),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_a2_1 ));
    CascadeMux I__1258 (
            .O(N__7052),
            .I(N__7048));
    InMux I__1257 (
            .O(N__7051),
            .I(N__7043));
    InMux I__1256 (
            .O(N__7048),
            .I(N__7043));
    LocalMux I__1255 (
            .O(N__7043),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_a2_2 ));
    IoInMux I__1254 (
            .O(N__7040),
            .I(N__7037));
    LocalMux I__1253 (
            .O(N__7037),
            .I(N__7034));
    Span4Mux_s3_v I__1252 (
            .O(N__7034),
            .I(N__7031));
    Sp12to4 I__1251 (
            .O(N__7031),
            .I(N__7027));
    InMux I__1250 (
            .O(N__7030),
            .I(N__7024));
    Span12Mux_h I__1249 (
            .O(N__7027),
            .I(N__7019));
    LocalMux I__1248 (
            .O(N__7024),
            .I(N__7016));
    InMux I__1247 (
            .O(N__7023),
            .I(N__7013));
    InMux I__1246 (
            .O(N__7022),
            .I(N__7010));
    Odrv12 I__1245 (
            .O(N__7019),
            .I(DBENn_c));
    Odrv4 I__1244 (
            .O(N__7016),
            .I(DBENn_c));
    LocalMux I__1243 (
            .O(N__7013),
            .I(DBENn_c));
    LocalMux I__1242 (
            .O(N__7010),
            .I(DBENn_c));
    CascadeMux I__1241 (
            .O(N__7001),
            .I(N__6998));
    InMux I__1240 (
            .O(N__6998),
            .I(N__6991));
    InMux I__1239 (
            .O(N__6997),
            .I(N__6988));
    InMux I__1238 (
            .O(N__6996),
            .I(N__6985));
    InMux I__1237 (
            .O(N__6995),
            .I(N__6982));
    InMux I__1236 (
            .O(N__6994),
            .I(N__6979));
    LocalMux I__1235 (
            .O(N__6991),
            .I(N__6974));
    LocalMux I__1234 (
            .O(N__6988),
            .I(N__6971));
    LocalMux I__1233 (
            .O(N__6985),
            .I(N__6968));
    LocalMux I__1232 (
            .O(N__6982),
            .I(N__6965));
    LocalMux I__1231 (
            .O(N__6979),
            .I(N__6962));
    InMux I__1230 (
            .O(N__6978),
            .I(N__6959));
    InMux I__1229 (
            .O(N__6977),
            .I(N__6956));
    Span4Mux_v I__1228 (
            .O(N__6974),
            .I(N__6949));
    Span4Mux_h I__1227 (
            .O(N__6971),
            .I(N__6949));
    Span4Mux_v I__1226 (
            .O(N__6968),
            .I(N__6949));
    Span4Mux_v I__1225 (
            .O(N__6965),
            .I(N__6942));
    Span4Mux_v I__1224 (
            .O(N__6962),
            .I(N__6942));
    LocalMux I__1223 (
            .O(N__6959),
            .I(N__6942));
    LocalMux I__1222 (
            .O(N__6956),
            .I(DMA_CYCLEm));
    Odrv4 I__1221 (
            .O(N__6949),
            .I(DMA_CYCLEm));
    Odrv4 I__1220 (
            .O(N__6942),
            .I(DMA_CYCLEm));
    InMux I__1219 (
            .O(N__6935),
            .I(N__6932));
    LocalMux I__1218 (
            .O(N__6932),
            .I(\U712_CYCLE_TERM.N_321 ));
    IoInMux I__1217 (
            .O(N__6929),
            .I(N__6925));
    IoInMux I__1216 (
            .O(N__6928),
            .I(N__6922));
    LocalMux I__1215 (
            .O(N__6925),
            .I(N__6918));
    LocalMux I__1214 (
            .O(N__6922),
            .I(N__6915));
    IoInMux I__1213 (
            .O(N__6921),
            .I(N__6912));
    IoSpan4Mux I__1212 (
            .O(N__6918),
            .I(N__6909));
    IoSpan4Mux I__1211 (
            .O(N__6915),
            .I(N__6906));
    LocalMux I__1210 (
            .O(N__6912),
            .I(N__6903));
    Span4Mux_s1_h I__1209 (
            .O(N__6909),
            .I(N__6900));
    Sp12to4 I__1208 (
            .O(N__6906),
            .I(N__6897));
    Span4Mux_s3_v I__1207 (
            .O(N__6903),
            .I(N__6894));
    Sp12to4 I__1206 (
            .O(N__6900),
            .I(N__6891));
    Span12Mux_s3_v I__1205 (
            .O(N__6897),
            .I(N__6888));
    Sp12to4 I__1204 (
            .O(N__6894),
            .I(N__6885));
    Span12Mux_h I__1203 (
            .O(N__6891),
            .I(N__6881));
    Span12Mux_h I__1202 (
            .O(N__6888),
            .I(N__6876));
    Span12Mux_h I__1201 (
            .O(N__6885),
            .I(N__6876));
    InMux I__1200 (
            .O(N__6884),
            .I(N__6873));
    Odrv12 I__1199 (
            .O(N__6881),
            .I(TACK_EN));
    Odrv12 I__1198 (
            .O(N__6876),
            .I(TACK_EN));
    LocalMux I__1197 (
            .O(N__6873),
            .I(TACK_EN));
    InMux I__1196 (
            .O(N__6866),
            .I(N__6863));
    LocalMux I__1195 (
            .O(N__6863),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__1194 (
            .O(N__6860),
            .I(N__6857));
    LocalMux I__1193 (
            .O(N__6857),
            .I(N__6854));
    IoSpan4Mux I__1192 (
            .O(N__6854),
            .I(N__6851));
    Sp12to4 I__1191 (
            .O(N__6851),
            .I(N__6848));
    Odrv12 I__1190 (
            .O(N__6848),
            .I(CMA_c_2));
    InMux I__1189 (
            .O(N__6845),
            .I(N__6842));
    LocalMux I__1188 (
            .O(N__6842),
            .I(N__6839));
    Span12Mux_h I__1187 (
            .O(N__6839),
            .I(N__6836));
    Odrv12 I__1186 (
            .O(N__6836),
            .I(A_c_13));
    InMux I__1185 (
            .O(N__6833),
            .I(N__6830));
    LocalMux I__1184 (
            .O(N__6830),
            .I(N__6827));
    Odrv12 I__1183 (
            .O(N__6827),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ));
    CascadeMux I__1182 (
            .O(N__6824),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ));
    InMux I__1181 (
            .O(N__6821),
            .I(N__6813));
    InMux I__1180 (
            .O(N__6820),
            .I(N__6813));
    InMux I__1179 (
            .O(N__6819),
            .I(N__6810));
    InMux I__1178 (
            .O(N__6818),
            .I(N__6807));
    LocalMux I__1177 (
            .O(N__6813),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    LocalMux I__1176 (
            .O(N__6810),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    LocalMux I__1175 (
            .O(N__6807),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    CascadeMux I__1174 (
            .O(N__6800),
            .I(\U712_CHIP_RAM.N_442_cascade_ ));
    InMux I__1173 (
            .O(N__6797),
            .I(N__6791));
    InMux I__1172 (
            .O(N__6796),
            .I(N__6791));
    LocalMux I__1171 (
            .O(N__6791),
            .I(\U712_CHIP_RAM.N_441 ));
    InMux I__1170 (
            .O(N__6788),
            .I(N__6785));
    LocalMux I__1169 (
            .O(N__6785),
            .I(N__6782));
    Span4Mux_h I__1168 (
            .O(N__6782),
            .I(N__6779));
    Odrv4 I__1167 (
            .O(N__6779),
            .I(\U712_CHIP_RAM.CPU_TACK_8_iv_i_a2_1 ));
    CascadeMux I__1166 (
            .O(N__6776),
            .I(N__6772));
    CascadeMux I__1165 (
            .O(N__6775),
            .I(N__6769));
    InMux I__1164 (
            .O(N__6772),
            .I(N__6762));
    InMux I__1163 (
            .O(N__6769),
            .I(N__6762));
    InMux I__1162 (
            .O(N__6768),
            .I(N__6756));
    InMux I__1161 (
            .O(N__6767),
            .I(N__6753));
    LocalMux I__1160 (
            .O(N__6762),
            .I(N__6750));
    InMux I__1159 (
            .O(N__6761),
            .I(N__6745));
    InMux I__1158 (
            .O(N__6760),
            .I(N__6745));
    InMux I__1157 (
            .O(N__6759),
            .I(N__6742));
    LocalMux I__1156 (
            .O(N__6756),
            .I(\U712_CHIP_RAM.N_295 ));
    LocalMux I__1155 (
            .O(N__6753),
            .I(\U712_CHIP_RAM.N_295 ));
    Odrv4 I__1154 (
            .O(N__6750),
            .I(\U712_CHIP_RAM.N_295 ));
    LocalMux I__1153 (
            .O(N__6745),
            .I(\U712_CHIP_RAM.N_295 ));
    LocalMux I__1152 (
            .O(N__6742),
            .I(\U712_CHIP_RAM.N_295 ));
    InMux I__1151 (
            .O(N__6731),
            .I(N__6728));
    LocalMux I__1150 (
            .O(N__6728),
            .I(N__6724));
    InMux I__1149 (
            .O(N__6727),
            .I(N__6720));
    Span4Mux_v I__1148 (
            .O(N__6724),
            .I(N__6717));
    InMux I__1147 (
            .O(N__6723),
            .I(N__6714));
    LocalMux I__1146 (
            .O(N__6720),
            .I(N__6707));
    Sp12to4 I__1145 (
            .O(N__6717),
            .I(N__6707));
    LocalMux I__1144 (
            .O(N__6714),
            .I(N__6707));
    Span12Mux_h I__1143 (
            .O(N__6707),
            .I(N__6704));
    Span12Mux_v I__1142 (
            .O(N__6704),
            .I(N__6701));
    Odrv12 I__1141 (
            .O(N__6701),
            .I(AWEn_c));
    InMux I__1140 (
            .O(N__6698),
            .I(N__6693));
    InMux I__1139 (
            .O(N__6697),
            .I(N__6690));
    InMux I__1138 (
            .O(N__6696),
            .I(N__6687));
    LocalMux I__1137 (
            .O(N__6693),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    LocalMux I__1136 (
            .O(N__6690),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    LocalMux I__1135 (
            .O(N__6687),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    InMux I__1134 (
            .O(N__6680),
            .I(N__6677));
    LocalMux I__1133 (
            .O(N__6677),
            .I(N__6672));
    InMux I__1132 (
            .O(N__6676),
            .I(N__6669));
    InMux I__1131 (
            .O(N__6675),
            .I(N__6666));
    Odrv4 I__1130 (
            .O(N__6672),
            .I(\U712_CHIP_RAM.N_551 ));
    LocalMux I__1129 (
            .O(N__6669),
            .I(\U712_CHIP_RAM.N_551 ));
    LocalMux I__1128 (
            .O(N__6666),
            .I(\U712_CHIP_RAM.N_551 ));
    CascadeMux I__1127 (
            .O(N__6659),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_ ));
    CEMux I__1126 (
            .O(N__6656),
            .I(N__6653));
    LocalMux I__1125 (
            .O(N__6653),
            .I(N__6650));
    Span4Mux_v I__1124 (
            .O(N__6650),
            .I(N__6647));
    Odrv4 I__1123 (
            .O(N__6647),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ));
    InMux I__1122 (
            .O(N__6644),
            .I(N__6639));
    CascadeMux I__1121 (
            .O(N__6643),
            .I(N__6636));
    InMux I__1120 (
            .O(N__6642),
            .I(N__6630));
    LocalMux I__1119 (
            .O(N__6639),
            .I(N__6627));
    InMux I__1118 (
            .O(N__6636),
            .I(N__6624));
    InMux I__1117 (
            .O(N__6635),
            .I(N__6617));
    InMux I__1116 (
            .O(N__6634),
            .I(N__6617));
    InMux I__1115 (
            .O(N__6633),
            .I(N__6614));
    LocalMux I__1114 (
            .O(N__6630),
            .I(N__6607));
    Span4Mux_v I__1113 (
            .O(N__6627),
            .I(N__6607));
    LocalMux I__1112 (
            .O(N__6624),
            .I(N__6607));
    InMux I__1111 (
            .O(N__6623),
            .I(N__6602));
    InMux I__1110 (
            .O(N__6622),
            .I(N__6602));
    LocalMux I__1109 (
            .O(N__6617),
            .I(\U712_CHIP_RAM.N_458 ));
    LocalMux I__1108 (
            .O(N__6614),
            .I(\U712_CHIP_RAM.N_458 ));
    Odrv4 I__1107 (
            .O(N__6607),
            .I(\U712_CHIP_RAM.N_458 ));
    LocalMux I__1106 (
            .O(N__6602),
            .I(\U712_CHIP_RAM.N_458 ));
    InMux I__1105 (
            .O(N__6593),
            .I(N__6590));
    LocalMux I__1104 (
            .O(N__6590),
            .I(N__6587));
    Span4Mux_h I__1103 (
            .O(N__6587),
            .I(N__6584));
    Odrv4 I__1102 (
            .O(N__6584),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_0_0_0_a2_1 ));
    InMux I__1101 (
            .O(N__6581),
            .I(N__6578));
    LocalMux I__1100 (
            .O(N__6578),
            .I(N__6575));
    Odrv4 I__1099 (
            .O(N__6575),
            .I(\U712_CHIP_RAM.N_428 ));
    CascadeMux I__1098 (
            .O(N__6572),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_0_cascade_ ));
    CascadeMux I__1097 (
            .O(N__6569),
            .I(N__6566));
    InMux I__1096 (
            .O(N__6566),
            .I(N__6563));
    LocalMux I__1095 (
            .O(N__6563),
            .I(N__6559));
    InMux I__1094 (
            .O(N__6562),
            .I(N__6556));
    Span4Mux_v I__1093 (
            .O(N__6559),
            .I(N__6551));
    LocalMux I__1092 (
            .O(N__6556),
            .I(N__6551));
    Odrv4 I__1091 (
            .O(N__6551),
            .I(\U712_CHIP_RAM.N_300 ));
    CascadeMux I__1090 (
            .O(N__6548),
            .I(N__6543));
    CascadeMux I__1089 (
            .O(N__6547),
            .I(N__6528));
    InMux I__1088 (
            .O(N__6546),
            .I(N__6520));
    InMux I__1087 (
            .O(N__6543),
            .I(N__6512));
    CascadeMux I__1086 (
            .O(N__6542),
            .I(N__6509));
    InMux I__1085 (
            .O(N__6541),
            .I(N__6506));
    InMux I__1084 (
            .O(N__6540),
            .I(N__6503));
    InMux I__1083 (
            .O(N__6539),
            .I(N__6498));
    InMux I__1082 (
            .O(N__6538),
            .I(N__6498));
    InMux I__1081 (
            .O(N__6537),
            .I(N__6495));
    InMux I__1080 (
            .O(N__6536),
            .I(N__6488));
    InMux I__1079 (
            .O(N__6535),
            .I(N__6488));
    InMux I__1078 (
            .O(N__6534),
            .I(N__6488));
    InMux I__1077 (
            .O(N__6533),
            .I(N__6479));
    InMux I__1076 (
            .O(N__6532),
            .I(N__6479));
    InMux I__1075 (
            .O(N__6531),
            .I(N__6479));
    InMux I__1074 (
            .O(N__6528),
            .I(N__6479));
    InMux I__1073 (
            .O(N__6527),
            .I(N__6471));
    InMux I__1072 (
            .O(N__6526),
            .I(N__6471));
    InMux I__1071 (
            .O(N__6525),
            .I(N__6464));
    InMux I__1070 (
            .O(N__6524),
            .I(N__6464));
    InMux I__1069 (
            .O(N__6523),
            .I(N__6464));
    LocalMux I__1068 (
            .O(N__6520),
            .I(N__6461));
    InMux I__1067 (
            .O(N__6519),
            .I(N__6450));
    InMux I__1066 (
            .O(N__6518),
            .I(N__6450));
    InMux I__1065 (
            .O(N__6517),
            .I(N__6450));
    InMux I__1064 (
            .O(N__6516),
            .I(N__6450));
    InMux I__1063 (
            .O(N__6515),
            .I(N__6450));
    LocalMux I__1062 (
            .O(N__6512),
            .I(N__6447));
    InMux I__1061 (
            .O(N__6509),
            .I(N__6444));
    LocalMux I__1060 (
            .O(N__6506),
            .I(N__6439));
    LocalMux I__1059 (
            .O(N__6503),
            .I(N__6439));
    LocalMux I__1058 (
            .O(N__6498),
            .I(N__6430));
    LocalMux I__1057 (
            .O(N__6495),
            .I(N__6430));
    LocalMux I__1056 (
            .O(N__6488),
            .I(N__6430));
    LocalMux I__1055 (
            .O(N__6479),
            .I(N__6430));
    InMux I__1054 (
            .O(N__6478),
            .I(N__6424));
    InMux I__1053 (
            .O(N__6477),
            .I(N__6424));
    InMux I__1052 (
            .O(N__6476),
            .I(N__6421));
    LocalMux I__1051 (
            .O(N__6471),
            .I(N__6416));
    LocalMux I__1050 (
            .O(N__6464),
            .I(N__6416));
    Span4Mux_v I__1049 (
            .O(N__6461),
            .I(N__6411));
    LocalMux I__1048 (
            .O(N__6450),
            .I(N__6411));
    Span4Mux_v I__1047 (
            .O(N__6447),
            .I(N__6402));
    LocalMux I__1046 (
            .O(N__6444),
            .I(N__6402));
    Span4Mux_v I__1045 (
            .O(N__6439),
            .I(N__6402));
    Span4Mux_v I__1044 (
            .O(N__6430),
            .I(N__6402));
    InMux I__1043 (
            .O(N__6429),
            .I(N__6399));
    LocalMux I__1042 (
            .O(N__6424),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1041 (
            .O(N__6421),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv12 I__1040 (
            .O(N__6416),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1039 (
            .O(N__6411),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1038 (
            .O(N__6402),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1037 (
            .O(N__6399),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    CascadeMux I__1036 (
            .O(N__6386),
            .I(N__6383));
    InMux I__1035 (
            .O(N__6383),
            .I(N__6380));
    LocalMux I__1034 (
            .O(N__6380),
            .I(\U712_CHIP_RAM.N_438 ));
    IoInMux I__1033 (
            .O(N__6377),
            .I(N__6374));
    LocalMux I__1032 (
            .O(N__6374),
            .I(N__6371));
    Span4Mux_s3_v I__1031 (
            .O(N__6371),
            .I(N__6367));
    InMux I__1030 (
            .O(N__6370),
            .I(N__6364));
    Span4Mux_v I__1029 (
            .O(N__6367),
            .I(N__6361));
    LocalMux I__1028 (
            .O(N__6364),
            .I(N__6358));
    Span4Mux_h I__1027 (
            .O(N__6361),
            .I(N__6355));
    Span4Mux_v I__1026 (
            .O(N__6358),
            .I(N__6352));
    Odrv4 I__1025 (
            .O(N__6355),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1024 (
            .O(N__6352),
            .I(CONSTANT_ONE_NET));
    IoInMux I__1023 (
            .O(N__6347),
            .I(N__6344));
    LocalMux I__1022 (
            .O(N__6344),
            .I(N__6341));
    IoSpan4Mux I__1021 (
            .O(N__6341),
            .I(N__6338));
    Span4Mux_s2_v I__1020 (
            .O(N__6338),
            .I(N__6334));
    InMux I__1019 (
            .O(N__6337),
            .I(N__6331));
    Sp12to4 I__1018 (
            .O(N__6334),
            .I(N__6328));
    LocalMux I__1017 (
            .O(N__6331),
            .I(N__6325));
    Span12Mux_s8_v I__1016 (
            .O(N__6328),
            .I(N__6322));
    Span4Mux_v I__1015 (
            .O(N__6325),
            .I(N__6319));
    Span12Mux_v I__1014 (
            .O(N__6322),
            .I(N__6316));
    Sp12to4 I__1013 (
            .O(N__6319),
            .I(N__6313));
    Span12Mux_h I__1012 (
            .O(N__6316),
            .I(N__6310));
    Span12Mux_h I__1011 (
            .O(N__6313),
            .I(N__6307));
    Odrv12 I__1010 (
            .O(N__6310),
            .I(A_c_11));
    Odrv12 I__1009 (
            .O(N__6307),
            .I(A_c_11));
    InMux I__1008 (
            .O(N__6302),
            .I(N__6299));
    LocalMux I__1007 (
            .O(N__6299),
            .I(N__6296));
    Span4Mux_v I__1006 (
            .O(N__6296),
            .I(N__6293));
    Odrv4 I__1005 (
            .O(N__6293),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ));
    CascadeMux I__1004 (
            .O(N__6290),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ));
    IoInMux I__1003 (
            .O(N__6287),
            .I(N__6284));
    LocalMux I__1002 (
            .O(N__6284),
            .I(N__6281));
    Span4Mux_s3_v I__1001 (
            .O(N__6281),
            .I(N__6278));
    Span4Mux_h I__1000 (
            .O(N__6278),
            .I(N__6275));
    Span4Mux_h I__999 (
            .O(N__6275),
            .I(N__6272));
    Sp12to4 I__998 (
            .O(N__6272),
            .I(N__6269));
    Span12Mux_v I__997 (
            .O(N__6269),
            .I(N__6265));
    InMux I__996 (
            .O(N__6268),
            .I(N__6262));
    Odrv12 I__995 (
            .O(N__6265),
            .I(LATCH_CLK_c));
    LocalMux I__994 (
            .O(N__6262),
            .I(LATCH_CLK_c));
    InMux I__993 (
            .O(N__6257),
            .I(N__6254));
    LocalMux I__992 (
            .O(N__6254),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_a2_0_1 ));
    CascadeMux I__991 (
            .O(N__6251),
            .I(N__6246));
    InMux I__990 (
            .O(N__6250),
            .I(N__6243));
    InMux I__989 (
            .O(N__6249),
            .I(N__6240));
    InMux I__988 (
            .O(N__6246),
            .I(N__6237));
    LocalMux I__987 (
            .O(N__6243),
            .I(\U712_CHIP_RAM.N_533 ));
    LocalMux I__986 (
            .O(N__6240),
            .I(\U712_CHIP_RAM.N_533 ));
    LocalMux I__985 (
            .O(N__6237),
            .I(\U712_CHIP_RAM.N_533 ));
    CascadeMux I__984 (
            .O(N__6230),
            .I(\U712_CHIP_RAM.N_296_cascade_ ));
    CascadeMux I__983 (
            .O(N__6227),
            .I(N__6224));
    InMux I__982 (
            .O(N__6224),
            .I(N__6221));
    LocalMux I__981 (
            .O(N__6221),
            .I(N__6217));
    InMux I__980 (
            .O(N__6220),
            .I(N__6214));
    Odrv4 I__979 (
            .O(N__6217),
            .I(\U712_CHIP_RAM.N_550 ));
    LocalMux I__978 (
            .O(N__6214),
            .I(\U712_CHIP_RAM.N_550 ));
    CascadeMux I__977 (
            .O(N__6209),
            .I(N__6206));
    InMux I__976 (
            .O(N__6206),
            .I(N__6202));
    CascadeMux I__975 (
            .O(N__6205),
            .I(N__6199));
    LocalMux I__974 (
            .O(N__6202),
            .I(N__6196));
    InMux I__973 (
            .O(N__6199),
            .I(N__6187));
    Span4Mux_v I__972 (
            .O(N__6196),
            .I(N__6184));
    InMux I__971 (
            .O(N__6195),
            .I(N__6177));
    InMux I__970 (
            .O(N__6194),
            .I(N__6177));
    InMux I__969 (
            .O(N__6193),
            .I(N__6177));
    InMux I__968 (
            .O(N__6192),
            .I(N__6170));
    InMux I__967 (
            .O(N__6191),
            .I(N__6170));
    InMux I__966 (
            .O(N__6190),
            .I(N__6170));
    LocalMux I__965 (
            .O(N__6187),
            .I(\U712_CHIP_RAM.N_463 ));
    Odrv4 I__964 (
            .O(N__6184),
            .I(\U712_CHIP_RAM.N_463 ));
    LocalMux I__963 (
            .O(N__6177),
            .I(\U712_CHIP_RAM.N_463 ));
    LocalMux I__962 (
            .O(N__6170),
            .I(\U712_CHIP_RAM.N_463 ));
    InMux I__961 (
            .O(N__6161),
            .I(N__6158));
    LocalMux I__960 (
            .O(N__6158),
            .I(N__6154));
    InMux I__959 (
            .O(N__6157),
            .I(N__6151));
    Span4Mux_h I__958 (
            .O(N__6154),
            .I(N__6148));
    LocalMux I__957 (
            .O(N__6151),
            .I(N__6145));
    Odrv4 I__956 (
            .O(N__6148),
            .I(\U712_CHIP_RAM.N_546 ));
    Odrv4 I__955 (
            .O(N__6145),
            .I(\U712_CHIP_RAM.N_546 ));
    InMux I__954 (
            .O(N__6140),
            .I(N__6137));
    LocalMux I__953 (
            .O(N__6137),
            .I(N__6134));
    Span4Mux_h I__952 (
            .O(N__6134),
            .I(N__6122));
    InMux I__951 (
            .O(N__6133),
            .I(N__6119));
    InMux I__950 (
            .O(N__6132),
            .I(N__6116));
    InMux I__949 (
            .O(N__6131),
            .I(N__6111));
    InMux I__948 (
            .O(N__6130),
            .I(N__6111));
    InMux I__947 (
            .O(N__6129),
            .I(N__6106));
    InMux I__946 (
            .O(N__6128),
            .I(N__6106));
    InMux I__945 (
            .O(N__6127),
            .I(N__6099));
    InMux I__944 (
            .O(N__6126),
            .I(N__6099));
    InMux I__943 (
            .O(N__6125),
            .I(N__6099));
    Odrv4 I__942 (
            .O(N__6122),
            .I(\U712_CHIP_RAM.N_464 ));
    LocalMux I__941 (
            .O(N__6119),
            .I(\U712_CHIP_RAM.N_464 ));
    LocalMux I__940 (
            .O(N__6116),
            .I(\U712_CHIP_RAM.N_464 ));
    LocalMux I__939 (
            .O(N__6111),
            .I(\U712_CHIP_RAM.N_464 ));
    LocalMux I__938 (
            .O(N__6106),
            .I(\U712_CHIP_RAM.N_464 ));
    LocalMux I__937 (
            .O(N__6099),
            .I(\U712_CHIP_RAM.N_464 ));
    InMux I__936 (
            .O(N__6086),
            .I(N__6081));
    InMux I__935 (
            .O(N__6085),
            .I(N__6078));
    InMux I__934 (
            .O(N__6084),
            .I(N__6075));
    LocalMux I__933 (
            .O(N__6081),
            .I(\U712_CHIP_RAM.N_465 ));
    LocalMux I__932 (
            .O(N__6078),
            .I(\U712_CHIP_RAM.N_465 ));
    LocalMux I__931 (
            .O(N__6075),
            .I(\U712_CHIP_RAM.N_465 ));
    CascadeMux I__930 (
            .O(N__6068),
            .I(\U712_CHIP_RAM.N_465_cascade_ ));
    InMux I__929 (
            .O(N__6065),
            .I(N__6062));
    LocalMux I__928 (
            .O(N__6062),
            .I(N__6059));
    Span12Mux_v I__927 (
            .O(N__6059),
            .I(N__6056));
    Span12Mux_h I__926 (
            .O(N__6056),
            .I(N__6053));
    Odrv12 I__925 (
            .O(N__6053),
            .I(A_c_20));
    InMux I__924 (
            .O(N__6050),
            .I(N__6047));
    LocalMux I__923 (
            .O(N__6047),
            .I(N__6043));
    InMux I__922 (
            .O(N__6046),
            .I(N__6040));
    Odrv4 I__921 (
            .O(N__6043),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    LocalMux I__920 (
            .O(N__6040),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    InMux I__919 (
            .O(N__6035),
            .I(N__6031));
    InMux I__918 (
            .O(N__6034),
            .I(N__6028));
    LocalMux I__917 (
            .O(N__6031),
            .I(N__6025));
    LocalMux I__916 (
            .O(N__6028),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    Odrv12 I__915 (
            .O(N__6025),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    InMux I__914 (
            .O(N__6020),
            .I(N__6017));
    LocalMux I__913 (
            .O(N__6017),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0 ));
    CascadeMux I__912 (
            .O(N__6014),
            .I(N__6011));
    InMux I__911 (
            .O(N__6011),
            .I(N__6008));
    LocalMux I__910 (
            .O(N__6008),
            .I(N__6005));
    Odrv4 I__909 (
            .O(N__6005),
            .I(\U712_CHIP_RAM.DBENn_8_0_0 ));
    IoInMux I__908 (
            .O(N__6002),
            .I(N__5999));
    LocalMux I__907 (
            .O(N__5999),
            .I(N__5996));
    Span4Mux_s2_v I__906 (
            .O(N__5996),
            .I(N__5993));
    Span4Mux_v I__905 (
            .O(N__5993),
            .I(N__5990));
    Span4Mux_v I__904 (
            .O(N__5990),
            .I(N__5987));
    Span4Mux_v I__903 (
            .O(N__5987),
            .I(N__5983));
    InMux I__902 (
            .O(N__5986),
            .I(N__5980));
    Odrv4 I__901 (
            .O(N__5983),
            .I(DBDIR_c));
    LocalMux I__900 (
            .O(N__5980),
            .I(DBDIR_c));
    IoInMux I__899 (
            .O(N__5975),
            .I(N__5971));
    IoInMux I__898 (
            .O(N__5974),
            .I(N__5968));
    LocalMux I__897 (
            .O(N__5971),
            .I(N__5965));
    LocalMux I__896 (
            .O(N__5968),
            .I(N__5962));
    Span4Mux_s0_v I__895 (
            .O(N__5965),
            .I(N__5959));
    Span4Mux_s3_v I__894 (
            .O(N__5962),
            .I(N__5956));
    Span4Mux_v I__893 (
            .O(N__5959),
            .I(N__5953));
    Span4Mux_h I__892 (
            .O(N__5956),
            .I(N__5950));
    Sp12to4 I__891 (
            .O(N__5953),
            .I(N__5946));
    Span4Mux_h I__890 (
            .O(N__5950),
            .I(N__5943));
    IoInMux I__889 (
            .O(N__5949),
            .I(N__5940));
    Span12Mux_s11_h I__888 (
            .O(N__5946),
            .I(N__5935));
    Sp12to4 I__887 (
            .O(N__5943),
            .I(N__5935));
    LocalMux I__886 (
            .O(N__5940),
            .I(N__5932));
    Span12Mux_v I__885 (
            .O(N__5935),
            .I(N__5927));
    Span12Mux_s8_h I__884 (
            .O(N__5932),
            .I(N__5927));
    Odrv12 I__883 (
            .O(N__5927),
            .I(CLK40_PLL_i_i));
    IoInMux I__882 (
            .O(N__5924),
            .I(N__5921));
    LocalMux I__881 (
            .O(N__5921),
            .I(N__5918));
    IoSpan4Mux I__880 (
            .O(N__5918),
            .I(N__5915));
    Span4Mux_s3_v I__879 (
            .O(N__5915),
            .I(N__5912));
    Span4Mux_v I__878 (
            .O(N__5912),
            .I(N__5909));
    Odrv4 I__877 (
            .O(N__5909),
            .I(N_167_i));
    CascadeMux I__876 (
            .O(N__5906),
            .I(\U712_CHIP_RAM.N_533_cascade_ ));
    InMux I__875 (
            .O(N__5903),
            .I(N__5900));
    LocalMux I__874 (
            .O(N__5900),
            .I(\U712_CHIP_RAM.N_370 ));
    CascadeMux I__873 (
            .O(N__5897),
            .I(\U712_CHIP_RAM.N_391_cascade_ ));
    CascadeMux I__872 (
            .O(N__5894),
            .I(N__5891));
    InMux I__871 (
            .O(N__5891),
            .I(N__5888));
    LocalMux I__870 (
            .O(N__5888),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0 ));
    IoInMux I__869 (
            .O(N__5885),
            .I(N__5882));
    LocalMux I__868 (
            .O(N__5882),
            .I(N__5879));
    Span12Mux_s6_h I__867 (
            .O(N__5879),
            .I(N__5876));
    Span12Mux_h I__866 (
            .O(N__5876),
            .I(N__5873));
    Odrv12 I__865 (
            .O(N__5873),
            .I(CLK_EN_c));
    InMux I__864 (
            .O(N__5870),
            .I(N__5866));
    InMux I__863 (
            .O(N__5869),
            .I(N__5863));
    LocalMux I__862 (
            .O(N__5866),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__861 (
            .O(N__5863),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__860 (
            .O(N__5858),
            .I(N__5854));
    InMux I__859 (
            .O(N__5857),
            .I(N__5851));
    LocalMux I__858 (
            .O(N__5854),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__857 (
            .O(N__5851),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__856 (
            .O(N__5846),
            .I(N__5842));
    InMux I__855 (
            .O(N__5845),
            .I(N__5839));
    InMux I__854 (
            .O(N__5842),
            .I(N__5836));
    LocalMux I__853 (
            .O(N__5839),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__852 (
            .O(N__5836),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__851 (
            .O(N__5831),
            .I(N__5827));
    InMux I__850 (
            .O(N__5830),
            .I(N__5824));
    LocalMux I__849 (
            .O(N__5827),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__848 (
            .O(N__5824),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    CascadeMux I__847 (
            .O(N__5819),
            .I(\U712_CHIP_RAM.N_295_cascade_ ));
    CascadeMux I__846 (
            .O(N__5816),
            .I(N__5812));
    InMux I__845 (
            .O(N__5815),
            .I(N__5807));
    InMux I__844 (
            .O(N__5812),
            .I(N__5807));
    LocalMux I__843 (
            .O(N__5807),
            .I(N__5802));
    InMux I__842 (
            .O(N__5806),
            .I(N__5794));
    InMux I__841 (
            .O(N__5805),
            .I(N__5791));
    Span4Mux_h I__840 (
            .O(N__5802),
            .I(N__5788));
    InMux I__839 (
            .O(N__5801),
            .I(N__5785));
    InMux I__838 (
            .O(N__5800),
            .I(N__5782));
    InMux I__837 (
            .O(N__5799),
            .I(N__5777));
    InMux I__836 (
            .O(N__5798),
            .I(N__5777));
    InMux I__835 (
            .O(N__5797),
            .I(N__5774));
    LocalMux I__834 (
            .O(N__5794),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__833 (
            .O(N__5791),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__832 (
            .O(N__5788),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__831 (
            .O(N__5785),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__830 (
            .O(N__5782),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__829 (
            .O(N__5777),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__828 (
            .O(N__5774),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__827 (
            .O(N__5759),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_cascade_ ));
    InMux I__826 (
            .O(N__5756),
            .I(N__5753));
    LocalMux I__825 (
            .O(N__5753),
            .I(N__5749));
    InMux I__824 (
            .O(N__5752),
            .I(N__5746));
    Span4Mux_v I__823 (
            .O(N__5749),
            .I(N__5738));
    LocalMux I__822 (
            .O(N__5746),
            .I(N__5738));
    InMux I__821 (
            .O(N__5745),
            .I(N__5733));
    InMux I__820 (
            .O(N__5744),
            .I(N__5733));
    InMux I__819 (
            .O(N__5743),
            .I(N__5730));
    Odrv4 I__818 (
            .O(N__5738),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__817 (
            .O(N__5733),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__816 (
            .O(N__5730),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    CascadeMux I__815 (
            .O(N__5723),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_ ));
    CEMux I__814 (
            .O(N__5720),
            .I(N__5717));
    LocalMux I__813 (
            .O(N__5717),
            .I(N__5714));
    Span4Mux_h I__812 (
            .O(N__5714),
            .I(N__5711));
    Odrv4 I__811 (
            .O(N__5711),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_1 ));
    InMux I__810 (
            .O(N__5708),
            .I(N__5704));
    InMux I__809 (
            .O(N__5707),
            .I(N__5700));
    LocalMux I__808 (
            .O(N__5704),
            .I(N__5693));
    InMux I__807 (
            .O(N__5703),
            .I(N__5690));
    LocalMux I__806 (
            .O(N__5700),
            .I(N__5687));
    InMux I__805 (
            .O(N__5699),
            .I(N__5684));
    InMux I__804 (
            .O(N__5698),
            .I(N__5679));
    InMux I__803 (
            .O(N__5697),
            .I(N__5679));
    CascadeMux I__802 (
            .O(N__5696),
            .I(N__5674));
    Span4Mux_h I__801 (
            .O(N__5693),
            .I(N__5671));
    LocalMux I__800 (
            .O(N__5690),
            .I(N__5666));
    Span4Mux_h I__799 (
            .O(N__5687),
            .I(N__5666));
    LocalMux I__798 (
            .O(N__5684),
            .I(N__5661));
    LocalMux I__797 (
            .O(N__5679),
            .I(N__5661));
    InMux I__796 (
            .O(N__5678),
            .I(N__5658));
    InMux I__795 (
            .O(N__5677),
            .I(N__5653));
    InMux I__794 (
            .O(N__5674),
            .I(N__5653));
    Odrv4 I__793 (
            .O(N__5671),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__792 (
            .O(N__5666),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__791 (
            .O(N__5661),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__790 (
            .O(N__5658),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__789 (
            .O(N__5653),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CascadeMux I__788 (
            .O(N__5642),
            .I(\U712_CHIP_RAM.N_463_cascade_ ));
    CascadeMux I__787 (
            .O(N__5639),
            .I(N__5636));
    InMux I__786 (
            .O(N__5636),
            .I(N__5632));
    InMux I__785 (
            .O(N__5635),
            .I(N__5629));
    LocalMux I__784 (
            .O(N__5632),
            .I(N__5625));
    LocalMux I__783 (
            .O(N__5629),
            .I(N__5622));
    CascadeMux I__782 (
            .O(N__5628),
            .I(N__5619));
    Span4Mux_h I__781 (
            .O(N__5625),
            .I(N__5615));
    Span4Mux_h I__780 (
            .O(N__5622),
            .I(N__5612));
    InMux I__779 (
            .O(N__5619),
            .I(N__5607));
    InMux I__778 (
            .O(N__5618),
            .I(N__5607));
    Odrv4 I__777 (
            .O(N__5615),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__776 (
            .O(N__5612),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__775 (
            .O(N__5607),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    CascadeMux I__774 (
            .O(N__5600),
            .I(\U712_CHIP_RAM.N_385_cascade_ ));
    InMux I__773 (
            .O(N__5597),
            .I(N__5594));
    LocalMux I__772 (
            .O(N__5594),
            .I(\U712_CHIP_RAM.N_384 ));
    CascadeMux I__771 (
            .O(N__5591),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0_cascade_ ));
    InMux I__770 (
            .O(N__5588),
            .I(N__5585));
    LocalMux I__769 (
            .O(N__5585),
            .I(\U712_CHIP_RAM.N_461 ));
    CascadeMux I__768 (
            .O(N__5582),
            .I(N__5579));
    InMux I__767 (
            .O(N__5579),
            .I(N__5576));
    LocalMux I__766 (
            .O(N__5576),
            .I(N__5573));
    Span4Mux_v I__765 (
            .O(N__5573),
            .I(N__5568));
    InMux I__764 (
            .O(N__5572),
            .I(N__5563));
    InMux I__763 (
            .O(N__5571),
            .I(N__5563));
    Odrv4 I__762 (
            .O(N__5568),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    LocalMux I__761 (
            .O(N__5563),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    CascadeMux I__760 (
            .O(N__5558),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0_a2_0_cascade_ ));
    CEMux I__759 (
            .O(N__5555),
            .I(N__5550));
    CEMux I__758 (
            .O(N__5554),
            .I(N__5547));
    CEMux I__757 (
            .O(N__5553),
            .I(N__5544));
    LocalMux I__756 (
            .O(N__5550),
            .I(N__5541));
    LocalMux I__755 (
            .O(N__5547),
            .I(N__5538));
    LocalMux I__754 (
            .O(N__5544),
            .I(N__5535));
    Span4Mux_h I__753 (
            .O(N__5541),
            .I(N__5530));
    Span4Mux_h I__752 (
            .O(N__5538),
            .I(N__5530));
    Span4Mux_v I__751 (
            .O(N__5535),
            .I(N__5527));
    Odrv4 I__750 (
            .O(N__5530),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__749 (
            .O(N__5527),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__748 (
            .O(N__5522),
            .I(N__5519));
    LocalMux I__747 (
            .O(N__5519),
            .I(N__5516));
    Span4Mux_h I__746 (
            .O(N__5516),
            .I(N__5513));
    Odrv4 I__745 (
            .O(N__5513),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0_a2_0 ));
    CascadeMux I__744 (
            .O(N__5510),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_1_cascade_ ));
    InMux I__743 (
            .O(N__5507),
            .I(N__5504));
    LocalMux I__742 (
            .O(N__5504),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    CascadeMux I__741 (
            .O(N__5501),
            .I(N__5495));
    CascadeMux I__740 (
            .O(N__5500),
            .I(N__5492));
    InMux I__739 (
            .O(N__5499),
            .I(N__5482));
    InMux I__738 (
            .O(N__5498),
            .I(N__5482));
    InMux I__737 (
            .O(N__5495),
            .I(N__5482));
    InMux I__736 (
            .O(N__5492),
            .I(N__5482));
    InMux I__735 (
            .O(N__5491),
            .I(N__5477));
    LocalMux I__734 (
            .O(N__5482),
            .I(N__5474));
    InMux I__733 (
            .O(N__5481),
            .I(N__5471));
    InMux I__732 (
            .O(N__5480),
            .I(N__5468));
    LocalMux I__731 (
            .O(N__5477),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    Odrv4 I__730 (
            .O(N__5474),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__729 (
            .O(N__5471),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__728 (
            .O(N__5468),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__727 (
            .O(N__5459),
            .I(N__5456));
    LocalMux I__726 (
            .O(N__5456),
            .I(\U712_CHIP_RAM.N_419 ));
    InMux I__725 (
            .O(N__5453),
            .I(N__5450));
    LocalMux I__724 (
            .O(N__5450),
            .I(N__5447));
    Odrv12 I__723 (
            .O(N__5447),
            .I(\U712_BYTE_ENABLE.N_326 ));
    InMux I__722 (
            .O(N__5444),
            .I(N__5441));
    LocalMux I__721 (
            .O(N__5441),
            .I(N__5438));
    Odrv4 I__720 (
            .O(N__5438),
            .I(\U712_BYTE_ENABLE.N_323 ));
    InMux I__719 (
            .O(N__5435),
            .I(N__5432));
    LocalMux I__718 (
            .O(N__5432),
            .I(N__5429));
    Odrv12 I__717 (
            .O(N__5429),
            .I(\U712_BYTE_ENABLE.N_324 ));
    InMux I__716 (
            .O(N__5426),
            .I(N__5423));
    LocalMux I__715 (
            .O(N__5423),
            .I(N__5420));
    Span4Mux_h I__714 (
            .O(N__5420),
            .I(N__5417));
    Sp12to4 I__713 (
            .O(N__5417),
            .I(N__5414));
    Span12Mux_v I__712 (
            .O(N__5414),
            .I(N__5411));
    Odrv12 I__711 (
            .O(N__5411),
            .I(A_c_17));
    InMux I__710 (
            .O(N__5408),
            .I(N__5399));
    InMux I__709 (
            .O(N__5407),
            .I(N__5392));
    InMux I__708 (
            .O(N__5406),
            .I(N__5392));
    InMux I__707 (
            .O(N__5405),
            .I(N__5392));
    InMux I__706 (
            .O(N__5404),
            .I(N__5385));
    InMux I__705 (
            .O(N__5403),
            .I(N__5385));
    InMux I__704 (
            .O(N__5402),
            .I(N__5385));
    LocalMux I__703 (
            .O(N__5399),
            .I(N__5382));
    LocalMux I__702 (
            .O(N__5392),
            .I(\U712_CHIP_RAM.N_90_i ));
    LocalMux I__701 (
            .O(N__5385),
            .I(\U712_CHIP_RAM.N_90_i ));
    Odrv4 I__700 (
            .O(N__5382),
            .I(\U712_CHIP_RAM.N_90_i ));
    InMux I__699 (
            .O(N__5375),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    IoInMux I__698 (
            .O(N__5372),
            .I(N__5369));
    LocalMux I__697 (
            .O(N__5369),
            .I(N__5366));
    IoSpan4Mux I__696 (
            .O(N__5366),
            .I(N__5363));
    Span4Mux_s2_v I__695 (
            .O(N__5363),
            .I(N__5360));
    Sp12to4 I__694 (
            .O(N__5360),
            .I(N__5357));
    Odrv12 I__693 (
            .O(N__5357),
            .I(N_188_i));
    InMux I__692 (
            .O(N__5354),
            .I(N__5350));
    InMux I__691 (
            .O(N__5353),
            .I(N__5347));
    LocalMux I__690 (
            .O(N__5350),
            .I(N__5342));
    LocalMux I__689 (
            .O(N__5347),
            .I(N__5342));
    Odrv4 I__688 (
            .O(N__5342),
            .I(\U712_CHIP_RAM.N_302 ));
    CascadeMux I__687 (
            .O(N__5339),
            .I(N__5336));
    InMux I__686 (
            .O(N__5336),
            .I(N__5332));
    InMux I__685 (
            .O(N__5335),
            .I(N__5329));
    LocalMux I__684 (
            .O(N__5332),
            .I(N__5324));
    LocalMux I__683 (
            .O(N__5329),
            .I(N__5324));
    Span4Mux_v I__682 (
            .O(N__5324),
            .I(N__5321));
    Odrv4 I__681 (
            .O(N__5321),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ));
    InMux I__680 (
            .O(N__5318),
            .I(N__5315));
    LocalMux I__679 (
            .O(N__5315),
            .I(\U712_CHIP_RAM.N_455 ));
    CascadeMux I__678 (
            .O(N__5312),
            .I(\U712_CHIP_RAM.N_417_cascade_ ));
    InMux I__677 (
            .O(N__5309),
            .I(N__5306));
    LocalMux I__676 (
            .O(N__5306),
            .I(N__5303));
    Span12Mux_h I__675 (
            .O(N__5303),
            .I(N__5300));
    Span12Mux_v I__674 (
            .O(N__5300),
            .I(N__5297));
    Odrv12 I__673 (
            .O(N__5297),
            .I(RAMSPACEn_c));
    InMux I__672 (
            .O(N__5294),
            .I(N__5291));
    LocalMux I__671 (
            .O(N__5291),
            .I(N__5285));
    InMux I__670 (
            .O(N__5290),
            .I(N__5278));
    InMux I__669 (
            .O(N__5289),
            .I(N__5278));
    InMux I__668 (
            .O(N__5288),
            .I(N__5278));
    Odrv4 I__667 (
            .O(N__5285),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__666 (
            .O(N__5278),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__665 (
            .O(N__5273),
            .I(N__5270));
    LocalMux I__664 (
            .O(N__5270),
            .I(N__5266));
    InMux I__663 (
            .O(N__5269),
            .I(N__5263));
    Span4Mux_h I__662 (
            .O(N__5266),
            .I(N__5260));
    LocalMux I__661 (
            .O(N__5263),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv4 I__660 (
            .O(N__5260),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__659 (
            .O(N__5255),
            .I(N__5252));
    LocalMux I__658 (
            .O(N__5252),
            .I(N__5249));
    Span4Mux_h I__657 (
            .O(N__5249),
            .I(N__5246));
    Odrv4 I__656 (
            .O(N__5246),
            .I(\U712_CHIP_RAM.REFRESH5lto7_0 ));
    InMux I__655 (
            .O(N__5243),
            .I(N__5240));
    LocalMux I__654 (
            .O(N__5240),
            .I(N__5237));
    Span4Mux_h I__653 (
            .O(N__5237),
            .I(N__5234));
    Odrv4 I__652 (
            .O(N__5234),
            .I(\U712_CHIP_RAM.REFRESH5lt7 ));
    InMux I__651 (
            .O(N__5231),
            .I(N__5228));
    LocalMux I__650 (
            .O(N__5228),
            .I(N__5224));
    InMux I__649 (
            .O(N__5227),
            .I(N__5221));
    Odrv4 I__648 (
            .O(N__5224),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0 ));
    LocalMux I__647 (
            .O(N__5221),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0 ));
    InMux I__646 (
            .O(N__5216),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__645 (
            .O(N__5213),
            .I(N__5210));
    LocalMux I__644 (
            .O(N__5210),
            .I(N__5207));
    Odrv4 I__643 (
            .O(N__5207),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__642 (
            .O(N__5204),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__641 (
            .O(N__5201),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__640 (
            .O(N__5198),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__639 (
            .O(N__5195),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__638 (
            .O(N__5192),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__637 (
            .O(N__5189),
            .I(N__5183));
    InMux I__636 (
            .O(N__5188),
            .I(N__5183));
    LocalMux I__635 (
            .O(N__5183),
            .I(N__5180));
    Odrv4 I__634 (
            .O(N__5180),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ));
    IoInMux I__633 (
            .O(N__5177),
            .I(N__5174));
    LocalMux I__632 (
            .O(N__5174),
            .I(N__5171));
    IoSpan4Mux I__631 (
            .O(N__5171),
            .I(N__5168));
    Sp12to4 I__630 (
            .O(N__5168),
            .I(N__5165));
    Span12Mux_s7_h I__629 (
            .O(N__5165),
            .I(N__5162));
    Odrv12 I__628 (
            .O(N__5162),
            .I(N_176_i));
    InMux I__627 (
            .O(N__5159),
            .I(N__5156));
    LocalMux I__626 (
            .O(N__5156),
            .I(N__5153));
    Odrv12 I__625 (
            .O(N__5153),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ));
    InMux I__624 (
            .O(N__5150),
            .I(N__5147));
    LocalMux I__623 (
            .O(N__5147),
            .I(N__5144));
    Span4Mux_v I__622 (
            .O(N__5144),
            .I(N__5141));
    Span4Mux_h I__621 (
            .O(N__5141),
            .I(N__5138));
    Sp12to4 I__620 (
            .O(N__5138),
            .I(N__5135));
    Odrv12 I__619 (
            .O(N__5135),
            .I(A_c_12));
    InMux I__618 (
            .O(N__5132),
            .I(N__5129));
    LocalMux I__617 (
            .O(N__5129),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER19 ));
    CascadeMux I__616 (
            .O(N__5126),
            .I(\U712_CHIP_RAM.N_464_cascade_ ));
    CascadeMux I__615 (
            .O(N__5123),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ));
    InMux I__614 (
            .O(N__5120),
            .I(N__5117));
    LocalMux I__613 (
            .O(N__5117),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0 ));
    InMux I__612 (
            .O(N__5114),
            .I(N__5111));
    LocalMux I__611 (
            .O(N__5111),
            .I(\U712_CHIP_RAM.N_390 ));
    InMux I__610 (
            .O(N__5108),
            .I(N__5105));
    LocalMux I__609 (
            .O(N__5105),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ));
    InMux I__608 (
            .O(N__5102),
            .I(N__5098));
    InMux I__607 (
            .O(N__5101),
            .I(N__5095));
    LocalMux I__606 (
            .O(N__5098),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ));
    LocalMux I__605 (
            .O(N__5095),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ));
    CascadeMux I__604 (
            .O(N__5090),
            .I(N__5087));
    InMux I__603 (
            .O(N__5087),
            .I(N__5084));
    LocalMux I__602 (
            .O(N__5084),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3 ));
    InMux I__601 (
            .O(N__5081),
            .I(N__5077));
    InMux I__600 (
            .O(N__5080),
            .I(N__5074));
    LocalMux I__599 (
            .O(N__5077),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ));
    LocalMux I__598 (
            .O(N__5074),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ));
    InMux I__597 (
            .O(N__5069),
            .I(N__5065));
    CascadeMux I__596 (
            .O(N__5068),
            .I(N__5062));
    LocalMux I__595 (
            .O(N__5065),
            .I(N__5059));
    InMux I__594 (
            .O(N__5062),
            .I(N__5056));
    Odrv4 I__593 (
            .O(N__5059),
            .I(DBR_SYNC_i_1));
    LocalMux I__592 (
            .O(N__5056),
            .I(DBR_SYNC_i_1));
    InMux I__591 (
            .O(N__5051),
            .I(N__5048));
    LocalMux I__590 (
            .O(N__5048),
            .I(DBR_SYNCZ0Z_0));
    InMux I__589 (
            .O(N__5045),
            .I(N__5042));
    LocalMux I__588 (
            .O(N__5042),
            .I(N__5039));
    Span4Mux_h I__587 (
            .O(N__5039),
            .I(N__5036));
    Sp12to4 I__586 (
            .O(N__5036),
            .I(N__5033));
    Span12Mux_v I__585 (
            .O(N__5033),
            .I(N__5030));
    Odrv12 I__584 (
            .O(N__5030),
            .I(A_c_5));
    CEMux I__583 (
            .O(N__5027),
            .I(N__5023));
    CEMux I__582 (
            .O(N__5026),
            .I(N__5018));
    LocalMux I__581 (
            .O(N__5023),
            .I(N__5015));
    CEMux I__580 (
            .O(N__5022),
            .I(N__5012));
    CEMux I__579 (
            .O(N__5021),
            .I(N__5009));
    LocalMux I__578 (
            .O(N__5018),
            .I(N__5006));
    Span4Mux_v I__577 (
            .O(N__5015),
            .I(N__5001));
    LocalMux I__576 (
            .O(N__5012),
            .I(N__5001));
    LocalMux I__575 (
            .O(N__5009),
            .I(N__4998));
    Span4Mux_h I__574 (
            .O(N__5006),
            .I(N__4995));
    Span4Mux_h I__573 (
            .O(N__5001),
            .I(N__4992));
    Span4Mux_v I__572 (
            .O(N__4998),
            .I(N__4989));
    Odrv4 I__571 (
            .O(N__4995),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    Odrv4 I__570 (
            .O(N__4992),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    Odrv4 I__569 (
            .O(N__4989),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    InMux I__568 (
            .O(N__4982),
            .I(N__4979));
    LocalMux I__567 (
            .O(N__4979),
            .I(N__4976));
    Sp12to4 I__566 (
            .O(N__4976),
            .I(N__4973));
    Span12Mux_v I__565 (
            .O(N__4973),
            .I(N__4970));
    Span12Mux_h I__564 (
            .O(N__4970),
            .I(N__4967));
    Odrv12 I__563 (
            .O(N__4967),
            .I(A_c_16));
    InMux I__562 (
            .O(N__4964),
            .I(N__4961));
    LocalMux I__561 (
            .O(N__4961),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ));
    InMux I__560 (
            .O(N__4958),
            .I(N__4955));
    LocalMux I__559 (
            .O(N__4955),
            .I(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a3_0_a2_0 ));
    IoInMux I__558 (
            .O(N__4952),
            .I(N__4949));
    LocalMux I__557 (
            .O(N__4949),
            .I(N__4946));
    IoSpan4Mux I__556 (
            .O(N__4946),
            .I(N__4943));
    Sp12to4 I__555 (
            .O(N__4943),
            .I(N__4940));
    Span12Mux_s7_h I__554 (
            .O(N__4940),
            .I(N__4937));
    Span12Mux_h I__553 (
            .O(N__4937),
            .I(N__4934));
    Odrv12 I__552 (
            .O(N__4934),
            .I(N_178_i));
    InMux I__551 (
            .O(N__4931),
            .I(N__4925));
    InMux I__550 (
            .O(N__4930),
            .I(N__4925));
    LocalMux I__549 (
            .O(N__4925),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ));
    CascadeMux I__548 (
            .O(N__4922),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_ ));
    InMux I__547 (
            .O(N__4919),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ));
    InMux I__546 (
            .O(N__4916),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ));
    InMux I__545 (
            .O(N__4913),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ));
    InMux I__544 (
            .O(N__4910),
            .I(N__4907));
    LocalMux I__543 (
            .O(N__4907),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ));
    CascadeMux I__542 (
            .O(N__4904),
            .I(N__4900));
    InMux I__541 (
            .O(N__4903),
            .I(N__4897));
    InMux I__540 (
            .O(N__4900),
            .I(N__4894));
    LocalMux I__539 (
            .O(N__4897),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ));
    LocalMux I__538 (
            .O(N__4894),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ));
    CascadeMux I__537 (
            .O(N__4889),
            .I(N__4886));
    InMux I__536 (
            .O(N__4886),
            .I(N__4883));
    LocalMux I__535 (
            .O(N__4883),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ));
    InMux I__534 (
            .O(N__4880),
            .I(N__4876));
    InMux I__533 (
            .O(N__4879),
            .I(N__4873));
    LocalMux I__532 (
            .O(N__4876),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_1 ));
    LocalMux I__531 (
            .O(N__4873),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_1 ));
    CascadeMux I__530 (
            .O(N__4868),
            .I(\U712_CHIP_RAM.N_298_cascade_ ));
    CascadeMux I__529 (
            .O(N__4865),
            .I(\U712_CHIP_RAM.N_300_cascade_ ));
    InMux I__528 (
            .O(N__4862),
            .I(N__4859));
    LocalMux I__527 (
            .O(N__4859),
            .I(N__4856));
    Odrv4 I__526 (
            .O(N__4856),
            .I(\U712_CHIP_RAM.N_310 ));
    CascadeMux I__525 (
            .O(N__4853),
            .I(\U712_CHIP_RAM.N_310_cascade_ ));
    InMux I__524 (
            .O(N__4850),
            .I(N__4846));
    InMux I__523 (
            .O(N__4849),
            .I(N__4843));
    LocalMux I__522 (
            .O(N__4846),
            .I(\U712_CHIP_RAM.N_313 ));
    LocalMux I__521 (
            .O(N__4843),
            .I(\U712_CHIP_RAM.N_313 ));
    InMux I__520 (
            .O(N__4838),
            .I(N__4835));
    LocalMux I__519 (
            .O(N__4835),
            .I(\U712_CHIP_RAM.N_389 ));
    InMux I__518 (
            .O(N__4832),
            .I(N__4829));
    LocalMux I__517 (
            .O(N__4829),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_5 ));
    InMux I__516 (
            .O(N__4826),
            .I(N__4823));
    LocalMux I__515 (
            .O(N__4823),
            .I(N__4820));
    Span4Mux_h I__514 (
            .O(N__4820),
            .I(N__4817));
    Sp12to4 I__513 (
            .O(N__4817),
            .I(N__4814));
    Span12Mux_v I__512 (
            .O(N__4814),
            .I(N__4811));
    Odrv12 I__511 (
            .O(N__4811),
            .I(A_c_18));
    CEMux I__510 (
            .O(N__4808),
            .I(N__4805));
    LocalMux I__509 (
            .O(N__4805),
            .I(N__4802));
    Odrv4 I__508 (
            .O(N__4802),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0 ));
    InMux I__507 (
            .O(N__4799),
            .I(N__4796));
    LocalMux I__506 (
            .O(N__4796),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    CascadeMux I__505 (
            .O(N__4793),
            .I(N__4790));
    InMux I__504 (
            .O(N__4790),
            .I(N__4787));
    LocalMux I__503 (
            .O(N__4787),
            .I(N__4784));
    Odrv4 I__502 (
            .O(N__4784),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_a2_1_0 ));
    CascadeMux I__501 (
            .O(N__4781),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_165_i_i_0_cascade_ ));
    InMux I__500 (
            .O(N__4778),
            .I(N__4775));
    LocalMux I__499 (
            .O(N__4775),
            .I(N__4772));
    Odrv4 I__498 (
            .O(N__4772),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    CascadeMux I__497 (
            .O(N__4769),
            .I(\U712_CHIP_RAM.N_90_i_cascade_ ));
    InMux I__496 (
            .O(N__4766),
            .I(N__4763));
    LocalMux I__495 (
            .O(N__4763),
            .I(N__4760));
    Span4Mux_v I__494 (
            .O(N__4760),
            .I(N__4757));
    Span4Mux_v I__493 (
            .O(N__4757),
            .I(N__4754));
    Sp12to4 I__492 (
            .O(N__4754),
            .I(N__4751));
    Odrv12 I__491 (
            .O(N__4751),
            .I(A_c_7));
    InMux I__490 (
            .O(N__4748),
            .I(N__4745));
    LocalMux I__489 (
            .O(N__4745),
            .I(N__4742));
    Span4Mux_v I__488 (
            .O(N__4742),
            .I(N__4739));
    Span4Mux_v I__487 (
            .O(N__4739),
            .I(N__4736));
    Sp12to4 I__486 (
            .O(N__4736),
            .I(N__4733));
    Odrv12 I__485 (
            .O(N__4733),
            .I(A_c_8));
    CEMux I__484 (
            .O(N__4730),
            .I(N__4727));
    LocalMux I__483 (
            .O(N__4727),
            .I(N__4724));
    Span4Mux_v I__482 (
            .O(N__4724),
            .I(N__4721));
    Odrv4 I__481 (
            .O(N__4721),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0 ));
    InMux I__480 (
            .O(N__4718),
            .I(N__4715));
    LocalMux I__479 (
            .O(N__4715),
            .I(N__4711));
    InMux I__478 (
            .O(N__4714),
            .I(N__4708));
    Span4Mux_v I__477 (
            .O(N__4711),
            .I(N__4703));
    LocalMux I__476 (
            .O(N__4708),
            .I(N__4703));
    Span4Mux_v I__475 (
            .O(N__4703),
            .I(N__4700));
    Sp12to4 I__474 (
            .O(N__4700),
            .I(N__4697));
    Span12Mux_h I__473 (
            .O(N__4697),
            .I(N__4694));
    Odrv12 I__472 (
            .O(N__4694),
            .I(DBRn_c));
    IoInMux I__471 (
            .O(N__4691),
            .I(N__4688));
    LocalMux I__470 (
            .O(N__4688),
            .I(N__4685));
    Span12Mux_s9_v I__469 (
            .O(N__4685),
            .I(N__4682));
    Odrv12 I__468 (
            .O(N__4682),
            .I(VBENn_c));
    InMux I__467 (
            .O(N__4679),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__466 (
            .O(N__4676),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__465 (
            .O(N__4673),
            .I(N__4649));
    ClkMux I__464 (
            .O(N__4672),
            .I(N__4649));
    ClkMux I__463 (
            .O(N__4671),
            .I(N__4649));
    ClkMux I__462 (
            .O(N__4670),
            .I(N__4649));
    ClkMux I__461 (
            .O(N__4669),
            .I(N__4649));
    ClkMux I__460 (
            .O(N__4668),
            .I(N__4649));
    ClkMux I__459 (
            .O(N__4667),
            .I(N__4649));
    ClkMux I__458 (
            .O(N__4666),
            .I(N__4649));
    GlobalMux I__457 (
            .O(N__4649),
            .I(N__4646));
    gio2CtrlBuf I__456 (
            .O(N__4646),
            .I(C1_c_g));
    InMux I__455 (
            .O(N__4643),
            .I(N__4639));
    InMux I__454 (
            .O(N__4642),
            .I(N__4636));
    LocalMux I__453 (
            .O(N__4639),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__452 (
            .O(N__4636),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__451 (
            .O(N__4631),
            .I(N__4627));
    InMux I__450 (
            .O(N__4630),
            .I(N__4624));
    LocalMux I__449 (
            .O(N__4627),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__448 (
            .O(N__4624),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    CascadeMux I__447 (
            .O(N__4619),
            .I(N__4615));
    InMux I__446 (
            .O(N__4618),
            .I(N__4612));
    InMux I__445 (
            .O(N__4615),
            .I(N__4609));
    LocalMux I__444 (
            .O(N__4612),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__443 (
            .O(N__4609),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__442 (
            .O(N__4604),
            .I(N__4600));
    InMux I__441 (
            .O(N__4603),
            .I(N__4597));
    LocalMux I__440 (
            .O(N__4600),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__439 (
            .O(N__4597),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__438 (
            .O(N__4592),
            .I(N__4588));
    InMux I__437 (
            .O(N__4591),
            .I(N__4585));
    LocalMux I__436 (
            .O(N__4588),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__435 (
            .O(N__4585),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__434 (
            .O(N__4580),
            .I(N__4576));
    InMux I__433 (
            .O(N__4579),
            .I(N__4573));
    LocalMux I__432 (
            .O(N__4576),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__431 (
            .O(N__4573),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__430 (
            .O(N__4568),
            .I(N__4565));
    LocalMux I__429 (
            .O(N__4565),
            .I(N__4562));
    Span4Mux_v I__428 (
            .O(N__4562),
            .I(N__4559));
    Span4Mux_v I__427 (
            .O(N__4559),
            .I(N__4556));
    Sp12to4 I__426 (
            .O(N__4556),
            .I(N__4553));
    Odrv12 I__425 (
            .O(N__4553),
            .I(A_c_6));
    InMux I__424 (
            .O(N__4550),
            .I(N__4547));
    LocalMux I__423 (
            .O(N__4547),
            .I(N__4544));
    Span4Mux_v I__422 (
            .O(N__4544),
            .I(N__4541));
    Sp12to4 I__421 (
            .O(N__4541),
            .I(N__4538));
    Span12Mux_v I__420 (
            .O(N__4538),
            .I(N__4535));
    Odrv12 I__419 (
            .O(N__4535),
            .I(A_c_2));
    InMux I__418 (
            .O(N__4532),
            .I(N__4529));
    LocalMux I__417 (
            .O(N__4529),
            .I(N__4526));
    Span4Mux_v I__416 (
            .O(N__4526),
            .I(N__4523));
    Sp12to4 I__415 (
            .O(N__4523),
            .I(N__4520));
    Span12Mux_h I__414 (
            .O(N__4520),
            .I(N__4517));
    Span12Mux_v I__413 (
            .O(N__4517),
            .I(N__4514));
    Odrv12 I__412 (
            .O(N__4514),
            .I(A_c_3));
    InMux I__411 (
            .O(N__4511),
            .I(N__4508));
    LocalMux I__410 (
            .O(N__4508),
            .I(N__4505));
    Span4Mux_h I__409 (
            .O(N__4505),
            .I(N__4502));
    Sp12to4 I__408 (
            .O(N__4502),
            .I(N__4499));
    Span12Mux_v I__407 (
            .O(N__4499),
            .I(N__4496));
    Odrv12 I__406 (
            .O(N__4496),
            .I(A_c_4));
    IoInMux I__405 (
            .O(N__4493),
            .I(N__4490));
    LocalMux I__404 (
            .O(N__4490),
            .I(N__4487));
    Odrv12 I__403 (
            .O(N__4487),
            .I(DBRn_c_i_0));
    IoInMux I__402 (
            .O(N__4484),
            .I(N__4481));
    LocalMux I__401 (
            .O(N__4481),
            .I(N__4478));
    IoSpan4Mux I__400 (
            .O(N__4478),
            .I(N__4475));
    Span4Mux_s3_v I__399 (
            .O(N__4475),
            .I(N__4472));
    Odrv4 I__398 (
            .O(N__4472),
            .I(CLK80_PLL_i_i));
    InMux I__397 (
            .O(N__4469),
            .I(N__4466));
    LocalMux I__396 (
            .O(N__4466),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__395 (
            .O(N__4463),
            .I(bfn_6_7_0_));
    InMux I__394 (
            .O(N__4460),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__393 (
            .O(N__4457),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__392 (
            .O(N__4454),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__391 (
            .O(N__4451),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__390 (
            .O(N__4448),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    IoInMux I__389 (
            .O(N__4445),
            .I(N__4442));
    LocalMux I__388 (
            .O(N__4442),
            .I(N__4439));
    Span4Mux_s0_v I__387 (
            .O(N__4439),
            .I(N__4436));
    Span4Mux_v I__386 (
            .O(N__4436),
            .I(N__4433));
    Sp12to4 I__385 (
            .O(N__4433),
            .I(N__4430));
    Span12Mux_h I__384 (
            .O(N__4430),
            .I(N__4427));
    Span12Mux_v I__383 (
            .O(N__4427),
            .I(N__4424));
    Odrv12 I__382 (
            .O(N__4424),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__4670));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .I(N__4671));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__4672));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__4669));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__4667));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__4668));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .I(N__4666));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_12_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__8602),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7997),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4493),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__8237),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_6 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_11_6  (
            .in0(N__8155),
            .in1(N__11576),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_2_1_2.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_2_1_2.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_2_1_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_2_1_2 (
            .in0(N__11060),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_6_7_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_6_7_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_6_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(N__4469),
            .in2(_gnd_net_),
            .in3(N__4463),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__4673),
            .ce(),
            .sr(N__7553));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_6_7_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_6_7_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_6_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_6_7_1  (
            .in0(_gnd_net_),
            .in1(N__4631),
            .in2(_gnd_net_),
            .in3(N__4460),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__4673),
            .ce(),
            .sr(N__7553));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_6_7_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_6_7_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_6_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(N__4604),
            .in2(_gnd_net_),
            .in3(N__4457),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__4673),
            .ce(),
            .sr(N__7553));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_6_7_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_6_7_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_6_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_6_7_3  (
            .in0(_gnd_net_),
            .in1(N__4643),
            .in2(_gnd_net_),
            .in3(N__4454),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__4673),
            .ce(),
            .sr(N__7553));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_6_7_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_6_7_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_6_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(N__4618),
            .in2(_gnd_net_),
            .in3(N__4451),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__4673),
            .ce(),
            .sr(N__7553));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_6_7_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_6_7_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_6_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_6_7_5  (
            .in0(_gnd_net_),
            .in1(N__4580),
            .in2(_gnd_net_),
            .in3(N__4448),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__4673),
            .ce(),
            .sr(N__7553));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_6_7_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_6_7_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_6_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_6_7_6  (
            .in0(_gnd_net_),
            .in1(N__4592),
            .in2(_gnd_net_),
            .in3(N__4679),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__4673),
            .ce(),
            .sr(N__7553));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_6_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_6_7_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_6_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_6_7_7  (
            .in0(_gnd_net_),
            .in1(N__5269),
            .in2(_gnd_net_),
            .in3(N__4676),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4673),
            .ce(),
            .sr(N__7553));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_6_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_6_8_0 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_6_8_0  (
            .in0(N__4642),
            .in1(N__4630),
            .in2(N__4619),
            .in3(N__4603),
            .lcout(\U712_CHIP_RAM.REFRESH5lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_6_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_6_8_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_6_8_2  (
            .in0(_gnd_net_),
            .in1(N__4591),
            .in2(_gnd_net_),
            .in3(N__4579),
            .lcout(\U712_CHIP_RAM.REFRESH5lto7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_6_12_0.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_6_12_0.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_6_12_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_6_12_0 (
            .in0(N__4718),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_7_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_7_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_7_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_7_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4568),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11023),
            .ce(N__5026),
            .sr(N__11538));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_7_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_7_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_7_6_0  (
            .in0(N__4550),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11029),
            .ce(N__5022),
            .sr(N__11535));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_7_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_7_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4532),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11029),
            .ce(N__5022),
            .sr(N__11535));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_7_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_7_6_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__4511),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11029),
            .ce(N__5022),
            .sr(N__11535));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_7_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_7_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4766),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11029),
            .ce(N__5022),
            .sr(N__11535));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_7_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_7_6_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_7_6_4  (
            .in0(N__4748),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11029),
            .ce(N__5022),
            .sr(N__11535));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_7_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_7_7_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_7_7_0  (
            .in0(N__6723),
            .in1(N__10880),
            .in2(_gnd_net_),
            .in3(N__5708),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11035),
            .ce(N__4730),
            .sr(N__11529));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_8_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_8_0  (
            .in0(N__6140),
            .in1(N__5707),
            .in2(N__6548),
            .in3(N__6644),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11040),
            .ce(N__5720),
            .sr(N__11518));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_7_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_7_8_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(N__11575),
            .in2(_gnd_net_),
            .in3(N__4799),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_0_LC_7_14_4.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_7_14_4.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_7_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_7_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4714),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11055),
            .ce(),
            .sr(N__11488));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_4 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(N__8393),
            .in2(_gnd_net_),
            .in3(N__9075),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_5_1 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_5_1  (
            .in0(N__4958),
            .in1(N__5408),
            .in2(N__6209),
            .in3(N__5213),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11017),
            .ce(N__5553),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ8AQ_LC_8_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ8AQ_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ8AQ_LC_8_5_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ8AQ_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(N__6476),
            .in2(_gnd_net_),
            .in3(N__5801),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_8_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_8_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_8_5_4  (
            .in0(_gnd_net_),
            .in1(N__6370),
            .in2(_gnd_net_),
            .in3(N__7369),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_8_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_8_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4826),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11024),
            .ce(N__5027),
            .sr(N__11530));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI09RS_LC_8_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI09RS_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI09RS_LC_8_6_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI09RS_LC_8_6_6  (
            .in0(N__5743),
            .in1(N__6429),
            .in2(_gnd_net_),
            .in3(N__8997),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_7_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_8_7_1  (
            .in0(N__11573),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5120),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_8_7_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__11574),
            .in2(_gnd_net_),
            .in3(N__6046),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_8_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_8_7_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_8_7_5  (
            .in0(N__6129),
            .in1(N__6527),
            .in2(N__5339),
            .in3(N__6642),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11030),
            .ce(N__4808),
            .sr(N__11519));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_8_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_8_7_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_8_7_7  (
            .in0(N__6128),
            .in1(N__5353),
            .in2(N__6643),
            .in3(N__6526),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI722C3_1_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI722C3_1_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI722C3_1_LC_8_8_0 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI722C3_1_LC_8_8_0  (
            .in0(N__7139),
            .in1(N__11334),
            .in2(N__4793),
            .in3(N__4849),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_165_i_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI30J08_1_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI30J08_1_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI30J08_1_LC_8_8_1 .LUT_INIT=16'b0000010100001101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI30J08_1_LC_8_8_1  (
            .in0(N__11333),
            .in1(N__4862),
            .in2(N__4781),
            .in3(N__5227),
            .lcout(\U712_CHIP_RAM.N_90_i ),
            .ltout(\U712_CHIP_RAM.N_90_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_8_2 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_8_2  (
            .in0(N__4778),
            .in1(N__5114),
            .in2(N__4769),
            .in3(N__4838),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11036),
            .ce(N__5555),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_8_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_8_8_3 .LUT_INIT=16'b0000010000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_8_8_3  (
            .in0(N__7211),
            .in1(N__6523),
            .in2(N__7145),
            .in3(N__7318),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_298_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_8_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_8_8_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4868),
            .in3(N__5815),
            .lcout(\U712_CHIP_RAM.N_546 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIVFJO_LC_8_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIVFJO_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIVFJO_LC_8_8_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIVFJO_LC_8_8_5  (
            .in0(N__5745),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7317),
            .lcout(\U712_CHIP_RAM.N_300 ),
            .ltout(\U712_CHIP_RAM.N_300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_8_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_8_6  (
            .in0(N__6525),
            .in1(N__7131),
            .in2(N__4865),
            .in3(N__7212),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_0_0_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIPOTI1_LC_8_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIPOTI1_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIPOTI1_LC_8_8_7 .LUT_INIT=16'b0000001100011111;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIPOTI1_LC_8_8_7  (
            .in0(N__5744),
            .in1(N__6524),
            .in2(N__5816),
            .in3(N__7319),
            .lcout(\U712_CHIP_RAM.N_313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_8_9_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_8_9_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_8_9_4  (
            .in0(N__7030),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6977),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_8_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_8_9_5 .LUT_INIT=16'b1100110000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_8_9_5  (
            .in0(N__7320),
            .in1(N__7213),
            .in2(_gnd_net_),
            .in3(N__7132),
            .lcout(\U712_CHIP_RAM.N_310 ),
            .ltout(\U712_CHIP_RAM.N_310_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_9_6 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_9_6  (
            .in0(N__11332),
            .in1(N__5231),
            .in2(N__4853),
            .in3(N__4850),
            .lcout(\U712_CHIP_RAM.N_389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_8_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_5_LC_8_10_2  (
            .in0(N__11291),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4931),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11044),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_10_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_10_6  (
            .in0(N__4832),
            .in1(N__4930),
            .in2(_gnd_net_),
            .in3(N__5481),
            .lcout(\U712_CHIP_RAM.N_455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_8_10_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_4_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(N__11290),
            .in2(_gnd_net_),
            .in3(N__8024),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11044),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_8_11_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_8_11_2  (
            .in0(N__5080),
            .in1(N__5480),
            .in2(N__4904),
            .in3(N__5102),
            .lcout(),
            .ltout(\U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_8_11_3 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__4880),
            .in2(N__4922),
            .in3(N__8329),
            .lcout(\U712_CHIP_RAM.N_419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_8_12_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_8_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(N__5101),
            .in2(N__5068),
            .in3(N__5069),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_8_12_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_8_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(N__4879),
            .in2(_gnd_net_),
            .in3(N__4919),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_8_12_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_8_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__4903),
            .in2(_gnd_net_),
            .in3(N__4916),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_8_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_8_12_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__5081),
            .in2(_gnd_net_),
            .in3(N__4913),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_8_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_8_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_8_12_4 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_2_LC_8_12_4  (
            .in0(N__11251),
            .in1(N__4910),
            .in2(N__5501),
            .in3(N__8333),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11050),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_8_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_8_12_5 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_1_LC_8_12_5  (
            .in0(N__8330),
            .in1(N__5498),
            .in2(N__4889),
            .in3(N__11250),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11050),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_8_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_8_12_6 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_0_LC_8_12_6  (
            .in0(N__11249),
            .in1(N__5108),
            .in2(N__5500),
            .in3(N__8332),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11050),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_8_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_8_12_7 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_3_LC_8_12_7  (
            .in0(N__8331),
            .in1(N__5499),
            .in2(N__5090),
            .in3(N__11252),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11050),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_RNITKK4_1_LC_8_13_1.C_ON=1'b0;
    defparam DBR_SYNC_RNITKK4_1_LC_8_13_1.SEQ_MODE=4'b0000;
    defparam DBR_SYNC_RNITKK4_1_LC_8_13_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBR_SYNC_RNITKK4_1_LC_8_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8299),
            .lcout(DBR_SYNC_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_1_LC_8_14_4.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_8_14_4.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_8_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_8_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5051),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11053),
            .ce(),
            .sr(N__11484));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_9_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_9_4_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_9_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_9_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5045),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11005),
            .ce(N__5021),
            .sr(N__11536));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_5_3  (
            .in0(N__4982),
            .in1(N__4964),
            .in2(_gnd_net_),
            .in3(N__10541),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_6_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_6_0  (
            .in0(N__5132),
            .in1(N__11359),
            .in2(_gnd_net_),
            .in3(N__5806),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11018),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_6_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_6_1  (
            .in0(N__5354),
            .in1(N__6133),
            .in2(_gnd_net_),
            .in3(N__6478),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a3_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_178_i_LC_9_6_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_178_i_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_178_i_LC_9_6_2 .LUT_INIT=16'b0101000111110011;
    LogicCell40 \U712_BYTE_ENABLE.N_178_i_LC_9_6_2  (
            .in0(N__9002),
            .in1(N__5189),
            .in2(N__10775),
            .in3(N__5435),
            .lcout(N_178_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_176_i_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_176_i_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_176_i_LC_9_6_4 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \U712_BYTE_ENABLE.N_176_i_LC_9_6_4  (
            .in0(N__10689),
            .in1(N__5188),
            .in2(N__9035),
            .in3(N__5453),
            .lcout(N_176_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_6_5  (
            .in0(N__5159),
            .in1(N__5150),
            .in2(_gnd_net_),
            .in3(N__10554),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_6_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_6_7  (
            .in0(N__7373),
            .in1(N__8998),
            .in2(N__7240),
            .in3(N__6477),
            .lcout(\U712_CHIP_RAM.CPU_TACK_8_iv_i_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_7_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_9_7_0  (
            .in0(N__6085),
            .in1(N__7296),
            .in2(N__6776),
            .in3(N__6518),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_9_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_9_7_1  (
            .in0(N__6515),
            .in1(N__5798),
            .in2(_gnd_net_),
            .in3(N__7111),
            .lcout(\U712_CHIP_RAM.N_370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_9_7_2 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_9_7_2  (
            .in0(N__7110),
            .in1(_gnd_net_),
            .in2(N__7222),
            .in3(N__7294),
            .lcout(\U712_CHIP_RAM.N_464 ),
            .ltout(\U712_CHIP_RAM.N_464_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7TF5_2_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7TF5_2_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7TF5_2_LC_9_7_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7TF5_2_LC_9_7_3  (
            .in0(N__6516),
            .in1(N__5335),
            .in2(N__5126),
            .in3(N__6633),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_7_4 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_7_4  (
            .in0(N__5752),
            .in1(N__6517),
            .in2(N__5123),
            .in3(N__6675),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_7_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_9_7_5  (
            .in0(N__6519),
            .in1(N__11358),
            .in2(_gnd_net_),
            .in3(N__7112),
            .lcout(\U712_CHIP_RAM.N_390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIBERN2_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIBERN2_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIBERN2_LC_9_7_6 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNIBERN2_LC_9_7_6  (
            .in0(N__5799),
            .in1(N__6996),
            .in2(N__6775),
            .in3(N__7295),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIHSKQ_LC_9_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIHSKQ_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIHSKQ_LC_9_7_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIHSKQ_LC_9_7_7  (
            .in0(N__5635),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5294),
            .lcout(\U712_CHIP_RAM.N_461 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_9_8_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_9_8_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__7316),
            .in2(_gnd_net_),
            .in3(N__7406),
            .lcout(\U712_CHIP_RAM.N_551 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_8_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_8_1  (
            .in0(N__5405),
            .in1(N__7140),
            .in2(_gnd_net_),
            .in3(N__5216),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__11031),
            .ce(N__5554),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_9_8_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_9_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__6546),
            .in2(_gnd_net_),
            .in3(N__5204),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_8_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_8_3  (
            .in0(N__5406),
            .in1(N__7221),
            .in2(_gnd_net_),
            .in3(N__5201),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__11031),
            .ce(N__5554),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_8_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_8_4  (
            .in0(N__5402),
            .in1(N__5845),
            .in2(_gnd_net_),
            .in3(N__5198),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__11031),
            .ce(N__5554),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_8_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_8_5  (
            .in0(N__5407),
            .in1(N__5858),
            .in2(_gnd_net_),
            .in3(N__5195),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__11031),
            .ce(N__5554),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_8_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_8_6  (
            .in0(N__5403),
            .in1(N__5870),
            .in2(_gnd_net_),
            .in3(N__5192),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__11031),
            .ce(N__5554),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_8_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_8_7  (
            .in0(N__5831),
            .in1(N__5404),
            .in2(_gnd_net_),
            .in3(N__5375),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11031),
            .ce(N__5554),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_188_i_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_188_i_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_188_i_LC_9_9_1 .LUT_INIT=16'b0101000111110011;
    LogicCell40 \U712_BYTE_ENABLE.N_188_i_LC_9_9_1  (
            .in0(N__5444),
            .in1(N__7799),
            .in2(N__10771),
            .in3(N__9074),
            .lcout(N_188_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_9_2 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_9_2  (
            .in0(N__5289),
            .in1(N__5677),
            .in2(N__5628),
            .in3(N__5572),
            .lcout(\U712_CHIP_RAM.N_302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_0_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_0_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_0_LC_9_9_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_0_LC_9_9_3  (
            .in0(N__5571),
            .in1(N__5288),
            .in2(N__5696),
            .in3(N__5618),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_4 .LUT_INIT=16'b1100110000001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_4  (
            .in0(N__5703),
            .in1(N__11352),
            .in2(N__7001),
            .in3(N__5318),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11037),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__5290),
            .in2(_gnd_net_),
            .in3(N__9073),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_417_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_6 .LUT_INIT=16'b1100000011000100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_6  (
            .in0(N__8053),
            .in1(N__11351),
            .in2(N__5312),
            .in3(N__5309),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11037),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_9_9_7 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_9_9_7  (
            .in0(N__5273),
            .in1(N__5255),
            .in2(N__11360),
            .in3(N__5243),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11037),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_10_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_9_10_1  (
            .in0(N__11349),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5507),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11041),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_9_10_4 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_9_10_4  (
            .in0(N__10679),
            .in1(N__11348),
            .in2(_gnd_net_),
            .in3(N__10764),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11041),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_10_6 .LUT_INIT=16'b0010001100000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_10_6  (
            .in0(N__5491),
            .in1(N__5459),
            .in2(N__8344),
            .in3(N__11350),
            .lcout(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11041),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UUBE_i_o2_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_i_o2_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_i_o2_LC_9_11_2 .LUT_INIT=16'b1111000100011111;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_i_o2_LC_9_11_2  (
            .in0(N__9612),
            .in1(N__9766),
            .in2(N__9528),
            .in3(N__9702),
            .lcout(\U712_BYTE_ENABLE.N_326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_LC_9_11_7 .LUT_INIT=16'b1111100010101111;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_i_o2_LC_9_11_7  (
            .in0(N__9765),
            .in1(N__9611),
            .in2(N__9706),
            .in3(N__9515),
            .lcout(\U712_BYTE_ENABLE.N_323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_i_o2_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_i_o2_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_i_o2_LC_9_12_2 .LUT_INIT=16'b1011101101110101;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_i_o2_LC_9_12_2  (
            .in0(N__9475),
            .in1(N__9756),
            .in2(N__9623),
            .in3(N__9684),
            .lcout(\U712_BYTE_ENABLE.N_324 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_5_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_5_0  (
            .in0(N__5426),
            .in1(N__6035),
            .in2(_gnd_net_),
            .in3(N__10542),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_5_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_5_3  (
            .in0(N__7236),
            .in1(N__5805),
            .in2(N__6542),
            .in3(N__7368),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_6_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_6_0  (
            .in0(N__6194),
            .in1(N__6536),
            .in2(N__7241),
            .in3(N__7374),
            .lcout(\U712_CHIP_RAM.N_384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIR80N2_LC_10_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIR80N2_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIR80N2_LC_10_6_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIR80N2_LC_10_6_1  (
            .in0(N__11357),
            .in1(N__5800),
            .in2(_gnd_net_),
            .in3(N__6759),
            .lcout(\U712_CHIP_RAM.N_463 ),
            .ltout(\U712_CHIP_RAM.N_463_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_10_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_10_6_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(N__6535),
            .in2(N__5642),
            .in3(N__7146),
            .lcout(\U712_CHIP_RAM.N_550 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_10_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_10_6_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_10_6_3  (
            .in0(N__6131),
            .in1(N__5698),
            .in2(N__5639),
            .in3(N__6195),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_385_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_6_4 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_6_4  (
            .in0(N__6161),
            .in1(_gnd_net_),
            .in2(N__5600),
            .in3(N__6250),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_6_5 .LUT_INIT=16'b1100110100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_6_5  (
            .in0(N__5597),
            .in1(N__6818),
            .in2(N__5591),
            .in3(N__10548),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11010),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNICG3P2_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNICG3P2_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNICG3P2_LC_10_6_6 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNICG3P2_LC_10_6_6  (
            .in0(N__5588),
            .in1(N__6130),
            .in2(N__5582),
            .in3(N__6534),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0_a2_0 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_10_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_10_6_7 .LUT_INIT=16'b1100111111111111;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_10_6_7  (
            .in0(_gnd_net_),
            .in1(N__5697),
            .in2(N__5558),
            .in3(N__6193),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI36AQC_2_LC_10_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI36AQC_2_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI36AQC_2_LC_10_7_0 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI36AQC_2_LC_10_7_0  (
            .in0(N__6538),
            .in1(N__6191),
            .in2(N__5894),
            .in3(N__6132),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNINN3QI_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNINN3QI_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNINN3QI_LC_10_7_1 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNINN3QI_LC_10_7_1  (
            .in0(N__6192),
            .in1(N__5522),
            .in2(N__5510),
            .in3(N__5699),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_10_7_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__11338),
            .in2(_gnd_net_),
            .in3(N__6760),
            .lcout(\U712_CHIP_RAM.N_533 ),
            .ltout(\U712_CHIP_RAM.N_533_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_3_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_3_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_3_LC_10_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_3_LC_10_7_3  (
            .in0(N__7363),
            .in1(N__7214),
            .in2(N__5906),
            .in3(N__5903),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_391_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIEVI78_3_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIEVI78_3_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIEVI78_3_LC_10_7_4 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIEVI78_3_LC_10_7_4  (
            .in0(_gnd_net_),
            .in1(N__6190),
            .in2(N__5897),
            .in3(N__6084),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_10_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_10_7_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_10_7_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_LC_10_7_5  (
            .in0(N__6761),
            .in1(N__6539),
            .in2(N__7375),
            .in3(N__6086),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11019),
            .ce(N__6656),
            .sr(N__11505));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_7_6  (
            .in0(N__5869),
            .in1(N__5857),
            .in2(N__5846),
            .in3(N__5830),
            .lcout(\U712_CHIP_RAM.N_295 ),
            .ltout(\U712_CHIP_RAM.N_295_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_7_7 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5819),
            .in3(N__5797),
            .lcout(\U712_CHIP_RAM.N_458 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNILJ788_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNILJ788_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNILJ788_LC_10_8_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNILJ788_LC_10_8_0  (
            .in0(N__6978),
            .in1(N__6696),
            .in2(N__7362),
            .in3(N__7407),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_10_8_1 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_10_8_1  (
            .in0(N__6531),
            .in1(N__6676),
            .in2(N__5759),
            .in3(N__5756),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_8_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5723),
            .in3(N__11571),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_8_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_8_3  (
            .in0(N__5678),
            .in1(N__6125),
            .in2(N__6547),
            .in3(N__6623),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIF4EE6_2_LC_10_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIF4EE6_2_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIF4EE6_2_LC_10_8_4 .LUT_INIT=16'b1111000000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIF4EE6_2_LC_10_8_4  (
            .in0(N__6126),
            .in1(N__6533),
            .in2(N__6251),
            .in3(N__6157),
            .lcout(\U712_CHIP_RAM.N_441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_10_8_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_10_8_5  (
            .in0(N__6532),
            .in1(N__6127),
            .in2(_gnd_net_),
            .in3(N__6768),
            .lcout(\U712_CHIP_RAM.DBENn_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_8_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_8_6  (
            .in0(N__7201),
            .in1(N__7109),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_465 ),
            .ltout(\U712_CHIP_RAM.N_465_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_10_8_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_3_LC_10_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6068),
            .in3(N__6622),
            .lcout(\U712_CHIP_RAM.N_469 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_9_0 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_10_9_0  (
            .in0(N__6065),
            .in1(N__6034),
            .in2(N__11837),
            .in3(N__6050),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11032),
            .ce(),
            .sr(N__11492));
    defparam \U712_CHIP_RAM.DBENn_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_10_9_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_10_9_1 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_10_9_1  (
            .in0(N__6020),
            .in1(N__7022),
            .in2(N__6014),
            .in3(N__10178),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11032),
            .ce(),
            .sr(N__11492));
    defparam \U712_CHIP_RAM.DBDIR_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_10_9_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_10_9_3 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_10_9_3  (
            .in0(N__6731),
            .in1(N__5986),
            .in2(_gnd_net_),
            .in3(N__6697),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11032),
            .ce(),
            .sr(N__11492));
    defparam pll_RNI8MQ3_LC_10_10_1.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_10_10_1.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_10_10_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 pll_RNI8MQ3_LC_10_10_1 (
            .in0(N__7718),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.N_167_i_LC_10_19_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_167_i_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_167_i_LC_10_19_2 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \U712_BUFFERS.N_167_i_LC_10_19_2  (
            .in0(N__10807),
            .in1(N__10667),
            .in2(_gnd_net_),
            .in3(N__10762),
            .lcout(N_167_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_11_3_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_3_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_3_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_3_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_4_4  (
            .in0(N__6337),
            .in1(N__6302),
            .in2(_gnd_net_),
            .in3(N__10586),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_5  (
            .in0(N__10587),
            .in1(N__9084),
            .in2(N__6290),
            .in3(N__10139),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_11_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_11_5_6 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_11_5_6  (
            .in0(N__6994),
            .in1(N__6268),
            .in2(N__7376),
            .in3(N__7385),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11002),
            .ce(),
            .sr(N__11511));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_6_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_6_3  (
            .in0(N__10502),
            .in1(N__9163),
            .in2(N__12174),
            .in3(N__10411),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_6_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_6_6  (
            .in0(N__6257),
            .in1(N__6249),
            .in2(N__6569),
            .in3(N__6220),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_296_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_6_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__6819),
            .in2(N__6230),
            .in3(N__9164),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11006),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_11_7_1 .LUT_INIT=16'b1010101000000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_11_7_1  (
            .in0(N__12173),
            .in1(N__6797),
            .in2(N__6227),
            .in3(N__6821),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11011),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_11_7_2  (
            .in0(N__6541),
            .in1(N__7148),
            .in2(N__6205),
            .in3(N__7367),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_442_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_7_3 .LUT_INIT=16'b1000100010001011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_7_3  (
            .in0(N__10421),
            .in1(N__6820),
            .in2(N__6800),
            .in3(N__6796),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11011),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_7_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__6788),
            .in2(_gnd_net_),
            .in3(N__6767),
            .lcout(\U712_CHIP_RAM.N_428 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_11_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_11_7_7 .LUT_INIT=16'b0101000011000000;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_11_7_7  (
            .in0(N__6727),
            .in1(N__10788),
            .in2(N__11356),
            .in3(N__6698),
            .lcout(DMA_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11011),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_11_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_11_8_0 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_11_8_0  (
            .in0(N__6540),
            .in1(N__6634),
            .in2(N__7052),
            .in3(N__6680),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_11_8_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6659),
            .in3(N__11570),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_8_2 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_8_2  (
            .in0(N__7051),
            .in1(N__6635),
            .in2(N__6386),
            .in3(N__6593),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_11_8_3 .LUT_INIT=16'b1100101011111010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_11_8_3  (
            .in0(N__7754),
            .in1(N__6581),
            .in2(N__6572),
            .in3(N__7144),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11020),
            .ce(),
            .sr(N__11493));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_2_LC_11_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_2_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_2_LC_11_8_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_2_LC_11_8_4  (
            .in0(N__6562),
            .in1(N__6537),
            .in2(_gnd_net_),
            .in3(N__7408),
            .lcout(\U712_CHIP_RAM.N_438 ),
            .ltout(\U712_CHIP_RAM.N_438_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_11_8_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_11_8_5  (
            .in0(N__7409),
            .in1(N__6997),
            .in2(N__7388),
            .in3(N__7338),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIREK92_3_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIREK92_3_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIREK92_3_LC_11_8_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIREK92_3_LC_11_8_7  (
            .in0(N__7334),
            .in1(N__7226),
            .in2(N__7147),
            .in3(N__7064),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_9_2 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_9_2  (
            .in0(N__7844),
            .in1(N__7860),
            .in2(_gnd_net_),
            .in3(N__7753),
            .lcout(\U712_CYCLE_TERM.N_321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_11_9_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_11_9_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_11_9_7  (
            .in0(N__7023),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6995),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_11_10_0 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_LC_11_10_0  (
            .in0(N__7877),
            .in1(N__6884),
            .in2(_gnd_net_),
            .in3(N__6935),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11033),
            .ce(),
            .sr(N__11489));
    defparam \U712_BYTE_ENABLE.LMBE_i_o2_LC_11_11_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LMBE_i_o2_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LMBE_i_o2_LC_11_11_1 .LUT_INIT=16'b1111001000101111;
    LogicCell40 \U712_BYTE_ENABLE.LMBE_i_o2_LC_11_11_1  (
            .in0(N__9767),
            .in1(N__9624),
            .in2(N__9707),
            .in3(N__9519),
            .lcout(\U712_BYTE_ENABLE.N_325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_4_0 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_12_4_0  (
            .in0(N__9368),
            .in1(N__11921),
            .in2(N__9329),
            .in3(N__6866),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11001),
            .ce(N__9244),
            .sr(N__11510));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_2  (
            .in0(N__10599),
            .in1(N__6845),
            .in2(_gnd_net_),
            .in3(N__6833),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_3  (
            .in0(N__9083),
            .in1(N__10600),
            .in2(N__6824),
            .in3(N__8618),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_5_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_5_7  (
            .in0(N__7583),
            .in1(N__7568),
            .in2(_gnd_net_),
            .in3(N__10598),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_12_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_12_6_0 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_12_6_0  (
            .in0(N__10549),
            .in1(N__12166),
            .in2(N__10422),
            .in3(N__7546),
            .lcout(\U712_CHIP_RAM.un1_CMA25_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_6_1  (
            .in0(N__7528),
            .in1(N__7505),
            .in2(_gnd_net_),
            .in3(N__10550),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_2  (
            .in0(N__10551),
            .in1(N__9081),
            .in2(N__7496),
            .in3(N__8702),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_6_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_12_6_5  (
            .in0(N__7474),
            .in1(N__7454),
            .in2(_gnd_net_),
            .in3(N__10552),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_6_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_6_6  (
            .in0(N__10415),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9165),
            .lcout(\U712_CHIP_RAM.N_305 ),
            .ltout(\U712_CHIP_RAM.N_305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_7 .LUT_INIT=16'b0100000000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_7  (
            .in0(N__9082),
            .in1(N__10267),
            .in2(N__7445),
            .in3(N__10553),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_7_2  (
            .in0(N__9079),
            .in1(N__7442),
            .in2(_gnd_net_),
            .in3(N__8720),
            .lcout(\U712_CHIP_RAM.N_346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_7_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_7_7  (
            .in0(N__7421),
            .in1(N__9080),
            .in2(_gnd_net_),
            .in3(N__8681),
            .lcout(\U712_CHIP_RAM.N_352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_186_i_LC_12_8_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_186_i_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_186_i_LC_12_8_2 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \U712_BYTE_ENABLE.N_186_i_LC_12_8_2  (
            .in0(N__10691),
            .in1(N__7798),
            .in2(N__7784),
            .in3(N__9085),
            .lcout(N_186_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_9_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_9_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__7845),
            .in2(_gnd_net_),
            .in3(N__7751),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_12_9_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_12_9_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_12_9_2  (
            .in0(N__7709),
            .in1(N__11245),
            .in2(_gnd_net_),
            .in3(N__7908),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11016),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_9_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_9_3 .LUT_INIT=16'b0000010100010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_9_3  (
            .in0(N__7907),
            .in1(N__7846),
            .in2(N__7865),
            .in3(N__7752),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_450_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_9_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_9_4 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_12_9_4  (
            .in0(N__7710),
            .in1(N__7864),
            .in2(N__7733),
            .in3(N__11244),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11016),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_12_9_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_12_9_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_12_9_5  (
            .in0(N__11246),
            .in1(_gnd_net_),
            .in2(N__7730),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11016),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_12_9_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_12_9_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(N__7665),
            .in2(_gnd_net_),
            .in3(N__7726),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_12_9_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_12_9_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_12_9_7  (
            .in0(N__11247),
            .in1(_gnd_net_),
            .in2(N__7670),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11016),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_12_10_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_12_10_1 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_12_10_1 .LUT_INIT=16'b1111111111000100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_12_10_1  (
            .in0(N__7910),
            .in1(N__7601),
            .in2(N__7714),
            .in3(N__7669),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11022),
            .ce(),
            .sr(N__11483));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_12_10_3 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_12_10_3 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_12_10_3  (
            .in0(N__7909),
            .in1(N__7892),
            .in2(N__7886),
            .in3(N__7876),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11022),
            .ce(),
            .sr(N__11483));
    defparam \U712_REG_SM.REG_TACK_LC_12_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_12_10_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_12_10_5  (
            .in0(N__8015),
            .in1(N__7847),
            .in2(N__8354),
            .in3(N__7826),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11022),
            .ce(),
            .sr(N__11483));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_12_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_12_10_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_12_10_6 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_12_10_6  (
            .in0(N__9983),
            .in1(N__8360),
            .in2(_gnd_net_),
            .in3(N__8915),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11022),
            .ce(),
            .sr(N__11483));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_12_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_12_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_12_11_3  (
            .in0(N__11194),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7805),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11025),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_12_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_12_11_4 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_12_11_4  (
            .in0(N__8889),
            .in1(N__7819),
            .in2(N__9979),
            .in3(N__8913),
            .lcout(\U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_7_LC_12_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_7_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_7_LC_12_11_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_7_LC_12_11_5  (
            .in0(N__11196),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7811),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11025),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_12_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_12_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__11195),
            .in2(_gnd_net_),
            .in3(N__7820),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11025),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_12_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_12_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_12_11_7  (
            .in0(N__11193),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8014),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11025),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_12_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_12_12_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_12_12_2  (
            .in0(N__10030),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8334),
            .lcout(\U712_REG_SM.N_320 ),
            .ltout(\U712_REG_SM.N_320_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_12_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_12_12_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_12_12_3  (
            .in0(N__8250),
            .in1(N__9978),
            .in2(N__8000),
            .in3(N__12304),
            .lcout(\U712_REG_SM.N_409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_7.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_7.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11248),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_5_3 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_5_3  (
            .in0(N__9119),
            .in1(N__7985),
            .in2(N__10370),
            .in3(N__10605),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_5_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_5_4  (
            .in0(N__10601),
            .in1(N__9120),
            .in2(N__7979),
            .in3(N__10127),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_13_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_13_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_13_5_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_13_5_5  (
            .in0(N__11572),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7964),
            .lcout(\U712_CHIP_RAM.un1_CMA25_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_13_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_13_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_13_5_6 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_13_5_6  (
            .in0(N__7958),
            .in1(N__9121),
            .in2(N__10612),
            .in3(N__8126),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_6_1 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_6_1  (
            .in0(N__9115),
            .in1(N__7949),
            .in2(N__10597),
            .in3(N__8690),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_6_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__7916),
            .in2(N__7943),
            .in3(N__7940),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11007),
            .ce(N__9250),
            .sr(N__11506));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_6_4 .LUT_INIT=16'b1101110111010101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_6_4  (
            .in0(N__10562),
            .in1(N__9355),
            .in2(N__9123),
            .in3(N__10268),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_7_0 .LUT_INIT=16'b1000111110000011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_13_7_0  (
            .in0(N__8189),
            .in1(N__9359),
            .in2(N__10616),
            .in3(N__8183),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11012),
            .ce(N__9240),
            .sr(N__11499));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_8_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_8_0  (
            .in0(N__11831),
            .in1(N__8156),
            .in2(N__11906),
            .in3(N__8125),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .ce(),
            .sr(N__11494));
    defparam \U712_BUFFERS.N_169_i_LC_13_9_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_169_i_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_169_i_LC_13_9_1 .LUT_INIT=16'b0000000011101010;
    LogicCell40 \U712_BUFFERS.N_169_i_LC_13_9_1  (
            .in0(N__9122),
            .in1(N__10690),
            .in2(N__10763),
            .in3(N__8386),
            .lcout(N_169_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_13_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_13_10_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__8935),
            .in2(_gnd_net_),
            .in3(N__8858),
            .lcout(),
            .ltout(\U712_REG_SM.N_397_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_13_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_13_10_3 .LUT_INIT=16'b1010000010100010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_13_10_3  (
            .in0(N__11301),
            .in1(N__8087),
            .in2(N__8063),
            .in3(N__8060),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11034),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_13_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_13_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_13_10_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_3_LC_13_10_7  (
            .in0(N__11300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10166),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11034),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIJUGT_3_LC_13_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIJUGT_3_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIJUGT_3_LC_13_11_0 .LUT_INIT=16'b0000100000001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIJUGT_3_LC_13_11_0  (
            .in0(N__10038),
            .in1(N__8275),
            .in2(N__12324),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.N_548 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_13_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_13_11_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__12297),
            .in2(_gnd_net_),
            .in3(N__10037),
            .lcout(\U712_REG_SM.N_319 ),
            .ltout(\U712_REG_SM.N_319_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_13_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_13_11_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_1_LC_13_11_2  (
            .in0(N__9883),
            .in1(N__8378),
            .in2(N__8003),
            .in3(N__9963),
            .lcout(),
            .ltout(\U712_REG_SM.REG_CYCLE_5_iv_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_13_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_13_11_3 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_13_11_3  (
            .in0(N__8379),
            .in1(N__11192),
            .in2(N__8402),
            .in3(N__8399),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11038),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_13_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_13_11_5 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_13_11_5  (
            .in0(N__8861),
            .in1(N__10039),
            .in2(N__12325),
            .in3(N__8888),
            .lcout(\U712_REG_SM.STATE_COUNTsr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_13_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_13_11_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_13_11_6  (
            .in0(N__9882),
            .in1(N__8274),
            .in2(_gnd_net_),
            .in3(N__9962),
            .lcout(\U712_REG_SM.N_328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_13_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_13_12_0 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_13_12_0  (
            .in0(N__10031),
            .in1(N__8276),
            .in2(N__8345),
            .in3(N__8251),
            .lcout(),
            .ltout(\U712_REG_SM.N_412_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_13_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_13_12_1 .LUT_INIT=16'b0000100000001010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_13_12_1  (
            .in0(N__11317),
            .in1(N__12307),
            .in2(N__8279),
            .in3(N__10033),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11042),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_13_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_13_12_5 .LUT_INIT=16'b1111010111000101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_13_12_5  (
            .in0(N__8252),
            .in1(N__12305),
            .in2(N__10082),
            .in3(N__10032),
            .lcout(),
            .ltout(\U712_REG_SM.N_360_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_13_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_13_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_13_12_6 .LUT_INIT=16'b0000110000000100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_13_12_6  (
            .in0(N__12306),
            .in1(N__11316),
            .in2(N__8261),
            .in3(N__8258),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11042),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_0_LC_13_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_13_13_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_13_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8224),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11045),
            .ce(),
            .sr(N__11479));
    defparam \U712_REG_SM.C3_SYNC_1_LC_13_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_13_13_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_13_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8195),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11045),
            .ce(),
            .sr(N__11479));
    defparam \U712_REG_SM.C1_SYNC_1_LC_13_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_13_14_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_13_14_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_13_14_4  (
            .in0(_gnd_net_),
            .in1(N__8567),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11049),
            .ce(),
            .sr(N__11478));
    defparam \U712_REG_SM.C1_SYNC_0_LC_13_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_13_15_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_13_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8603),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11051),
            .ce(),
            .sr(N__11477));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_4_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_4_2 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_14_4_2  (
            .in0(N__9390),
            .in1(N__9311),
            .in2(N__10115),
            .in3(N__8561),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11003),
            .ce(N__9249),
            .sr(N__11531));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_4_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_4_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_14_4_3  (
            .in0(N__12184),
            .in1(N__9391),
            .in2(_gnd_net_),
            .in3(N__10610),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11003),
            .ce(N__9249),
            .sr(N__11531));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_4_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_14_4_7 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_14_4_7  (
            .in0(N__8711),
            .in1(N__9392),
            .in2(N__9326),
            .in3(N__8513),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11003),
            .ce(N__9249),
            .sr(N__11531));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_5_0 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_14_5_0  (
            .in0(N__10151),
            .in1(N__9388),
            .in2(N__9328),
            .in3(N__8486),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11008),
            .ce(N__9245),
            .sr(N__11520));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_5_1 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_14_5_1  (
            .in0(N__9386),
            .in1(N__8729),
            .in2(N__9325),
            .in3(N__8456),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11008),
            .ce(N__9245),
            .sr(N__11520));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_14_5_4 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_14_5_4  (
            .in0(N__12026),
            .in1(N__9387),
            .in2(N__9327),
            .in3(N__8426),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11008),
            .ce(N__9245),
            .sr(N__11520));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_14_6_1  (
            .in0(N__9140),
            .in1(N__8771),
            .in2(N__9125),
            .in3(N__11660),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11013),
            .ce(N__9251),
            .sr(N__11512));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_1  (
            .in0(N__10313),
            .in1(N__11757),
            .in2(_gnd_net_),
            .in3(N__10353),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11648),
            .ce(N__11612),
            .sr(N__11507));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_4  (
            .in0(N__10354),
            .in1(N__11759),
            .in2(_gnd_net_),
            .in3(N__8668),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11648),
            .ce(N__11612),
            .sr(N__11507));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_7  (
            .in0(N__8669),
            .in1(N__11758),
            .in2(_gnd_net_),
            .in3(N__12122),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11648),
            .ce(N__11612),
            .sr(N__11507));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_8_1  (
            .in0(N__11760),
            .in1(N__12005),
            .in2(_gnd_net_),
            .in3(N__10249),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__11610),
            .sr(N__11500));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_8_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_8_2  (
            .in0(N__12006),
            .in1(N__11761),
            .in2(_gnd_net_),
            .in3(N__11965),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__11610),
            .sr(N__11500));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_8_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_8_7  (
            .in0(N__8666),
            .in1(N__11827),
            .in2(_gnd_net_),
            .in3(N__12121),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__11610),
            .sr(N__11500));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_9_7  (
            .in0(N__11812),
            .in1(N__8667),
            .in2(_gnd_net_),
            .in3(N__10352),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__11609),
            .sr(N__11495));
    defparam \U712_REG_SM.REGENn_LC_14_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_14_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_14_10_0 .LUT_INIT=16'b1100011011000100;
    LogicCell40 \U712_REG_SM.REGENn_LC_14_10_0  (
            .in0(N__8792),
            .in1(N__8811),
            .in2(N__12332),
            .in3(N__8896),
            .lcout(BLSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11039),
            .ce(),
            .sr(N__11490));
    defparam \U712_REG_SM.START_RST_LC_14_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_14_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_14_10_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \U712_REG_SM.START_RST_LC_14_10_6  (
            .in0(N__10078),
            .in1(N__8936),
            .in2(_gnd_net_),
            .in3(N__10099),
            .lcout(\U712_REG_SM.START_RSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11039),
            .ce(),
            .sr(N__11490));
    defparam \U712_REG_SM.STATE_COUNT_8_LC_14_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_8_LC_14_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_8_LC_14_11_1 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_8_LC_14_11_1  (
            .in0(N__8924),
            .in1(N__11265),
            .in2(N__9977),
            .in3(N__8914),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11043),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_14_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_14_11_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_14_11_2  (
            .in0(N__8859),
            .in1(N__10041),
            .in2(N__12329),
            .in3(N__8897),
            .lcout(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_14_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_14_11_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_14_11_3  (
            .in0(N__10042),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12314),
            .lcout(),
            .ltout(\U712_REG_SM.N_318_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_14_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_14_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_14_11_4 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_14_11_4  (
            .in0(N__11264),
            .in1(N__10100),
            .in2(N__8864),
            .in3(N__10079),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11043),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_RNO_0_LC_14_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_RNO_0_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REGENn_RNO_0_LC_14_11_6 .LUT_INIT=16'b0011000001000100;
    LogicCell40 \U712_REG_SM.REGENn_RNO_0_LC_14_11_6  (
            .in0(N__8860),
            .in1(N__10040),
            .in2(N__10081),
            .in3(N__8810),
            .lcout(\U712_REG_SM.REGENn_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDSn_RNO_0_LC_14_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_14_14_1 .LUT_INIT=16'b0000001000001000;
    LogicCell40 \U712_REG_SM.UDSn_RNO_0_LC_14_14_1  (
            .in0(N__9614),
            .in1(N__9532),
            .in2(N__10888),
            .in3(N__9683),
            .lcout(\U712_REG_SM.N_400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_RNO_0_LC_14_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_14_15_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_REG_SM.LDSn_RNO_0_LC_14_15_4  (
            .in0(N__10870),
            .in1(N__9613),
            .in2(N__9533),
            .in3(N__9682),
            .lcout(\U712_REG_SM.N_398 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_326_i_LC_14_20_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_326_i_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_326_i_LC_14_20_1 .LUT_INIT=16'b0101101001001000;
    LogicCell40 \U712_BYTE_ENABLE.N_326_i_LC_14_20_1  (
            .in0(N__9681),
            .in1(N__9755),
            .in2(N__9521),
            .in3(N__9622),
            .lcout(N_326_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_325_i_LC_14_20_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_325_i_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_325_i_LC_14_20_3 .LUT_INIT=16'b0101101000010010;
    LogicCell40 \U712_BYTE_ENABLE.N_325_i_LC_14_20_3  (
            .in0(N__9680),
            .in1(N__9754),
            .in2(N__9520),
            .in3(N__9621),
            .lcout(N_325_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_323_i_LC_14_20_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_323_i_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_323_i_LC_14_20_4 .LUT_INIT=16'b0001001101000100;
    LogicCell40 \U712_BYTE_ENABLE.N_323_i_LC_14_20_4  (
            .in0(N__9752),
            .in1(N__9678),
            .in2(N__9625),
            .in3(N__9502),
            .lcout(N_323_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_324_i_LC_14_20_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_324_i_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_324_i_LC_14_20_6 .LUT_INIT=16'b0010001110001000;
    LogicCell40 \U712_BYTE_ENABLE.N_324_i_LC_14_20_6  (
            .in0(N__9753),
            .in1(N__9679),
            .in2(N__9626),
            .in3(N__9503),
            .lcout(N_324_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WEn_LC_15_3_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_15_3_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_15_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_15_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9179),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11004),
            .ce(),
            .sr(N__11539));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_15_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_15_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_15_4_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_15_4_3  (
            .in0(_gnd_net_),
            .in1(N__9108),
            .in2(_gnd_net_),
            .in3(N__10609),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_15_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_15_5_2 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_15_5_2  (
            .in0(N__9389),
            .in1(N__8945),
            .in2(N__9324),
            .in3(N__8951),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11014),
            .ce(N__9233),
            .sr(N__11532));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_15_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_15_6_2 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_15_6_2  (
            .in0(N__10429),
            .in1(N__10560),
            .in2(_gnd_net_),
            .in3(N__9178),
            .lcout(\U712_CHIP_RAM.CMA_5_i_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_15_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_15_6_6 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_15_6_6  (
            .in0(N__9134),
            .in1(N__10561),
            .in2(N__9124),
            .in3(N__10274),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_1  (
            .in0(N__11799),
            .in1(N__10312),
            .in2(_gnd_net_),
            .in3(N__11969),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11647),
            .ce(N__11615),
            .sr(N__11513));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_7  (
            .in0(N__12071),
            .in1(N__11800),
            .in2(_gnd_net_),
            .in3(N__11902),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11647),
            .ce(N__11615),
            .sr(N__11513));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_8_1  (
            .in0(N__11823),
            .in1(N__10305),
            .in2(_gnd_net_),
            .in3(N__11964),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__11613),
            .sr(N__11508));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_8_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_8_7  (
            .in0(N__11895),
            .in1(_gnd_net_),
            .in2(N__11836),
            .in3(N__12070),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__11613),
            .sr(N__11508));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_9_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_9_2  (
            .in0(N__10202),
            .in1(N__11811),
            .in2(_gnd_net_),
            .in3(N__10239),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11643),
            .ce(N__11611),
            .sr(N__11501));
    defparam \U712_REG_SM.WRITE_CYCLE_LC_15_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_15_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_15_11_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_REG_SM.WRITE_CYCLE_LC_15_11_7  (
            .in0(N__10889),
            .in1(N__9878),
            .in2(_gnd_net_),
            .in3(N__10098),
            .lcout(\U712_REG_SM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11046),
            .ce(),
            .sr(N__11491));
    defparam \U712_REG_SM.STATE_COUNT_RNI3HF31_1_LC_15_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI3HF31_1_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI3HF31_1_LC_15_13_2 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI3HF31_1_LC_15_13_2  (
            .in0(N__10080),
            .in1(N__12320),
            .in2(N__10043),
            .in3(N__9967),
            .lcout(\U712_REG_SM.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDSn_LC_15_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_15_14_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_15_14_2 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \U712_REG_SM.UDSn_LC_15_14_2  (
            .in0(N__12318),
            .in1(N__9920),
            .in2(N__9901),
            .in3(N__12357),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11052),
            .ce(),
            .sr(N__11481));
    defparam \U712_REG_SM.PRnW_LC_15_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.PRnW_LC_15_14_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.PRnW_LC_15_14_5 .LUT_INIT=16'b1101111111010000;
    LogicCell40 \U712_REG_SM.PRnW_LC_15_14_5  (
            .in0(N__9884),
            .in1(N__12319),
            .in2(N__12359),
            .in3(N__9844),
            .lcout(PRnW_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11052),
            .ce(),
            .sr(N__11481));
    defparam \U712_REG_SM.LDSn_LC_15_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_15_15_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_15_15_0 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \U712_REG_SM.LDSn_LC_15_15_0  (
            .in0(N__9833),
            .in1(N__12358),
            .in2(N__9817),
            .in3(N__12330),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11054),
            .ce(),
            .sr(N__11480));
    defparam \U712_CHIP_RAM.CASn_LC_16_3_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_16_3_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_16_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_16_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10611),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11009),
            .ce(),
            .sr(N__11544));
    defparam \U712_CHIP_RAM.RASn_LC_16_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_16_4_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_16_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_16_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10433),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11015),
            .ce(),
            .sr(N__11540));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_16_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_16_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_16_6_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_16_6_4  (
            .in0(N__12069),
            .in1(N__11835),
            .in2(_gnd_net_),
            .in3(N__12119),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__11619),
            .sr(N__11533));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_16_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_16_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_16_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_16_7_2  (
            .in0(N__11798),
            .in1(N__10355),
            .in2(_gnd_net_),
            .in3(N__10304),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__11617),
            .sr(N__11521));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_16_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_16_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_16_8_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_16_8_7  (
            .in0(N__12013),
            .in1(N__11819),
            .in2(_gnd_net_),
            .in3(N__10250),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11644),
            .ce(N__11616),
            .sr(N__11514));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_16_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_16_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_16_9_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_16_9_1  (
            .in0(N__10238),
            .in1(N__11801),
            .in2(_gnd_net_),
            .in3(N__10201),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__11614),
            .sr(N__11509));
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_16_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_16_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_16_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_2_LC_16_10_0  (
            .in0(N__11243),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10157),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11047),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_16_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_16_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_16_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_16_10_2  (
            .in0(N__11242),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11066),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11047),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_RNO_LC_16_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_16_14_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_REG_SM.ASn_ess_RNO_LC_16_14_0  (
            .in0(N__11569),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12350),
            .lcout(\U712_REG_SM.N_152_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_LC_16_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_LC_16_15_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_ess_LC_16_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.ASn_ess_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12331),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11056),
            .ce(N__12197),
            .sr(N__11482));
    defparam \U712_CHIP_RAM.CRCSn_LC_17_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_17_4_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_17_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_17_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12185),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11021),
            .ce(),
            .sr(N__11545));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_6_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_6_4  (
            .in0(N__12120),
            .in1(N__11830),
            .in2(_gnd_net_),
            .in3(N__12068),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11646),
            .ce(N__11621),
            .sr(N__11537));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_17_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_17_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_17_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_17_7_7  (
            .in0(N__12014),
            .in1(N__11829),
            .in2(_gnd_net_),
            .in3(N__11947),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11645),
            .ce(N__11620),
            .sr(N__11534));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_8_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_8_4  (
            .in0(N__11885),
            .in1(N__11828),
            .in2(_gnd_net_),
            .in3(N__11089),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11642),
            .ce(N__11618),
            .sr(N__11522));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_9_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_17_9_7  (
            .in0(N__11263),
            .in1(N__11105),
            .in2(_gnd_net_),
            .in3(N__11093),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11048),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_0 .LUT_INIT=16'b0101001100110011;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_0  (
            .in0(N__10887),
            .in1(N__10808),
            .in2(N__10727),
            .in3(N__10666),
            .lcout(N_362),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

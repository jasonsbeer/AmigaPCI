-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 13 2025 15:27:47

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U400_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U400_TOP
entity U400_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    MA : out std_logic_vector(12 downto 0);
    A : in std_logic_vector(31 downto 0);
    LBENn : out std_logic;
    CS0n : out std_logic;
    UUBEn : out std_logic;
    TAn : out std_logic;
    CLK40 : in std_logic;
    RnW : in std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    WEn : out std_logic;
    LLBEn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    RASn : out std_logic;
    CS1n : out std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic);
end U400_TOP;

-- Architecture of U400_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U400_TOP is

signal \N__7125\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \CLK40_ibuf_gb_io_gb_input\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_28\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CONFIGUREDC_net\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a2_1_0_0_cascade_\ : std_logic;
signal \bfn_4_5_0_\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_1\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_2\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_3\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_4\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_5\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_6\ : std_logic;
signal \U400_SDRAM.un2_REFRESH_COUNTER_cry_7\ : std_logic;
signal \INVU400_SDRAM.REFRESH_COUNTER_2C_net\ : std_logic;
signal \bfn_4_6_0_\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_2C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_0_0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a2_1_0_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U400_SDRAM.N_97_cascade_\ : std_logic;
signal \U400_SDRAM.N_256_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \CS0n_c\ : std_logic;
signal \INVU400_SDRAM.CS0nC_net\ : std_logic;
signal \CASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \INVU400_SDRAM.CASnC_net\ : std_logic;
signal \RASn_c\ : std_logic;
signal \INVU400_SDRAM.RASnC_net\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_18\ : std_logic;
signal \MA_c_8\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_17\ : std_logic;
signal \MA_c_7\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_8C_net\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_16\ : std_logic;
signal \MA_c_6\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_6C_net\ : std_logic;
signal \U400_SDRAM.N_216\ : std_logic;
signal \U400_SDRAM.N_187\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_2_0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_0C_net\ : std_logic;
signal \U400_SDRAM.TACK_7_iv_i_i_2\ : std_logic;
signal \U400_SDRAM.TACK_7_iv_i_i_1_0_cascade_\ : std_logic;
signal \U400_SDRAM.N_258\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_0_1\ : std_logic;
signal \U400_SDRAM.N_258_cascade_\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_0_0\ : std_logic;
signal \U400_SDRAM.N_240_cascade_\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \INVU400_SDRAM.REFRESH_COUNTER_1C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2\ : std_logic;
signal \U400_SDRAM.CS0_EN_0_cascade_\ : std_logic;
signal \U400_SDRAM.CS0_ENZ0\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U400_SDRAM.CS1_EN_0_cascade_\ : std_logic;
signal \INVU400_SDRAM.CS0_ENC_net\ : std_logic;
signal \U400_SDRAM.N_114_cascade_\ : std_logic;
signal \U400_SDRAM.N_220\ : std_logic;
signal \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3Z0Z_0\ : std_logic;
signal \U400_SDRAM.N_230_cascade_\ : std_logic;
signal \A_c_19\ : std_logic;
signal \MA_c_9\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_9C_net\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_29\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0\ : std_logic;
signal \A_c_21\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \A_c_22\ : std_logic;
signal \U400_SDRAM.N_240\ : std_logic;
signal \BANK1_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U400_SDRAM.N_82\ : std_logic;
signal \U400_SDRAM.N_34\ : std_logic;
signal \INVU400_SDRAM.BANK0C_net\ : std_logic;
signal \U400_SDRAM.N_118_cascade_\ : std_logic;
signal \U400_SDRAM.N_215\ : std_logic;
signal \U400_SDRAM.RAM_CYCLEZ0\ : std_logic;
signal \U400_SDRAM.N_236_cascade_\ : std_logic;
signal \U400_SDRAM.N_23_i\ : std_logic;
signal \U400_SDRAM.N_23_i_cascade_\ : std_logic;
signal \U400_SDRAM.N_242\ : std_logic;
signal \U400_SDRAM.N_139\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_1\ : std_logic;
signal \U400_SDRAM.N_198\ : std_logic;
signal \U400_SDRAM.N_259\ : std_logic;
signal \U400_SDRAM.N_118\ : std_logic;
signal \U400_SDRAM.N_39\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_3\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_1C_net\ : std_logic;
signal \U400_SDRAM.N_219_i\ : std_logic;
signal \U400_SDRAM.N_239\ : std_logic;
signal \U400_SDRAM.N_207\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_5_1_cascade_\ : std_logic;
signal \U400_SDRAM.N_250\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_31_i_i_i_2_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_31_i_i_i_3_cascade_\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_1C_net\ : std_logic;
signal \U400_SDRAM.N_261\ : std_logic;
signal \U400_SDRAM.N_140\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_4_1\ : std_logic;
signal \U400_SDRAM.CS1_ENZ0\ : std_logic;
signal \CS1n_c\ : std_logic;
signal \INVU400_SDRAM.CS1nC_net\ : std_logic;
signal \A_c_26\ : std_logic;
signal \MA_c_12\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_12C_net\ : std_logic;
signal \TA_OUT\ : std_logic;
signal \N_66\ : std_logic;
signal \U400_SDRAM.BURSTZ0\ : std_logic;
signal \U400_SDRAM.TA_EN11_m\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER26_0_cascade_\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER26_2_0\ : std_logic;
signal \U400_SDRAM.TA_COUNTER27\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_3\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.CO1\ : std_logic;
signal \U400_SDRAM.TA_COUNTER23\ : std_logic;
signal \U400_SDRAM.TACKZ0\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_0_sqmuxa\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_0\ : std_logic;
signal \CLK40_c_g\ : std_logic;
signal \U400_SDRAM.N_189\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U400_SDRAM.un1_REFRESH_COUNTERlto7_5\ : std_logic;
signal \U400_SDRAM.un1_REFRESH_COUNTERlto7_4\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_8\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER52_2_0_i_1\ : std_logic;
signal \U400_SDRAM.N_195_cascade_\ : std_logic;
signal \U400_SDRAM.N_94\ : std_logic;
signal \U400_ADDRESS_DECODE_RAM_SPACE_i_o3_0_o2_1\ : std_logic;
signal \A_c_31\ : std_logic;
signal \U400_ADDRESS_DECODE_RAM_SPACE_i_o3_0_o2_2\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U400_SDRAM.N_225\ : std_logic;
signal \U400_SDRAM.N_236\ : std_logic;
signal \U400_SDRAM.RAM_CYCLE_STARTZ0\ : std_logic;
signal \U400_SDRAM.N_228\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_a2_2_0_1_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_1_1_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_2_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.WRITE_CYCLEZ0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.N_256\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_a2_0_1_0_cascade_\ : std_logic;
signal \U400_SDRAM.N_97\ : std_logic;
signal \U400_SDRAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_0_0\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_1_0_cascade_\ : std_logic;
signal \U400_SDRAM.N_114\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_ne_0C_net\ : std_logic;
signal \U400_SDRAM.N_71\ : std_logic;
signal \A_c_25\ : std_logic;
signal \MA_c_11\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_11C_net\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U400_SDRAM.MA_5_iv_0_5\ : std_logic;
signal \MA_c_5\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_5C_net\ : std_logic;
signal \U400_BYTE_ENABLE.N_101_i\ : std_logic;
signal \U400_BYTE_ENABLE.N_101_i_cascade_\ : std_logic;
signal \un1_LMBEn_i_0_0\ : std_logic;
signal \A_c_0\ : std_logic;
signal \RAM_SPACE_i_o3_0_o2dup\ : std_logic;
signal \A_c_20\ : std_logic;
signal \MA_c_10\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_10C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \N_63\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \U400_BYTE_ENABLE.N_168\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \un1_LLBEn_i_0_0\ : std_logic;
signal \TA_EN_i_ess\ : std_logic;
signal \N_526_i\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_13\ : std_logic;
signal \MA_c_3\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_3C_net\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_12\ : std_logic;
signal \MA_c_2\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_10\ : std_logic;
signal \MA_c_0\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \MA_c_4\ : std_logic;
signal \U400_SDRAM.MA_5_iv_0_1\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U400_SDRAM.MA19\ : std_logic;
signal \MA_c_1\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_2C_net\ : std_logic;
signal \U400_SDRAM.un1_MA20_0_i_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \MA_wire\ : std_logic_vector(12 downto 0);
signal \A_wire\ : std_logic_vector(31 downto 0);
signal \CASn_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \UUBEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \LLBEn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \TAn_wire\ : std_logic;
signal \LBENn_wire\ : std_logic;
signal \CS1n_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CS0n_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CLK40_wire\ : std_logic;

begin
    MA <= \MA_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    BANK1 <= \BANK1_wire\;
    UUBEn <= \UUBEn_wire\;
    \SIZ_wire\ <= SIZ;
    LLBEn <= \LLBEn_wire\;
    \TSn_wire\ <= TSn;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    TAn <= \TAn_wire\;
    LBENn <= \LBENn_wire\;
    CS1n <= \CS1n_wire\;
    WEn <= \WEn_wire\;
    \RnW_wire\ <= RnW;
    CS0n <= \CS0n_wire\;
    LMBEn <= \LMBEn_wire\;
    \CLK40_wire\ <= CLK40;

    \MA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7125\,
            DIN => \N__7124\,
            DOUT => \N__7123\,
            PACKAGEPIN => \MA_wire\(7)
        );

    \MA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7125\,
            PADOUT => \N__7124\,
            PADIN => \N__7123\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2774\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7116\,
            DIN => \N__7115\,
            DOUT => \N__7114\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7116\,
            PADOUT => \N__7115\,
            PADIN => \N__7114\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7107\,
            DIN => \N__7106\,
            DOUT => \N__7105\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7107\,
            PADOUT => \N__7106\,
            PADIN => \N__7105\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2870\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7098\,
            DIN => \N__7097\,
            DOUT => \N__7096\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7098\,
            PADOUT => \N__7097\,
            PADIN => \N__7096\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3329\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7089\,
            DIN => \N__7088\,
            DOUT => \N__7087\,
            PACKAGEPIN => \MA_wire\(8)
        );

    \MA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7089\,
            PADOUT => \N__7088\,
            PADIN => \N__7087\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2810\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7080\,
            DIN => \N__7079\,
            DOUT => \N__7078\,
            PACKAGEPIN => \MA_wire\(10)
        );

    \MA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7080\,
            PADOUT => \N__7079\,
            PADIN => \N__7078\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6086\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7071\,
            DIN => \N__7070\,
            DOUT => \N__7069\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7071\,
            PADOUT => \N__7070\,
            PADIN => \N__7069\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7062\,
            DIN => \N__7061\,
            DOUT => \N__7060\,
            PACKAGEPIN => \MA_wire\(2)
        );

    \MA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7062\,
            PADOUT => \N__7061\,
            PADIN => \N__7060\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5597\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7053\,
            DIN => \N__7052\,
            DOUT => \N__7051\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7053\,
            PADOUT => \N__7052\,
            PADIN => \N__7051\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7044\,
            DIN => \N__7043\,
            DOUT => \N__7042\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7044\,
            PADOUT => \N__7043\,
            PADIN => \N__7042\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7035\,
            DIN => \N__7034\,
            DOUT => \N__7033\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7035\,
            PADOUT => \N__7034\,
            PADIN => \N__7033\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3752\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7026\,
            DIN => \N__7025\,
            DOUT => \N__7024\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7026\,
            PADOUT => \N__7025\,
            PADIN => \N__7024\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7017\,
            DIN => \N__7016\,
            DOUT => \N__7015\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7017\,
            PADOUT => \N__7016\,
            PADIN => \N__7015\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7008\,
            DIN => \N__7007\,
            DOUT => \N__7006\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7008\,
            PADOUT => \N__7007\,
            PADIN => \N__7006\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6999\,
            DIN => \N__6998\,
            DOUT => \N__6997\,
            PACKAGEPIN => \MA_wire\(12)
        );

    \MA_obuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6999\,
            PADOUT => \N__6998\,
            PADIN => \N__6997\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3584\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6990\,
            DIN => \N__6989\,
            DOUT => \N__6988\,
            PACKAGEPIN => \MA_wire\(1)
        );

    \MA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6990\,
            PADOUT => \N__6989\,
            PADIN => \N__6988\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6278\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6981\,
            DIN => \N__6980\,
            DOUT => \N__6979\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6981\,
            PADOUT => \N__6980\,
            PADIN => \N__6979\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6972\,
            DIN => \N__6971\,
            DOUT => \N__6970\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6972\,
            PADOUT => \N__6971\,
            PADIN => \N__6970\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6963\,
            DIN => \N__6962\,
            DOUT => \N__6961\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6963\,
            PADOUT => \N__6962\,
            PADIN => \N__6961\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6954\,
            DIN => \N__6953\,
            DOUT => \N__6952\,
            PACKAGEPIN => \MA_wire\(4)
        );

    \MA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6954\,
            PADOUT => \N__6953\,
            PADIN => \N__6952\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6368\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6945\,
            DIN => \N__6944\,
            DOUT => \N__6943\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6945\,
            PADOUT => \N__6944\,
            PADIN => \N__6943\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6936\,
            DIN => \N__6935\,
            DOUT => \N__6934\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6936\,
            PADOUT => \N__6935\,
            PADIN => \N__6934\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6927\,
            DIN => \N__6926\,
            DOUT => \N__6925\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6927\,
            PADOUT => \N__6926\,
            PADIN => \N__6925\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5696\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6918\,
            DIN => \N__6917\,
            DOUT => \N__6916\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6918\,
            PADOUT => \N__6917\,
            PADIN => \N__6916\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6909\,
            DIN => \N__6908\,
            DOUT => \N__6907\,
            PACKAGEPIN => \MA_wire\(9)
        );

    \MA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6909\,
            PADOUT => \N__6908\,
            PADIN => \N__6907\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3227\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6900\,
            DIN => \N__6899\,
            DOUT => \N__6898\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6900\,
            PADOUT => \N__6899\,
            PADIN => \N__6898\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5876\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6891\,
            DIN => \N__6890\,
            DOUT => \N__6889\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6891\,
            PADOUT => \N__6890\,
            PADIN => \N__6889\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6882\,
            DIN => \N__6881\,
            DOUT => \N__6880\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6882\,
            PADOUT => \N__6881\,
            PADIN => \N__6880\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6873\,
            DIN => \N__6872\,
            DOUT => \N__6871\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6873\,
            PADOUT => \N__6872\,
            PADIN => \N__6871\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2636\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6864\,
            DIN => \N__6863\,
            DOUT => \N__6862\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6864\,
            PADOUT => \N__6863\,
            PADIN => \N__6862\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6855\,
            DIN => \N__6854\,
            DOUT => \N__6853\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6855\,
            PADOUT => \N__6854\,
            PADIN => \N__6853\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6846\,
            DIN => \N__6845\,
            DOUT => \N__6844\,
            PACKAGEPIN => \MA_wire\(3)
        );

    \MA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6846\,
            PADOUT => \N__6845\,
            PADIN => \N__6844\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5639\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6837\,
            DIN => \N__6836\,
            DOUT => \N__6835\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6837\,
            PADOUT => \N__6836\,
            PADIN => \N__6835\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6828\,
            DIN => \N__6827\,
            DOUT => \N__6826\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6828\,
            PADOUT => \N__6827\,
            PADIN => \N__6826\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6819\,
            DIN => \N__6818\,
            DOUT => \N__6817\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6819\,
            PADOUT => \N__6818\,
            PADIN => \N__6817\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6810\,
            DIN => \N__6809\,
            DOUT => \N__6808\,
            PACKAGEPIN => \MA_wire\(6)
        );

    \MA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6810\,
            PADOUT => \N__6809\,
            PADIN => \N__6808\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2939\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6801\,
            DIN => \N__6800\,
            DOUT => \N__6799\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6801\,
            PADOUT => \N__6800\,
            PADIN => \N__6799\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6792\,
            DIN => \N__6791\,
            DOUT => \N__6790\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6792\,
            PADOUT => \N__6791\,
            PADIN => \N__6790\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6783\,
            DIN => \N__6782\,
            DOUT => \N__6781\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6783\,
            PADOUT => \N__6782\,
            PADIN => \N__6781\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6774\,
            DIN => \N__6773\,
            DOUT => \N__6772\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6774\,
            PADOUT => \N__6773\,
            PADIN => \N__6772\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2852\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6765\,
            DIN => \N__6764\,
            DOUT => \N__6763\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6765\,
            PADOUT => \N__6764\,
            PADIN => \N__6763\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6756\,
            DIN => \N__6755\,
            DOUT => \N__6754\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6756\,
            PADOUT => \N__6755\,
            PADIN => \N__6754\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3380\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6747\,
            DIN => \N__6746\,
            DOUT => \N__6745\,
            PACKAGEPIN => \MA_wire\(11)
        );

    \MA_obuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6747\,
            PADOUT => \N__6746\,
            PADIN => \N__6745\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5321\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6738\,
            DIN => \N__6737\,
            DOUT => \N__6736\,
            PACKAGEPIN => \TAn_wire\
        );

    \TAn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6738\,
            PADOUT => \N__6737\,
            PADIN => \N__6736\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5672\,
            DIN0 => OPEN,
            DOUT0 => \N__3773\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6729\,
            DIN => \N__6728\,
            DOUT => \N__6727\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6729\,
            PADOUT => \N__6728\,
            PADIN => \N__6727\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6720\,
            DIN => \N__6719\,
            DOUT => \N__6718\,
            PACKAGEPIN => \MA_wire\(5)
        );

    \MA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6720\,
            PADOUT => \N__6719\,
            PADIN => \N__6718\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5282\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6711\,
            DIN => \N__6710\,
            DOUT => \N__6709\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6711\,
            PADOUT => \N__6710\,
            PADIN => \N__6709\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6702\,
            DIN => \N__6701\,
            DOUT => \N__6700\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6702\,
            PADOUT => \N__6701\,
            PADIN => \N__6700\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LBENn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6693\,
            DIN => \N__6692\,
            DOUT => \N__6691\,
            PACKAGEPIN => \LBENn_wire\
        );

    \LBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6693\,
            PADOUT => \N__6692\,
            PADIN => \N__6691\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5194\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6684\,
            DIN => \N__6683\,
            DOUT => \N__6682\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6684\,
            PADOUT => \N__6683\,
            PADIN => \N__6682\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6675\,
            DIN => \N__6674\,
            DOUT => \N__6673\,
            PACKAGEPIN => \CS1n_wire\
        );

    \CS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6675\,
            PADOUT => \N__6674\,
            PADIN => \N__6673\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3614\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6666\,
            DIN => \N__6665\,
            DOUT => \N__6664\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6666\,
            PADOUT => \N__6665\,
            PADIN => \N__6664\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6657\,
            DIN => \N__6656\,
            DOUT => \N__6655\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6657\,
            PADOUT => \N__6656\,
            PADIN => \N__6655\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6648\,
            DIN => \N__6647\,
            DOUT => \N__6646\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6648\,
            PADOUT => \N__6647\,
            PADIN => \N__6646\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6639\,
            DIN => \N__6638\,
            DOUT => \N__6637\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6639\,
            PADOUT => \N__6638\,
            PADIN => \N__6637\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6630\,
            DIN => \N__6629\,
            DOUT => \N__6628\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6630\,
            PADOUT => \N__6629\,
            PADIN => \N__6628\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2861\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6621\,
            DIN => \N__6620\,
            DOUT => \N__6619\,
            PACKAGEPIN => \MA_wire\(0)
        );

    \MA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6621\,
            PADOUT => \N__6620\,
            PADIN => \N__6619\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5564\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6612\,
            DIN => \N__6611\,
            DOUT => \N__6610\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6612\,
            PADOUT => \N__6611\,
            PADIN => \N__6610\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6603\,
            DIN => \N__6602\,
            DOUT => \N__6601\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6603\,
            PADOUT => \N__6602\,
            PADIN => \N__6601\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6594\,
            DIN => \N__6593\,
            DOUT => \N__6592\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6594\,
            PADOUT => \N__6593\,
            PADIN => \N__6592\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6585\,
            DIN => \N__6584\,
            DOUT => \N__6583\,
            PACKAGEPIN => \CS0n_wire\
        );

    \CS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6585\,
            PADOUT => \N__6584\,
            PADIN => \N__6583\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2882\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6576\,
            DIN => \N__6575\,
            DOUT => \N__6574\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6576\,
            PADOUT => \N__6575\,
            PADIN => \N__6574\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6567\,
            DIN => \N__6566\,
            DOUT => \N__6565\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6567\,
            PADOUT => \N__6566\,
            PADIN => \N__6565\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5258\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6558\,
            DIN => \N__6557\,
            DOUT => \N__6556\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6558\,
            PADOUT => \N__6557\,
            PADIN => \N__6556\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6549\,
            DIN => \N__6548\,
            DOUT => \N__6547\,
            PACKAGEPIN => \CLK40_wire\
        );

    \CLK40_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6549\,
            PADOUT => \N__6548\,
            PADIN => \N__6547\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_ibuf_gb_io_gb_input\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1554\ : InMux
    port map (
            O => \N__6530\,
            I => \N__6527\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__6527\,
            I => \N__6524\
        );

    \I__1552\ : Span4Mux_s3_v
    port map (
            O => \N__6524\,
            I => \N__6521\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__6521\,
            I => \A_c_6\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__6518\,
            I => \N__6515\
        );

    \I__1549\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6512\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__6512\,
            I => \N__6509\
        );

    \I__1547\ : IoSpan4Mux
    port map (
            O => \N__6509\,
            I => \N__6506\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__6506\,
            I => \A_c_14\
        );

    \I__1545\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6492\
        );

    \I__1544\ : InMux
    port map (
            O => \N__6502\,
            I => \N__6486\
        );

    \I__1543\ : InMux
    port map (
            O => \N__6501\,
            I => \N__6482\
        );

    \I__1542\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6479\
        );

    \I__1541\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6476\
        );

    \I__1540\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6469\
        );

    \I__1539\ : InMux
    port map (
            O => \N__6497\,
            I => \N__6469\
        );

    \I__1538\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6466\
        );

    \I__1537\ : InMux
    port map (
            O => \N__6495\,
            I => \N__6463\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__6492\,
            I => \N__6459\
        );

    \I__1535\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6454\
        );

    \I__1534\ : InMux
    port map (
            O => \N__6490\,
            I => \N__6454\
        );

    \I__1533\ : InMux
    port map (
            O => \N__6489\,
            I => \N__6451\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__6486\,
            I => \N__6447\
        );

    \I__1531\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6444\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__6482\,
            I => \N__6437\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__6479\,
            I => \N__6437\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__6476\,
            I => \N__6437\
        );

    \I__1527\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6432\
        );

    \I__1526\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6432\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__6469\,
            I => \N__6427\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__6466\,
            I => \N__6427\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__6463\,
            I => \N__6422\
        );

    \I__1522\ : InMux
    port map (
            O => \N__6462\,
            I => \N__6419\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__6459\,
            I => \N__6412\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__6454\,
            I => \N__6412\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__6451\,
            I => \N__6412\
        );

    \I__1518\ : InMux
    port map (
            O => \N__6450\,
            I => \N__6409\
        );

    \I__1517\ : Span4Mux_h
    port map (
            O => \N__6447\,
            I => \N__6400\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__6444\,
            I => \N__6400\
        );

    \I__1515\ : Span4Mux_v
    port map (
            O => \N__6437\,
            I => \N__6400\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__6432\,
            I => \N__6400\
        );

    \I__1513\ : Span12Mux_s8_v
    port map (
            O => \N__6427\,
            I => \N__6397\
        );

    \I__1512\ : InMux
    port map (
            O => \N__6426\,
            I => \N__6394\
        );

    \I__1511\ : InMux
    port map (
            O => \N__6425\,
            I => \N__6391\
        );

    \I__1510\ : Span12Mux_s6_h
    port map (
            O => \N__6422\,
            I => \N__6386\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__6419\,
            I => \N__6386\
        );

    \I__1508\ : Span4Mux_v
    port map (
            O => \N__6412\,
            I => \N__6379\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__6409\,
            I => \N__6379\
        );

    \I__1506\ : Span4Mux_v
    port map (
            O => \N__6400\,
            I => \N__6379\
        );

    \I__1505\ : Odrv12
    port map (
            O => \N__6397\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__6394\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__6391\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1502\ : Odrv12
    port map (
            O => \N__6386\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__6379\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1500\ : IoInMux
    port map (
            O => \N__6368\,
            I => \N__6365\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__6365\,
            I => \N__6362\
        );

    \I__1498\ : Span4Mux_s1_v
    port map (
            O => \N__6362\,
            I => \N__6359\
        );

    \I__1497\ : Span4Mux_h
    port map (
            O => \N__6359\,
            I => \N__6356\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__6356\,
            I => \MA_c_4\
        );

    \I__1495\ : InMux
    port map (
            O => \N__6353\,
            I => \N__6350\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__6350\,
            I => \U400_SDRAM.MA_5_iv_0_1\
        );

    \I__1493\ : InMux
    port map (
            O => \N__6347\,
            I => \N__6344\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__6344\,
            I => \N__6341\
        );

    \I__1491\ : Odrv4
    port map (
            O => \N__6341\,
            I => \A_c_11\
        );

    \I__1490\ : InMux
    port map (
            O => \N__6338\,
            I => \N__6328\
        );

    \I__1489\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6325\
        );

    \I__1488\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6316\
        );

    \I__1487\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6316\
        );

    \I__1486\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6316\
        );

    \I__1485\ : InMux
    port map (
            O => \N__6333\,
            I => \N__6316\
        );

    \I__1484\ : InMux
    port map (
            O => \N__6332\,
            I => \N__6311\
        );

    \I__1483\ : InMux
    port map (
            O => \N__6331\,
            I => \N__6311\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__6328\,
            I => \N__6307\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__6325\,
            I => \N__6304\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__6316\,
            I => \N__6301\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__6311\,
            I => \N__6298\
        );

    \I__1478\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6295\
        );

    \I__1477\ : Span4Mux_h
    port map (
            O => \N__6307\,
            I => \N__6290\
        );

    \I__1476\ : Span4Mux_s2_v
    port map (
            O => \N__6304\,
            I => \N__6290\
        );

    \I__1475\ : Span4Mux_s2_v
    port map (
            O => \N__6301\,
            I => \N__6287\
        );

    \I__1474\ : Odrv12
    port map (
            O => \N__6298\,
            I => \U400_SDRAM.MA19\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__6295\,
            I => \U400_SDRAM.MA19\
        );

    \I__1472\ : Odrv4
    port map (
            O => \N__6290\,
            I => \U400_SDRAM.MA19\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__6287\,
            I => \U400_SDRAM.MA19\
        );

    \I__1470\ : IoInMux
    port map (
            O => \N__6278\,
            I => \N__6275\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__6275\,
            I => \N__6272\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__6272\,
            I => \MA_c_1\
        );

    \I__1467\ : CEMux
    port map (
            O => \N__6269\,
            I => \N__6262\
        );

    \I__1466\ : CEMux
    port map (
            O => \N__6268\,
            I => \N__6259\
        );

    \I__1465\ : CEMux
    port map (
            O => \N__6267\,
            I => \N__6255\
        );

    \I__1464\ : CEMux
    port map (
            O => \N__6266\,
            I => \N__6251\
        );

    \I__1463\ : CEMux
    port map (
            O => \N__6265\,
            I => \N__6248\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__6262\,
            I => \N__6245\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__6259\,
            I => \N__6242\
        );

    \I__1460\ : CEMux
    port map (
            O => \N__6258\,
            I => \N__6238\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__6255\,
            I => \N__6234\
        );

    \I__1458\ : CEMux
    port map (
            O => \N__6254\,
            I => \N__6231\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__6251\,
            I => \N__6228\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__6248\,
            I => \N__6225\
        );

    \I__1455\ : Span4Mux_v
    port map (
            O => \N__6245\,
            I => \N__6220\
        );

    \I__1454\ : Span4Mux_h
    port map (
            O => \N__6242\,
            I => \N__6220\
        );

    \I__1453\ : CEMux
    port map (
            O => \N__6241\,
            I => \N__6217\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__6238\,
            I => \N__6214\
        );

    \I__1451\ : CEMux
    port map (
            O => \N__6237\,
            I => \N__6211\
        );

    \I__1450\ : Span4Mux_h
    port map (
            O => \N__6234\,
            I => \N__6206\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__6231\,
            I => \N__6206\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__6228\,
            I => \U400_SDRAM.un1_MA20_0_i_0\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__6225\,
            I => \U400_SDRAM.un1_MA20_0_i_0\
        );

    \I__1446\ : Odrv4
    port map (
            O => \N__6220\,
            I => \U400_SDRAM.un1_MA20_0_i_0\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__6217\,
            I => \U400_SDRAM.un1_MA20_0_i_0\
        );

    \I__1444\ : Odrv12
    port map (
            O => \N__6214\,
            I => \U400_SDRAM.un1_MA20_0_i_0\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__6211\,
            I => \U400_SDRAM.un1_MA20_0_i_0\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__6206\,
            I => \U400_SDRAM.un1_MA20_0_i_0\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__6191\,
            I => \N__6188\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6184\
        );

    \I__1439\ : InMux
    port map (
            O => \N__6187\,
            I => \N__6181\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__6184\,
            I => \N__6174\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__6181\,
            I => \N__6166\
        );

    \I__1436\ : SRMux
    port map (
            O => \N__6180\,
            I => \N__6116\
        );

    \I__1435\ : SRMux
    port map (
            O => \N__6179\,
            I => \N__6116\
        );

    \I__1434\ : SRMux
    port map (
            O => \N__6178\,
            I => \N__6116\
        );

    \I__1433\ : SRMux
    port map (
            O => \N__6177\,
            I => \N__6116\
        );

    \I__1432\ : Glb2LocalMux
    port map (
            O => \N__6174\,
            I => \N__6116\
        );

    \I__1431\ : SRMux
    port map (
            O => \N__6173\,
            I => \N__6116\
        );

    \I__1430\ : SRMux
    port map (
            O => \N__6172\,
            I => \N__6116\
        );

    \I__1429\ : SRMux
    port map (
            O => \N__6171\,
            I => \N__6116\
        );

    \I__1428\ : SRMux
    port map (
            O => \N__6170\,
            I => \N__6116\
        );

    \I__1427\ : SRMux
    port map (
            O => \N__6169\,
            I => \N__6116\
        );

    \I__1426\ : Glb2LocalMux
    port map (
            O => \N__6166\,
            I => \N__6116\
        );

    \I__1425\ : SRMux
    port map (
            O => \N__6165\,
            I => \N__6116\
        );

    \I__1424\ : SRMux
    port map (
            O => \N__6164\,
            I => \N__6116\
        );

    \I__1423\ : SRMux
    port map (
            O => \N__6163\,
            I => \N__6116\
        );

    \I__1422\ : SRMux
    port map (
            O => \N__6162\,
            I => \N__6116\
        );

    \I__1421\ : SRMux
    port map (
            O => \N__6161\,
            I => \N__6116\
        );

    \I__1420\ : SRMux
    port map (
            O => \N__6160\,
            I => \N__6116\
        );

    \I__1419\ : SRMux
    port map (
            O => \N__6159\,
            I => \N__6116\
        );

    \I__1418\ : SRMux
    port map (
            O => \N__6158\,
            I => \N__6116\
        );

    \I__1417\ : SRMux
    port map (
            O => \N__6157\,
            I => \N__6116\
        );

    \I__1416\ : GlobalMux
    port map (
            O => \N__6116\,
            I => \N__6113\
        );

    \I__1415\ : gio2CtrlBuf
    port map (
            O => \N__6113\,
            I => \RESETn_c_i_g\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__6110\,
            I => \N__6107\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6107\,
            I => \N__6104\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6104\,
            I => \N__6101\
        );

    \I__1411\ : Span4Mux_v
    port map (
            O => \N__6101\,
            I => \N__6098\
        );

    \I__1410\ : Span4Mux_v
    port map (
            O => \N__6098\,
            I => \N__6095\
        );

    \I__1409\ : Span4Mux_v
    port map (
            O => \N__6095\,
            I => \N__6092\
        );

    \I__1408\ : Sp12to4
    port map (
            O => \N__6092\,
            I => \N__6089\
        );

    \I__1407\ : Odrv12
    port map (
            O => \N__6089\,
            I => \A_c_20\
        );

    \I__1406\ : IoInMux
    port map (
            O => \N__6086\,
            I => \N__6083\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__6083\,
            I => \N__6080\
        );

    \I__1404\ : Odrv12
    port map (
            O => \N__6080\,
            I => \MA_c_10\
        );

    \I__1403\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6071\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6064\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6075\,
            I => \N__6059\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6074\,
            I => \N__6056\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6071\,
            I => \N__6053\
        );

    \I__1398\ : InMux
    port map (
            O => \N__6070\,
            I => \N__6050\
        );

    \I__1397\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6047\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6068\,
            I => \N__6044\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6041\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6064\,
            I => \N__6037\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6063\,
            I => \N__6032\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6062\,
            I => \N__6032\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6059\,
            I => \N__6022\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6056\,
            I => \N__6022\
        );

    \I__1389\ : Span4Mux_h
    port map (
            O => \N__6053\,
            I => \N__6022\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6050\,
            I => \N__6022\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__6047\,
            I => \N__6017\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__6044\,
            I => \N__6017\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__6041\,
            I => \N__6014\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6040\,
            I => \N__6011\
        );

    \I__1383\ : Span4Mux_v
    port map (
            O => \N__6037\,
            I => \N__6006\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__6032\,
            I => \N__6006\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6031\,
            I => \N__6003\
        );

    \I__1380\ : Span4Mux_v
    port map (
            O => \N__6022\,
            I => \N__6000\
        );

    \I__1379\ : Span4Mux_v
    port map (
            O => \N__6017\,
            I => \N__5991\
        );

    \I__1378\ : Span4Mux_h
    port map (
            O => \N__6014\,
            I => \N__5991\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__6011\,
            I => \N__5991\
        );

    \I__1376\ : Span4Mux_v
    port map (
            O => \N__6006\,
            I => \N__5991\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__6003\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__6000\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__5991\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__5984\,
            I => \N__5981\
        );

    \I__1371\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5978\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__5978\,
            I => \N__5975\
        );

    \I__1369\ : Span4Mux_h
    port map (
            O => \N__5975\,
            I => \N__5972\
        );

    \I__1368\ : Odrv4
    port map (
            O => \N__5972\,
            I => \A_c_3\
        );

    \I__1367\ : CascadeMux
    port map (
            O => \N__5969\,
            I => \N__5964\
        );

    \I__1366\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5961\
        );

    \I__1365\ : InMux
    port map (
            O => \N__5967\,
            I => \N__5951\
        );

    \I__1364\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5948\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__5961\,
            I => \N__5945\
        );

    \I__1362\ : InMux
    port map (
            O => \N__5960\,
            I => \N__5942\
        );

    \I__1361\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5939\
        );

    \I__1360\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5936\
        );

    \I__1359\ : InMux
    port map (
            O => \N__5957\,
            I => \N__5933\
        );

    \I__1358\ : InMux
    port map (
            O => \N__5956\,
            I => \N__5930\
        );

    \I__1357\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5925\
        );

    \I__1356\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5925\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__5951\,
            I => \N__5921\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__5948\,
            I => \N__5918\
        );

    \I__1353\ : Span4Mux_h
    port map (
            O => \N__5945\,
            I => \N__5913\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__5942\,
            I => \N__5913\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__5939\,
            I => \N__5906\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__5936\,
            I => \N__5906\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__5933\,
            I => \N__5906\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__5930\,
            I => \N__5901\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__5925\,
            I => \N__5901\
        );

    \I__1346\ : InMux
    port map (
            O => \N__5924\,
            I => \N__5898\
        );

    \I__1345\ : Span4Mux_h
    port map (
            O => \N__5921\,
            I => \N__5895\
        );

    \I__1344\ : Span4Mux_h
    port map (
            O => \N__5918\,
            I => \N__5890\
        );

    \I__1343\ : Span4Mux_v
    port map (
            O => \N__5913\,
            I => \N__5890\
        );

    \I__1342\ : Span4Mux_v
    port map (
            O => \N__5906\,
            I => \N__5885\
        );

    \I__1341\ : Span4Mux_v
    port map (
            O => \N__5901\,
            I => \N__5885\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__5898\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1339\ : Odrv4
    port map (
            O => \N__5895\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__5890\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1337\ : Odrv4
    port map (
            O => \N__5885\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1336\ : IoInMux
    port map (
            O => \N__5876\,
            I => \N__5873\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__5873\,
            I => \N__5870\
        );

    \I__1334\ : Odrv4
    port map (
            O => \N__5870\,
            I => \N_63\
        );

    \I__1333\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5861\
        );

    \I__1332\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5861\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__5861\,
            I => \N__5858\
        );

    \I__1330\ : Span4Mux_v
    port map (
            O => \N__5858\,
            I => \N__5854\
        );

    \I__1329\ : InMux
    port map (
            O => \N__5857\,
            I => \N__5850\
        );

    \I__1328\ : Span4Mux_v
    port map (
            O => \N__5854\,
            I => \N__5847\
        );

    \I__1327\ : InMux
    port map (
            O => \N__5853\,
            I => \N__5844\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__5850\,
            I => \N__5841\
        );

    \I__1325\ : Span4Mux_v
    port map (
            O => \N__5847\,
            I => \N__5838\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__5844\,
            I => \N__5833\
        );

    \I__1323\ : Sp12to4
    port map (
            O => \N__5841\,
            I => \N__5833\
        );

    \I__1322\ : Sp12to4
    port map (
            O => \N__5838\,
            I => \N__5828\
        );

    \I__1321\ : Span12Mux_v
    port map (
            O => \N__5833\,
            I => \N__5828\
        );

    \I__1320\ : Odrv12
    port map (
            O => \N__5828\,
            I => \A_c_1\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__5825\,
            I => \N__5819\
        );

    \I__1318\ : InMux
    port map (
            O => \N__5824\,
            I => \N__5816\
        );

    \I__1317\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5813\
        );

    \I__1316\ : InMux
    port map (
            O => \N__5822\,
            I => \N__5808\
        );

    \I__1315\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5805\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__5816\,
            I => \N__5800\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5813\,
            I => \N__5800\
        );

    \I__1312\ : InMux
    port map (
            O => \N__5812\,
            I => \N__5795\
        );

    \I__1311\ : InMux
    port map (
            O => \N__5811\,
            I => \N__5795\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__5808\,
            I => \N__5790\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__5805\,
            I => \N__5790\
        );

    \I__1308\ : Span4Mux_v
    port map (
            O => \N__5800\,
            I => \N__5787\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__5795\,
            I => \N__5784\
        );

    \I__1306\ : Span4Mux_v
    port map (
            O => \N__5790\,
            I => \N__5781\
        );

    \I__1305\ : Span4Mux_h
    port map (
            O => \N__5787\,
            I => \N__5776\
        );

    \I__1304\ : Span4Mux_v
    port map (
            O => \N__5784\,
            I => \N__5776\
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__5781\,
            I => \SIZ_c_1\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__5776\,
            I => \SIZ_c_1\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__5771\,
            I => \N__5767\
        );

    \I__1300\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5762\
        );

    \I__1299\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5762\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__5762\,
            I => \U400_BYTE_ENABLE.N_168\
        );

    \I__1297\ : InMux
    port map (
            O => \N__5759\,
            I => \N__5752\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__5758\,
            I => \N__5749\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5757\,
            I => \N__5745\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5742\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5739\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5752\,
            I => \N__5736\
        );

    \I__1291\ : InMux
    port map (
            O => \N__5749\,
            I => \N__5731\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5731\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5745\,
            I => \N__5728\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__5742\,
            I => \N__5725\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5739\,
            I => \N__5718\
        );

    \I__1286\ : Span4Mux_v
    port map (
            O => \N__5736\,
            I => \N__5718\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__5731\,
            I => \N__5718\
        );

    \I__1284\ : Span4Mux_v
    port map (
            O => \N__5728\,
            I => \N__5715\
        );

    \I__1283\ : Span4Mux_v
    port map (
            O => \N__5725\,
            I => \N__5712\
        );

    \I__1282\ : Span4Mux_h
    port map (
            O => \N__5718\,
            I => \N__5709\
        );

    \I__1281\ : Span4Mux_h
    port map (
            O => \N__5715\,
            I => \N__5704\
        );

    \I__1280\ : Span4Mux_h
    port map (
            O => \N__5712\,
            I => \N__5704\
        );

    \I__1279\ : Span4Mux_v
    port map (
            O => \N__5709\,
            I => \N__5701\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__5704\,
            I => \SIZ_c_0\
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__5701\,
            I => \SIZ_c_0\
        );

    \I__1276\ : IoInMux
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5693\,
            I => \N__5690\
        );

    \I__1274\ : Span4Mux_s2_v
    port map (
            O => \N__5690\,
            I => \N__5687\
        );

    \I__1273\ : Odrv4
    port map (
            O => \N__5687\,
            I => \un1_LLBEn_i_0_0\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5684\,
            I => \N__5681\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__5681\,
            I => \N__5678\
        );

    \I__1270\ : Span4Mux_v
    port map (
            O => \N__5678\,
            I => \N__5675\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__5675\,
            I => \TA_EN_i_ess\
        );

    \I__1268\ : IoInMux
    port map (
            O => \N__5672\,
            I => \N__5669\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__5669\,
            I => \N__5666\
        );

    \I__1266\ : Odrv4
    port map (
            O => \N__5666\,
            I => \N_526_i\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5660\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5660\,
            I => \N__5657\
        );

    \I__1263\ : Odrv4
    port map (
            O => \N__5657\,
            I => \A_c_5\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__5654\,
            I => \N__5651\
        );

    \I__1261\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5648\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5648\,
            I => \N__5645\
        );

    \I__1259\ : Span4Mux_v
    port map (
            O => \N__5645\,
            I => \N__5642\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__5642\,
            I => \A_c_13\
        );

    \I__1257\ : IoInMux
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__5636\,
            I => \N__5633\
        );

    \I__1255\ : IoSpan4Mux
    port map (
            O => \N__5633\,
            I => \N__5630\
        );

    \I__1254\ : Span4Mux_s3_h
    port map (
            O => \N__5630\,
            I => \N__5627\
        );

    \I__1253\ : Span4Mux_h
    port map (
            O => \N__5627\,
            I => \N__5624\
        );

    \I__1252\ : Odrv4
    port map (
            O => \N__5624\,
            I => \MA_c_3\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5621\,
            I => \N__5618\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5618\,
            I => \N__5615\
        );

    \I__1249\ : Span4Mux_v
    port map (
            O => \N__5615\,
            I => \N__5612\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__5612\,
            I => \A_c_4\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__5609\,
            I => \N__5606\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5606\,
            I => \N__5603\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__5603\,
            I => \N__5600\
        );

    \I__1244\ : Odrv4
    port map (
            O => \N__5600\,
            I => \A_c_12\
        );

    \I__1243\ : IoInMux
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5594\,
            I => \N__5591\
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__5591\,
            I => \MA_c_2\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5588\,
            I => \N__5585\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__5585\,
            I => \N__5582\
        );

    \I__1238\ : Span4Mux_h
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__5579\,
            I => \A_c_2\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5573\,
            I => \N__5570\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5570\,
            I => \N__5567\
        );

    \I__1233\ : Odrv4
    port map (
            O => \N__5567\,
            I => \A_c_10\
        );

    \I__1232\ : IoInMux
    port map (
            O => \N__5564\,
            I => \N__5561\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__1230\ : Span4Mux_s1_v
    port map (
            O => \N__5558\,
            I => \N__5555\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__5555\,
            I => \MA_c_0\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5552\,
            I => \N__5539\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5551\,
            I => \N__5539\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5550\,
            I => \N__5534\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5549\,
            I => \N__5534\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__5548\,
            I => \N__5530\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__5547\,
            I => \N__5524\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__5546\,
            I => \N__5517\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__5545\,
            I => \N__5513\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__5544\,
            I => \N__5510\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5539\,
            I => \N__5505\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5534\,
            I => \N__5505\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5500\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5530\,
            I => \N__5500\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5529\,
            I => \N__5497\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5528\,
            I => \N__5494\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5491\
        );

    \I__1212\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5484\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5484\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5484\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5477\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5477\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5477\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5516\,
            I => \N__5474\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5513\,
            I => \N__5471\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5468\
        );

    \I__1203\ : Span4Mux_h
    port map (
            O => \N__5505\,
            I => \N__5465\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5500\,
            I => \N__5458\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__5497\,
            I => \N__5458\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5494\,
            I => \N__5458\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5491\,
            I => \N__5449\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5484\,
            I => \N__5449\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5477\,
            I => \N__5449\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5474\,
            I => \N__5446\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5471\,
            I => \N__5441\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5468\,
            I => \N__5441\
        );

    \I__1193\ : Span4Mux_v
    port map (
            O => \N__5465\,
            I => \N__5436\
        );

    \I__1192\ : Span4Mux_v
    port map (
            O => \N__5458\,
            I => \N__5436\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5457\,
            I => \N__5431\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5431\
        );

    \I__1189\ : Span4Mux_v
    port map (
            O => \N__5449\,
            I => \N__5428\
        );

    \I__1188\ : Span4Mux_v
    port map (
            O => \N__5446\,
            I => \N__5423\
        );

    \I__1187\ : Span4Mux_h
    port map (
            O => \N__5441\,
            I => \N__5423\
        );

    \I__1186\ : Odrv4
    port map (
            O => \N__5436\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__5431\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1184\ : Odrv4
    port map (
            O => \N__5428\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1183\ : Odrv4
    port map (
            O => \N__5423\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5411\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_0_0\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__5408\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_1_0_cascade_\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5405\,
            I => \N__5402\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5402\,
            I => \N__5399\
        );

    \I__1177\ : Span4Mux_v
    port map (
            O => \N__5399\,
            I => \N__5388\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5398\,
            I => \N__5383\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5383\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5396\,
            I => \N__5380\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5377\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5370\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5370\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5392\,
            I => \N__5370\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5391\,
            I => \N__5367\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__5388\,
            I => \U400_SDRAM.N_114\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__5383\,
            I => \U400_SDRAM.N_114\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5380\,
            I => \U400_SDRAM.N_114\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5377\,
            I => \U400_SDRAM.N_114\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5370\,
            I => \U400_SDRAM.N_114\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5367\,
            I => \U400_SDRAM.N_114\
        );

    \I__1162\ : CEMux
    port map (
            O => \N__5354\,
            I => \N__5351\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5351\,
            I => \N__5346\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5341\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5341\
        );

    \I__1158\ : Odrv12
    port map (
            O => \N__5346\,
            I => \U400_SDRAM.N_71\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5341\,
            I => \U400_SDRAM.N_71\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__5336\,
            I => \N__5333\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5333\,
            I => \N__5330\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__1153\ : Span12Mux_s7_v
    port map (
            O => \N__5327\,
            I => \N__5324\
        );

    \I__1152\ : Odrv12
    port map (
            O => \N__5324\,
            I => \A_c_25\
        );

    \I__1151\ : IoInMux
    port map (
            O => \N__5321\,
            I => \N__5318\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5318\,
            I => \N__5315\
        );

    \I__1149\ : Odrv12
    port map (
            O => \N__5315\,
            I => \MA_c_11\
        );

    \I__1148\ : CascadeMux
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5306\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5306\,
            I => \N__5303\
        );

    \I__1145\ : Odrv12
    port map (
            O => \N__5303\,
            I => \A_c_7\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5297\,
            I => \N__5294\
        );

    \I__1142\ : IoSpan4Mux
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__5291\,
            I => \A_c_15\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5288\,
            I => \N__5285\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5285\,
            I => \U400_SDRAM.MA_5_iv_0_5\
        );

    \I__1138\ : IoInMux
    port map (
            O => \N__5282\,
            I => \N__5279\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5279\,
            I => \N__5276\
        );

    \I__1136\ : Span4Mux_s2_v
    port map (
            O => \N__5276\,
            I => \N__5273\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__5270\,
            I => \MA_c_5\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5264\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__5264\,
            I => \U400_BYTE_ENABLE.N_101_i\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__5261\,
            I => \U400_BYTE_ENABLE.N_101_i_cascade_\
        );

    \I__1130\ : IoInMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__5255\,
            I => \N__5252\
        );

    \I__1128\ : Span4Mux_s3_v
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__1127\ : Odrv4
    port map (
            O => \N__5249\,
            I => \un1_LMBEn_i_0_0\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5242\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5245\,
            I => \N__5239\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5242\,
            I => \N__5235\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__5239\,
            I => \N__5232\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5238\,
            I => \N__5229\
        );

    \I__1121\ : Span4Mux_v
    port map (
            O => \N__5235\,
            I => \N__5226\
        );

    \I__1120\ : Span4Mux_v
    port map (
            O => \N__5232\,
            I => \N__5223\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5229\,
            I => \N__5220\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__5226\,
            I => \N__5217\
        );

    \I__1117\ : Sp12to4
    port map (
            O => \N__5223\,
            I => \N__5214\
        );

    \I__1116\ : Span4Mux_h
    port map (
            O => \N__5220\,
            I => \N__5211\
        );

    \I__1115\ : Span4Mux_v
    port map (
            O => \N__5217\,
            I => \N__5208\
        );

    \I__1114\ : Span12Mux_s6_h
    port map (
            O => \N__5214\,
            I => \N__5203\
        );

    \I__1113\ : Sp12to4
    port map (
            O => \N__5211\,
            I => \N__5203\
        );

    \I__1112\ : Sp12to4
    port map (
            O => \N__5208\,
            I => \N__5198\
        );

    \I__1111\ : Span12Mux_v
    port map (
            O => \N__5203\,
            I => \N__5198\
        );

    \I__1110\ : Odrv12
    port map (
            O => \N__5198\,
            I => \A_c_0\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__5195\,
            I => \N__5190\
        );

    \I__1108\ : IoInMux
    port map (
            O => \N__5194\,
            I => \N__5187\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5184\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5190\,
            I => \N__5180\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5187\,
            I => \N__5177\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5184\,
            I => \N__5174\
        );

    \I__1103\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5171\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5180\,
            I => \N__5168\
        );

    \I__1101\ : Odrv12
    port map (
            O => \N__5177\,
            I => \RAM_SPACE_i_o3_0_o2dup\
        );

    \I__1100\ : Odrv4
    port map (
            O => \N__5174\,
            I => \RAM_SPACE_i_o3_0_o2dup\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5171\,
            I => \RAM_SPACE_i_o3_0_o2dup\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__5168\,
            I => \RAM_SPACE_i_o3_0_o2dup\
        );

    \I__1097\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5156\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5156\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER52_2_0_i_1\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__5153\,
            I => \U400_SDRAM.N_195_cascade_\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5147\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5147\,
            I => \U400_SDRAM.N_94\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__5144\,
            I => \N__5140\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5143\,
            I => \N__5137\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5140\,
            I => \N__5134\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5137\,
            I => \N__5131\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5134\,
            I => \N__5128\
        );

    \I__1087\ : Span4Mux_v
    port map (
            O => \N__5131\,
            I => \N__5123\
        );

    \I__1086\ : Span4Mux_v
    port map (
            O => \N__5128\,
            I => \N__5123\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__5123\,
            I => \U400_ADDRESS_DECODE_RAM_SPACE_i_o3_0_o2_1\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5117\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__5117\,
            I => \N__5113\
        );

    \I__1082\ : InMux
    port map (
            O => \N__5116\,
            I => \N__5110\
        );

    \I__1081\ : Span4Mux_h
    port map (
            O => \N__5113\,
            I => \N__5107\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__5110\,
            I => \N__5104\
        );

    \I__1079\ : Span4Mux_h
    port map (
            O => \N__5107\,
            I => \N__5101\
        );

    \I__1078\ : Span12Mux_s10_h
    port map (
            O => \N__5104\,
            I => \N__5098\
        );

    \I__1077\ : Span4Mux_v
    port map (
            O => \N__5101\,
            I => \N__5095\
        );

    \I__1076\ : Odrv12
    port map (
            O => \N__5098\,
            I => \A_c_31\
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__5095\,
            I => \A_c_31\
        );

    \I__1074\ : CascadeMux
    port map (
            O => \N__5090\,
            I => \N__5087\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5084\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5084\,
            I => \N__5080\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5083\,
            I => \N__5077\
        );

    \I__1070\ : Span4Mux_v
    port map (
            O => \N__5080\,
            I => \N__5072\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5077\,
            I => \N__5072\
        );

    \I__1068\ : Span4Mux_v
    port map (
            O => \N__5072\,
            I => \N__5069\
        );

    \I__1067\ : Sp12to4
    port map (
            O => \N__5069\,
            I => \N__5066\
        );

    \I__1066\ : Odrv12
    port map (
            O => \N__5066\,
            I => \U400_ADDRESS_DECODE_RAM_SPACE_i_o3_0_o2_2\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5060\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__5060\,
            I => \N__5057\
        );

    \I__1063\ : Odrv12
    port map (
            O => \N__5057\,
            I => \TSn_c\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5054\,
            I => \N__5051\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5051\,
            I => \U400_SDRAM.N_225\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__5048\,
            I => \N__5040\
        );

    \I__1059\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5036\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5046\,
            I => \N__5031\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5045\,
            I => \N__5031\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5028\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5025\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5022\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5019\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5036\,
            I => \N__5016\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5031\,
            I => \U400_SDRAM.N_236\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__5028\,
            I => \U400_SDRAM.N_236\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5025\,
            I => \U400_SDRAM.N_236\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5022\,
            I => \U400_SDRAM.N_236\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5019\,
            I => \U400_SDRAM.N_236\
        );

    \I__1046\ : Odrv4
    port map (
            O => \N__5016\,
            I => \U400_SDRAM.N_236\
        );

    \I__1045\ : InMux
    port map (
            O => \N__5003\,
            I => \N__4990\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5002\,
            I => \N__4990\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4987\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4984\
        );

    \I__1041\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4975\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4975\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4975\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4975\
        );

    \I__1037\ : InMux
    port map (
            O => \N__4995\,
            I => \N__4972\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4990\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__4987\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__4984\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__4975\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__4972\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__1031\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4958\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__4958\,
            I => \U400_SDRAM.N_228\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__4955\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_a2_2_0_1_cascade_\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__4952\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_1_1_cascade_\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__4949\,
            I => \N__4943\
        );

    \I__1026\ : InMux
    port map (
            O => \N__4948\,
            I => \N__4937\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4947\,
            I => \N__4932\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4946\,
            I => \N__4932\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4927\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4920\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4941\,
            I => \N__4920\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4940\,
            I => \N__4917\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__4937\,
            I => \N__4914\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4932\,
            I => \N__4911\
        );

    \I__1017\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4902\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4902\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__4927\,
            I => \N__4895\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4892\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4889\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__4920\,
            I => \N__4884\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4917\,
            I => \N__4884\
        );

    \I__1010\ : Span4Mux_h
    port map (
            O => \N__4914\,
            I => \N__4881\
        );

    \I__1009\ : Span4Mux_v
    port map (
            O => \N__4911\,
            I => \N__4878\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4871\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4909\,
            I => \N__4871\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4871\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4907\,
            I => \N__4868\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__4902\,
            I => \N__4865\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4901\,
            I => \N__4862\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4857\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4857\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4898\,
            I => \N__4854\
        );

    \I__999\ : Span4Mux_v
    port map (
            O => \N__4895\,
            I => \N__4845\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__4892\,
            I => \N__4845\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__4889\,
            I => \N__4845\
        );

    \I__996\ : Span4Mux_h
    port map (
            O => \N__4884\,
            I => \N__4845\
        );

    \I__995\ : Odrv4
    port map (
            O => \N__4881\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__4878\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4871\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__4868\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__991\ : Odrv12
    port map (
            O => \N__4865\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__4862\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4857\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4854\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__987\ : Odrv4
    port map (
            O => \N__4845\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__986\ : InMux
    port map (
            O => \N__4826\,
            I => \N__4823\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4823\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_2_1\
        );

    \I__984\ : InMux
    port map (
            O => \N__4820\,
            I => \N__4814\
        );

    \I__983\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4810\
        );

    \I__982\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4803\
        );

    \I__981\ : InMux
    port map (
            O => \N__4817\,
            I => \N__4800\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4814\,
            I => \N__4791\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__4813\,
            I => \N__4786\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4810\,
            I => \N__4782\
        );

    \I__977\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4775\
        );

    \I__976\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4775\
        );

    \I__975\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4775\
        );

    \I__974\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4770\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4803\,
            I => \N__4765\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4800\,
            I => \N__4765\
        );

    \I__971\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4760\
        );

    \I__970\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4760\
        );

    \I__969\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4757\
        );

    \I__968\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4754\
        );

    \I__967\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4751\
        );

    \I__966\ : InMux
    port map (
            O => \N__4794\,
            I => \N__4748\
        );

    \I__965\ : Span4Mux_h
    port map (
            O => \N__4791\,
            I => \N__4745\
        );

    \I__964\ : InMux
    port map (
            O => \N__4790\,
            I => \N__4742\
        );

    \I__963\ : InMux
    port map (
            O => \N__4789\,
            I => \N__4739\
        );

    \I__962\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4734\
        );

    \I__961\ : InMux
    port map (
            O => \N__4785\,
            I => \N__4734\
        );

    \I__960\ : Span4Mux_v
    port map (
            O => \N__4782\,
            I => \N__4731\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4775\,
            I => \N__4728\
        );

    \I__958\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4725\
        );

    \I__957\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4722\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4770\,
            I => \N__4717\
        );

    \I__955\ : Span4Mux_h
    port map (
            O => \N__4765\,
            I => \N__4717\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4760\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4757\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4754\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4751\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__4748\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__949\ : Odrv4
    port map (
            O => \N__4745\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4742\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4739\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4734\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__945\ : Odrv4
    port map (
            O => \N__4731\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__944\ : Odrv12
    port map (
            O => \N__4728\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4725\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4722\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__941\ : Odrv4
    port map (
            O => \N__4717\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__4688\,
            I => \N__4684\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__4687\,
            I => \N__4681\
        );

    \I__938\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4675\
        );

    \I__937\ : InMux
    port map (
            O => \N__4681\,
            I => \N__4672\
        );

    \I__936\ : InMux
    port map (
            O => \N__4680\,
            I => \N__4668\
        );

    \I__935\ : CascadeMux
    port map (
            O => \N__4679\,
            I => \N__4665\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__4678\,
            I => \N__4660\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4675\,
            I => \N__4656\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4672\,
            I => \N__4653\
        );

    \I__931\ : InMux
    port map (
            O => \N__4671\,
            I => \N__4650\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4668\,
            I => \N__4647\
        );

    \I__929\ : InMux
    port map (
            O => \N__4665\,
            I => \N__4640\
        );

    \I__928\ : InMux
    port map (
            O => \N__4664\,
            I => \N__4640\
        );

    \I__927\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4640\
        );

    \I__926\ : InMux
    port map (
            O => \N__4660\,
            I => \N__4635\
        );

    \I__925\ : InMux
    port map (
            O => \N__4659\,
            I => \N__4635\
        );

    \I__924\ : Span4Mux_v
    port map (
            O => \N__4656\,
            I => \N__4630\
        );

    \I__923\ : Span4Mux_v
    port map (
            O => \N__4653\,
            I => \N__4630\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__4650\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__4647\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4640\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__4635\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__918\ : Odrv4
    port map (
            O => \N__4630\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__4619\,
            I => \N__4612\
        );

    \I__916\ : InMux
    port map (
            O => \N__4618\,
            I => \N__4605\
        );

    \I__915\ : InMux
    port map (
            O => \N__4617\,
            I => \N__4602\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__4616\,
            I => \N__4599\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__4615\,
            I => \N__4593\
        );

    \I__912\ : InMux
    port map (
            O => \N__4612\,
            I => \N__4580\
        );

    \I__911\ : InMux
    port map (
            O => \N__4611\,
            I => \N__4580\
        );

    \I__910\ : InMux
    port map (
            O => \N__4610\,
            I => \N__4580\
        );

    \I__909\ : InMux
    port map (
            O => \N__4609\,
            I => \N__4575\
        );

    \I__908\ : InMux
    port map (
            O => \N__4608\,
            I => \N__4575\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4605\,
            I => \N__4569\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4602\,
            I => \N__4566\
        );

    \I__905\ : InMux
    port map (
            O => \N__4599\,
            I => \N__4561\
        );

    \I__904\ : InMux
    port map (
            O => \N__4598\,
            I => \N__4561\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__4597\,
            I => \N__4558\
        );

    \I__902\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4555\
        );

    \I__901\ : InMux
    port map (
            O => \N__4593\,
            I => \N__4550\
        );

    \I__900\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4550\
        );

    \I__899\ : InMux
    port map (
            O => \N__4591\,
            I => \N__4547\
        );

    \I__898\ : InMux
    port map (
            O => \N__4590\,
            I => \N__4540\
        );

    \I__897\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4540\
        );

    \I__896\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4540\
        );

    \I__895\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4537\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4580\,
            I => \N__4532\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4575\,
            I => \N__4532\
        );

    \I__892\ : InMux
    port map (
            O => \N__4574\,
            I => \N__4529\
        );

    \I__891\ : InMux
    port map (
            O => \N__4573\,
            I => \N__4524\
        );

    \I__890\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4524\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__4569\,
            I => \N__4517\
        );

    \I__888\ : Span4Mux_v
    port map (
            O => \N__4566\,
            I => \N__4517\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__4561\,
            I => \N__4517\
        );

    \I__886\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4514\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4555\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4550\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__4547\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4540\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__4537\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__880\ : Odrv4
    port map (
            O => \N__4532\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4529\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4524\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__877\ : Odrv4
    port map (
            O => \N__4517\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4514\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__875\ : InMux
    port map (
            O => \N__4493\,
            I => \N__4485\
        );

    \I__874\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4482\
        );

    \I__873\ : InMux
    port map (
            O => \N__4491\,
            I => \N__4479\
        );

    \I__872\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4474\
        );

    \I__871\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4474\
        );

    \I__870\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4470\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4485\,
            I => \N__4463\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4482\,
            I => \N__4463\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4479\,
            I => \N__4456\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4474\,
            I => \N__4456\
        );

    \I__865\ : InMux
    port map (
            O => \N__4473\,
            I => \N__4453\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4470\,
            I => \N__4450\
        );

    \I__863\ : InMux
    port map (
            O => \N__4469\,
            I => \N__4445\
        );

    \I__862\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4445\
        );

    \I__861\ : Span4Mux_v
    port map (
            O => \N__4463\,
            I => \N__4438\
        );

    \I__860\ : InMux
    port map (
            O => \N__4462\,
            I => \N__4435\
        );

    \I__859\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4432\
        );

    \I__858\ : Span4Mux_h
    port map (
            O => \N__4456\,
            I => \N__4429\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4453\,
            I => \N__4426\
        );

    \I__856\ : Span4Mux_v
    port map (
            O => \N__4450\,
            I => \N__4421\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4445\,
            I => \N__4421\
        );

    \I__854\ : InMux
    port map (
            O => \N__4444\,
            I => \N__4414\
        );

    \I__853\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4414\
        );

    \I__852\ : InMux
    port map (
            O => \N__4442\,
            I => \N__4414\
        );

    \I__851\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4411\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__4438\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4435\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4432\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__4429\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__846\ : Odrv4
    port map (
            O => \N__4426\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__845\ : Odrv4
    port map (
            O => \N__4421\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4414\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4411\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__842\ : InMux
    port map (
            O => \N__4394\,
            I => \N__4390\
        );

    \I__841\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4387\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4390\,
            I => \N__4382\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4387\,
            I => \N__4382\
        );

    \I__838\ : Span4Mux_h
    port map (
            O => \N__4382\,
            I => \N__4377\
        );

    \I__837\ : InMux
    port map (
            O => \N__4381\,
            I => \N__4374\
        );

    \I__836\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4371\
        );

    \I__835\ : Odrv4
    port map (
            O => \N__4377\,
            I => \U400_SDRAM.N_256\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4374\,
            I => \U400_SDRAM.N_256\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4371\,
            I => \U400_SDRAM.N_256\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__4364\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_a2_0_1_0_cascade_\
        );

    \I__831\ : InMux
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4358\,
            I => \N__4353\
        );

    \I__829\ : InMux
    port map (
            O => \N__4357\,
            I => \N__4350\
        );

    \I__828\ : InMux
    port map (
            O => \N__4356\,
            I => \N__4346\
        );

    \I__827\ : Span4Mux_v
    port map (
            O => \N__4353\,
            I => \N__4341\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4350\,
            I => \N__4341\
        );

    \I__825\ : InMux
    port map (
            O => \N__4349\,
            I => \N__4338\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4346\,
            I => \N__4328\
        );

    \I__823\ : Span4Mux_h
    port map (
            O => \N__4341\,
            I => \N__4325\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4338\,
            I => \N__4322\
        );

    \I__821\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4317\
        );

    \I__820\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4317\
        );

    \I__819\ : InMux
    port map (
            O => \N__4335\,
            I => \N__4308\
        );

    \I__818\ : InMux
    port map (
            O => \N__4334\,
            I => \N__4308\
        );

    \I__817\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4308\
        );

    \I__816\ : InMux
    port map (
            O => \N__4332\,
            I => \N__4308\
        );

    \I__815\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4305\
        );

    \I__814\ : Odrv4
    port map (
            O => \N__4328\,
            I => \U400_SDRAM.N_97\
        );

    \I__813\ : Odrv4
    port map (
            O => \N__4325\,
            I => \U400_SDRAM.N_97\
        );

    \I__812\ : Odrv4
    port map (
            O => \N__4322\,
            I => \U400_SDRAM.N_97\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4317\,
            I => \U400_SDRAM.N_97\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__4308\,
            I => \U400_SDRAM.N_97\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4305\,
            I => \U400_SDRAM.N_97\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__4292\,
            I => \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__4289\,
            I => \N__4285\
        );

    \I__806\ : InMux
    port map (
            O => \N__4288\,
            I => \N__4281\
        );

    \I__805\ : InMux
    port map (
            O => \N__4285\,
            I => \N__4273\
        );

    \I__804\ : InMux
    port map (
            O => \N__4284\,
            I => \N__4273\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4281\,
            I => \N__4270\
        );

    \I__802\ : InMux
    port map (
            O => \N__4280\,
            I => \N__4263\
        );

    \I__801\ : InMux
    port map (
            O => \N__4279\,
            I => \N__4263\
        );

    \I__800\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4263\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4273\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_2\
        );

    \I__798\ : Odrv4
    port map (
            O => \N__4270\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_2\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4263\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_2\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__4256\,
            I => \N__4250\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__4255\,
            I => \N__4246\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__4254\,
            I => \N__4243\
        );

    \I__793\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4240\
        );

    \I__792\ : InMux
    port map (
            O => \N__4250\,
            I => \N__4237\
        );

    \I__791\ : InMux
    port map (
            O => \N__4249\,
            I => \N__4230\
        );

    \I__790\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4230\
        );

    \I__789\ : InMux
    port map (
            O => \N__4243\,
            I => \N__4230\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4240\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_3\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4237\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_3\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4230\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_3\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__4223\,
            I => \N__4219\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__4222\,
            I => \N__4214\
        );

    \I__783\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4207\
        );

    \I__782\ : InMux
    port map (
            O => \N__4218\,
            I => \N__4207\
        );

    \I__781\ : InMux
    port map (
            O => \N__4217\,
            I => \N__4204\
        );

    \I__780\ : InMux
    port map (
            O => \N__4214\,
            I => \N__4197\
        );

    \I__779\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4197\
        );

    \I__778\ : InMux
    port map (
            O => \N__4212\,
            I => \N__4197\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4207\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4204\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4197\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__774\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4186\
        );

    \I__773\ : InMux
    port map (
            O => \N__4189\,
            I => \N__4183\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__4186\,
            I => \U400_SDRAM.CO1\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4183\,
            I => \U400_SDRAM.CO1\
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__4178\,
            I => \N__4174\
        );

    \I__769\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4168\
        );

    \I__768\ : InMux
    port map (
            O => \N__4174\,
            I => \N__4163\
        );

    \I__767\ : InMux
    port map (
            O => \N__4173\,
            I => \N__4163\
        );

    \I__766\ : InMux
    port map (
            O => \N__4172\,
            I => \N__4158\
        );

    \I__765\ : InMux
    port map (
            O => \N__4171\,
            I => \N__4158\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4168\,
            I => \U400_SDRAM.TA_COUNTER23\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__4163\,
            I => \U400_SDRAM.TA_COUNTER23\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4158\,
            I => \U400_SDRAM.TA_COUNTER23\
        );

    \I__761\ : InMux
    port map (
            O => \N__4151\,
            I => \N__4143\
        );

    \I__760\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4138\
        );

    \I__759\ : InMux
    port map (
            O => \N__4149\,
            I => \N__4138\
        );

    \I__758\ : InMux
    port map (
            O => \N__4148\,
            I => \N__4135\
        );

    \I__757\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4130\
        );

    \I__756\ : InMux
    port map (
            O => \N__4146\,
            I => \N__4130\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4143\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__4138\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4135\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__4130\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__4121\,
            I => \U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_\
        );

    \I__750\ : InMux
    port map (
            O => \N__4118\,
            I => \N__4112\
        );

    \I__749\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4112\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4112\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa\
        );

    \I__747\ : InMux
    port map (
            O => \N__4109\,
            I => \N__4095\
        );

    \I__746\ : InMux
    port map (
            O => \N__4108\,
            I => \N__4095\
        );

    \I__745\ : InMux
    port map (
            O => \N__4107\,
            I => \N__4095\
        );

    \I__744\ : InMux
    port map (
            O => \N__4106\,
            I => \N__4092\
        );

    \I__743\ : InMux
    port map (
            O => \N__4105\,
            I => \N__4083\
        );

    \I__742\ : InMux
    port map (
            O => \N__4104\,
            I => \N__4083\
        );

    \I__741\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4083\
        );

    \I__740\ : InMux
    port map (
            O => \N__4102\,
            I => \N__4083\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4095\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4092\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__4083\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__736\ : ClkMux
    port map (
            O => \N__4076\,
            I => \N__3995\
        );

    \I__735\ : ClkMux
    port map (
            O => \N__4075\,
            I => \N__3995\
        );

    \I__734\ : ClkMux
    port map (
            O => \N__4074\,
            I => \N__3995\
        );

    \I__733\ : ClkMux
    port map (
            O => \N__4073\,
            I => \N__3995\
        );

    \I__732\ : ClkMux
    port map (
            O => \N__4072\,
            I => \N__3995\
        );

    \I__731\ : ClkMux
    port map (
            O => \N__4071\,
            I => \N__3995\
        );

    \I__730\ : ClkMux
    port map (
            O => \N__4070\,
            I => \N__3995\
        );

    \I__729\ : ClkMux
    port map (
            O => \N__4069\,
            I => \N__3995\
        );

    \I__728\ : ClkMux
    port map (
            O => \N__4068\,
            I => \N__3995\
        );

    \I__727\ : ClkMux
    port map (
            O => \N__4067\,
            I => \N__3995\
        );

    \I__726\ : ClkMux
    port map (
            O => \N__4066\,
            I => \N__3995\
        );

    \I__725\ : ClkMux
    port map (
            O => \N__4065\,
            I => \N__3995\
        );

    \I__724\ : ClkMux
    port map (
            O => \N__4064\,
            I => \N__3995\
        );

    \I__723\ : ClkMux
    port map (
            O => \N__4063\,
            I => \N__3995\
        );

    \I__722\ : ClkMux
    port map (
            O => \N__4062\,
            I => \N__3995\
        );

    \I__721\ : ClkMux
    port map (
            O => \N__4061\,
            I => \N__3995\
        );

    \I__720\ : ClkMux
    port map (
            O => \N__4060\,
            I => \N__3995\
        );

    \I__719\ : ClkMux
    port map (
            O => \N__4059\,
            I => \N__3995\
        );

    \I__718\ : ClkMux
    port map (
            O => \N__4058\,
            I => \N__3995\
        );

    \I__717\ : ClkMux
    port map (
            O => \N__4057\,
            I => \N__3995\
        );

    \I__716\ : ClkMux
    port map (
            O => \N__4056\,
            I => \N__3995\
        );

    \I__715\ : ClkMux
    port map (
            O => \N__4055\,
            I => \N__3995\
        );

    \I__714\ : ClkMux
    port map (
            O => \N__4054\,
            I => \N__3995\
        );

    \I__713\ : ClkMux
    port map (
            O => \N__4053\,
            I => \N__3995\
        );

    \I__712\ : ClkMux
    port map (
            O => \N__4052\,
            I => \N__3995\
        );

    \I__711\ : ClkMux
    port map (
            O => \N__4051\,
            I => \N__3995\
        );

    \I__710\ : ClkMux
    port map (
            O => \N__4050\,
            I => \N__3995\
        );

    \I__709\ : GlobalMux
    port map (
            O => \N__3995\,
            I => \N__3992\
        );

    \I__708\ : gio2CtrlBuf
    port map (
            O => \N__3992\,
            I => \CLK40_c_g\
        );

    \I__707\ : InMux
    port map (
            O => \N__3989\,
            I => \N__3986\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3986\,
            I => \U400_SDRAM.N_189\
        );

    \I__705\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3977\
        );

    \I__704\ : InMux
    port map (
            O => \N__3982\,
            I => \N__3974\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__3981\,
            I => \N__3971\
        );

    \I__702\ : InMux
    port map (
            O => \N__3980\,
            I => \N__3962\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3977\,
            I => \N__3959\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__3974\,
            I => \N__3956\
        );

    \I__699\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3953\
        );

    \I__698\ : InMux
    port map (
            O => \N__3970\,
            I => \N__3943\
        );

    \I__697\ : InMux
    port map (
            O => \N__3969\,
            I => \N__3943\
        );

    \I__696\ : InMux
    port map (
            O => \N__3968\,
            I => \N__3943\
        );

    \I__695\ : InMux
    port map (
            O => \N__3967\,
            I => \N__3943\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__3966\,
            I => \N__3937\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__3965\,
            I => \N__3933\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__3962\,
            I => \N__3927\
        );

    \I__691\ : Span4Mux_v
    port map (
            O => \N__3959\,
            I => \N__3920\
        );

    \I__690\ : Span4Mux_v
    port map (
            O => \N__3956\,
            I => \N__3920\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3953\,
            I => \N__3920\
        );

    \I__688\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3917\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3943\,
            I => \N__3914\
        );

    \I__686\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3911\
        );

    \I__685\ : InMux
    port map (
            O => \N__3941\,
            I => \N__3908\
        );

    \I__684\ : InMux
    port map (
            O => \N__3940\,
            I => \N__3903\
        );

    \I__683\ : InMux
    port map (
            O => \N__3937\,
            I => \N__3903\
        );

    \I__682\ : InMux
    port map (
            O => \N__3936\,
            I => \N__3896\
        );

    \I__681\ : InMux
    port map (
            O => \N__3933\,
            I => \N__3896\
        );

    \I__680\ : InMux
    port map (
            O => \N__3932\,
            I => \N__3896\
        );

    \I__679\ : InMux
    port map (
            O => \N__3931\,
            I => \N__3893\
        );

    \I__678\ : InMux
    port map (
            O => \N__3930\,
            I => \N__3890\
        );

    \I__677\ : Span4Mux_v
    port map (
            O => \N__3927\,
            I => \N__3887\
        );

    \I__676\ : Span4Mux_h
    port map (
            O => \N__3920\,
            I => \N__3882\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3917\,
            I => \N__3882\
        );

    \I__674\ : Span4Mux_v
    port map (
            O => \N__3914\,
            I => \N__3877\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__3911\,
            I => \N__3877\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3908\,
            I => \N__3870\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3903\,
            I => \N__3870\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3896\,
            I => \N__3870\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3893\,
            I => \N__3865\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3890\,
            I => \N__3865\
        );

    \I__667\ : Span4Mux_h
    port map (
            O => \N__3887\,
            I => \N__3860\
        );

    \I__666\ : Span4Mux_v
    port map (
            O => \N__3882\,
            I => \N__3860\
        );

    \I__665\ : Span4Mux_v
    port map (
            O => \N__3877\,
            I => \N__3857\
        );

    \I__664\ : Span4Mux_v
    port map (
            O => \N__3870\,
            I => \N__3854\
        );

    \I__663\ : Span12Mux_s8_v
    port map (
            O => \N__3865\,
            I => \N__3851\
        );

    \I__662\ : Span4Mux_h
    port map (
            O => \N__3860\,
            I => \N__3848\
        );

    \I__661\ : Span4Mux_h
    port map (
            O => \N__3857\,
            I => \N__3845\
        );

    \I__660\ : Span4Mux_h
    port map (
            O => \N__3854\,
            I => \N__3842\
        );

    \I__659\ : Odrv12
    port map (
            O => \N__3851\,
            I => \RESETn_c\
        );

    \I__658\ : Odrv4
    port map (
            O => \N__3848\,
            I => \RESETn_c\
        );

    \I__657\ : Odrv4
    port map (
            O => \N__3845\,
            I => \RESETn_c\
        );

    \I__656\ : Odrv4
    port map (
            O => \N__3842\,
            I => \RESETn_c\
        );

    \I__655\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3830\,
            I => \N__3826\
        );

    \I__653\ : InMux
    port map (
            O => \N__3829\,
            I => \N__3823\
        );

    \I__652\ : Odrv4
    port map (
            O => \N__3826\,
            I => \U400_SDRAM.un1_REFRESH_COUNTERlto7_5\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3823\,
            I => \U400_SDRAM.un1_REFRESH_COUNTERlto7_5\
        );

    \I__650\ : InMux
    port map (
            O => \N__3818\,
            I => \N__3815\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3815\,
            I => \N__3811\
        );

    \I__648\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3808\
        );

    \I__647\ : Odrv4
    port map (
            O => \N__3811\,
            I => \U400_SDRAM.un1_REFRESH_COUNTERlto7_4\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3808\,
            I => \U400_SDRAM.un1_REFRESH_COUNTERlto7_4\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__3803\,
            I => \N__3800\
        );

    \I__644\ : InMux
    port map (
            O => \N__3800\,
            I => \N__3796\
        );

    \I__643\ : InMux
    port map (
            O => \N__3799\,
            I => \N__3793\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3796\,
            I => \N__3789\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3793\,
            I => \N__3786\
        );

    \I__640\ : InMux
    port map (
            O => \N__3792\,
            I => \N__3783\
        );

    \I__639\ : Span4Mux_h
    port map (
            O => \N__3789\,
            I => \N__3778\
        );

    \I__638\ : Span4Mux_h
    port map (
            O => \N__3786\,
            I => \N__3778\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__3783\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__3778\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\
        );

    \I__635\ : IoInMux
    port map (
            O => \N__3773\,
            I => \N__3770\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3770\,
            I => \N__3766\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__3769\,
            I => \N__3763\
        );

    \I__632\ : Span12Mux_s5_h
    port map (
            O => \N__3766\,
            I => \N__3760\
        );

    \I__631\ : InMux
    port map (
            O => \N__3763\,
            I => \N__3757\
        );

    \I__630\ : Odrv12
    port map (
            O => \N__3760\,
            I => \TA_OUT\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3757\,
            I => \TA_OUT\
        );

    \I__628\ : IoInMux
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3749\,
            I => \N__3746\
        );

    \I__626\ : Odrv4
    port map (
            O => \N__3746\,
            I => \N_66\
        );

    \I__625\ : CascadeMux
    port map (
            O => \N__3743\,
            I => \N__3740\
        );

    \I__624\ : InMux
    port map (
            O => \N__3740\,
            I => \N__3735\
        );

    \I__623\ : InMux
    port map (
            O => \N__3739\,
            I => \N__3732\
        );

    \I__622\ : InMux
    port map (
            O => \N__3738\,
            I => \N__3729\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3735\,
            I => \U400_SDRAM.BURSTZ0\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__3732\,
            I => \U400_SDRAM.BURSTZ0\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3729\,
            I => \U400_SDRAM.BURSTZ0\
        );

    \I__618\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3719\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3719\,
            I => \U400_SDRAM.TA_EN11_m\
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__3716\,
            I => \U400_SDRAM.un1_TA_COUNTER26_0_cascade_\
        );

    \I__615\ : InMux
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3710\,
            I => \U400_SDRAM.un1_TA_COUNTER26_2_0\
        );

    \I__613\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3703\
        );

    \I__612\ : InMux
    port map (
            O => \N__3706\,
            I => \N__3700\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3703\,
            I => \U400_SDRAM.TA_COUNTER27\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3700\,
            I => \U400_SDRAM.TA_COUNTER27\
        );

    \I__609\ : InMux
    port map (
            O => \N__3695\,
            I => \N__3692\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3692\,
            I => \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0\
        );

    \I__607\ : InMux
    port map (
            O => \N__3689\,
            I => \N__3686\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3686\,
            I => \N__3683\
        );

    \I__605\ : Odrv4
    port map (
            O => \N__3683\,
            I => \U400_SDRAM.N_207\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__3680\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_5_1_cascade_\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__3677\,
            I => \N__3674\
        );

    \I__602\ : InMux
    port map (
            O => \N__3674\,
            I => \N__3671\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3671\,
            I => \U400_SDRAM.N_250\
        );

    \I__600\ : CascadeMux
    port map (
            O => \N__3668\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_31_i_i_i_2_cascade_\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__3665\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_31_i_i_i_3_cascade_\
        );

    \I__598\ : InMux
    port map (
            O => \N__3662\,
            I => \N__3658\
        );

    \I__597\ : InMux
    port map (
            O => \N__3661\,
            I => \N__3655\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3658\,
            I => \U400_SDRAM.N_261\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3655\,
            I => \U400_SDRAM.N_261\
        );

    \I__594\ : InMux
    port map (
            O => \N__3650\,
            I => \N__3644\
        );

    \I__593\ : InMux
    port map (
            O => \N__3649\,
            I => \N__3644\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3644\,
            I => \U400_SDRAM.N_140\
        );

    \I__591\ : InMux
    port map (
            O => \N__3641\,
            I => \N__3638\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3638\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_4_1\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__3635\,
            I => \N__3632\
        );

    \I__588\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3628\
        );

    \I__587\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3625\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3628\,
            I => \N__3622\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3625\,
            I => \N__3619\
        );

    \I__584\ : Odrv4
    port map (
            O => \N__3622\,
            I => \U400_SDRAM.CS1_ENZ0\
        );

    \I__583\ : Odrv4
    port map (
            O => \N__3619\,
            I => \U400_SDRAM.CS1_ENZ0\
        );

    \I__582\ : IoInMux
    port map (
            O => \N__3614\,
            I => \N__3611\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3611\,
            I => \N__3608\
        );

    \I__580\ : Odrv12
    port map (
            O => \N__3608\,
            I => \CS1n_c\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__3605\,
            I => \N__3602\
        );

    \I__578\ : InMux
    port map (
            O => \N__3602\,
            I => \N__3599\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3599\,
            I => \N__3596\
        );

    \I__576\ : Span4Mux_v
    port map (
            O => \N__3596\,
            I => \N__3593\
        );

    \I__575\ : Span4Mux_v
    port map (
            O => \N__3593\,
            I => \N__3590\
        );

    \I__574\ : IoSpan4Mux
    port map (
            O => \N__3590\,
            I => \N__3587\
        );

    \I__573\ : Odrv4
    port map (
            O => \N__3587\,
            I => \A_c_26\
        );

    \I__572\ : IoInMux
    port map (
            O => \N__3584\,
            I => \N__3581\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3581\,
            I => \N__3578\
        );

    \I__570\ : Odrv12
    port map (
            O => \N__3578\,
            I => \MA_c_12\
        );

    \I__569\ : CascadeMux
    port map (
            O => \N__3575\,
            I => \U400_SDRAM.N_236_cascade_\
        );

    \I__568\ : InMux
    port map (
            O => \N__3572\,
            I => \N__3563\
        );

    \I__567\ : InMux
    port map (
            O => \N__3571\,
            I => \N__3563\
        );

    \I__566\ : InMux
    port map (
            O => \N__3570\,
            I => \N__3563\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__3563\,
            I => \U400_SDRAM.N_23_i\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__3560\,
            I => \U400_SDRAM.N_23_i_cascade_\
        );

    \I__563\ : InMux
    port map (
            O => \N__3557\,
            I => \N__3554\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3554\,
            I => \U400_SDRAM.N_242\
        );

    \I__561\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3545\
        );

    \I__560\ : InMux
    port map (
            O => \N__3550\,
            I => \N__3545\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3545\,
            I => \U400_SDRAM.N_139\
        );

    \I__558\ : InMux
    port map (
            O => \N__3542\,
            I => \N__3539\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3539\,
            I => \N__3536\
        );

    \I__556\ : Span4Mux_h
    port map (
            O => \N__3536\,
            I => \N__3533\
        );

    \I__555\ : Odrv4
    port map (
            O => \N__3533\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_1\
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__3530\,
            I => \N__3527\
        );

    \I__553\ : InMux
    port map (
            O => \N__3527\,
            I => \N__3524\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3524\,
            I => \U400_SDRAM.N_198\
        );

    \I__551\ : InMux
    port map (
            O => \N__3521\,
            I => \N__3515\
        );

    \I__550\ : InMux
    port map (
            O => \N__3520\,
            I => \N__3515\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3515\,
            I => \U400_SDRAM.N_259\
        );

    \I__548\ : CascadeMux
    port map (
            O => \N__3512\,
            I => \N__3508\
        );

    \I__547\ : InMux
    port map (
            O => \N__3511\,
            I => \N__3503\
        );

    \I__546\ : InMux
    port map (
            O => \N__3508\,
            I => \N__3503\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3503\,
            I => \U400_SDRAM.N_118\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__3500\,
            I => \N__3493\
        );

    \I__543\ : InMux
    port map (
            O => \N__3499\,
            I => \N__3487\
        );

    \I__542\ : InMux
    port map (
            O => \N__3498\,
            I => \N__3480\
        );

    \I__541\ : InMux
    port map (
            O => \N__3497\,
            I => \N__3480\
        );

    \I__540\ : InMux
    port map (
            O => \N__3496\,
            I => \N__3480\
        );

    \I__539\ : InMux
    port map (
            O => \N__3493\,
            I => \N__3475\
        );

    \I__538\ : InMux
    port map (
            O => \N__3492\,
            I => \N__3475\
        );

    \I__537\ : InMux
    port map (
            O => \N__3491\,
            I => \N__3470\
        );

    \I__536\ : InMux
    port map (
            O => \N__3490\,
            I => \N__3470\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3487\,
            I => \N__3467\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3480\,
            I => \U400_SDRAM.N_39\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3475\,
            I => \U400_SDRAM.N_39\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3470\,
            I => \U400_SDRAM.N_39\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__3467\,
            I => \U400_SDRAM.N_39\
        );

    \I__530\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3455\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3455\,
            I => \N__3452\
        );

    \I__528\ : Span4Mux_h
    port map (
            O => \N__3452\,
            I => \N__3449\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__3449\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_3\
        );

    \I__526\ : CEMux
    port map (
            O => \N__3446\,
            I => \N__3441\
        );

    \I__525\ : CEMux
    port map (
            O => \N__3445\,
            I => \N__3438\
        );

    \I__524\ : CEMux
    port map (
            O => \N__3444\,
            I => \N__3435\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3441\,
            I => \U400_SDRAM.N_219_i\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3438\,
            I => \U400_SDRAM.N_219_i\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3435\,
            I => \U400_SDRAM.N_219_i\
        );

    \I__520\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3425\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3425\,
            I => \N__3422\
        );

    \I__518\ : Span4Mux_h
    port map (
            O => \N__3422\,
            I => \N__3416\
        );

    \I__517\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3413\
        );

    \I__516\ : InMux
    port map (
            O => \N__3420\,
            I => \N__3410\
        );

    \I__515\ : InMux
    port map (
            O => \N__3419\,
            I => \N__3407\
        );

    \I__514\ : Odrv4
    port map (
            O => \N__3416\,
            I => \U400_SDRAM.N_239\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3413\,
            I => \U400_SDRAM.N_239\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3410\,
            I => \U400_SDRAM.N_239\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3407\,
            I => \U400_SDRAM.N_239\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__3398\,
            I => \N__3395\
        );

    \I__509\ : InMux
    port map (
            O => \N__3395\,
            I => \N__3392\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3392\,
            I => \N__3389\
        );

    \I__507\ : Span4Mux_v
    port map (
            O => \N__3389\,
            I => \N__3386\
        );

    \I__506\ : Sp12to4
    port map (
            O => \N__3386\,
            I => \N__3383\
        );

    \I__505\ : Odrv12
    port map (
            O => \N__3383\,
            I => \A_c_21\
        );

    \I__504\ : IoInMux
    port map (
            O => \N__3380\,
            I => \N__3377\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3377\,
            I => \N__3374\
        );

    \I__502\ : IoSpan4Mux
    port map (
            O => \N__3374\,
            I => \N__3371\
        );

    \I__501\ : Span4Mux_s3_h
    port map (
            O => \N__3371\,
            I => \N__3368\
        );

    \I__500\ : Span4Mux_v
    port map (
            O => \N__3368\,
            I => \N__3364\
        );

    \I__499\ : InMux
    port map (
            O => \N__3367\,
            I => \N__3361\
        );

    \I__498\ : Odrv4
    port map (
            O => \N__3364\,
            I => \BANK0_c\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3361\,
            I => \BANK0_c\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__3356\,
            I => \N__3353\
        );

    \I__495\ : InMux
    port map (
            O => \N__3353\,
            I => \N__3350\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3350\,
            I => \N__3347\
        );

    \I__493\ : Span12Mux_s9_h
    port map (
            O => \N__3347\,
            I => \N__3344\
        );

    \I__492\ : Odrv12
    port map (
            O => \N__3344\,
            I => \A_c_22\
        );

    \I__491\ : InMux
    port map (
            O => \N__3341\,
            I => \N__3337\
        );

    \I__490\ : InMux
    port map (
            O => \N__3340\,
            I => \N__3334\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3337\,
            I => \U400_SDRAM.N_240\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3334\,
            I => \U400_SDRAM.N_240\
        );

    \I__487\ : IoInMux
    port map (
            O => \N__3329\,
            I => \N__3326\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3326\,
            I => \N__3323\
        );

    \I__485\ : IoSpan4Mux
    port map (
            O => \N__3323\,
            I => \N__3320\
        );

    \I__484\ : IoSpan4Mux
    port map (
            O => \N__3320\,
            I => \N__3317\
        );

    \I__483\ : Span4Mux_s3_h
    port map (
            O => \N__3317\,
            I => \N__3313\
        );

    \I__482\ : InMux
    port map (
            O => \N__3316\,
            I => \N__3310\
        );

    \I__481\ : Odrv4
    port map (
            O => \N__3313\,
            I => \BANK1_c\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3310\,
            I => \BANK1_c\
        );

    \I__479\ : InMux
    port map (
            O => \N__3305\,
            I => \N__3302\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3302\,
            I => \N__3299\
        );

    \I__477\ : Span12Mux_v
    port map (
            O => \N__3299\,
            I => \N__3296\
        );

    \I__476\ : Odrv12
    port map (
            O => \N__3296\,
            I => \RnW_c\
        );

    \I__475\ : InMux
    port map (
            O => \N__3293\,
            I => \N__3290\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3290\,
            I => \U400_SDRAM.N_82\
        );

    \I__473\ : InMux
    port map (
            O => \N__3287\,
            I => \N__3284\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3284\,
            I => \U400_SDRAM.N_34\
        );

    \I__471\ : CascadeMux
    port map (
            O => \N__3281\,
            I => \U400_SDRAM.N_118_cascade_\
        );

    \I__470\ : InMux
    port map (
            O => \N__3278\,
            I => \N__3275\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3275\,
            I => \U400_SDRAM.N_215\
        );

    \I__468\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3268\
        );

    \I__467\ : InMux
    port map (
            O => \N__3271\,
            I => \N__3265\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3268\,
            I => \U400_SDRAM.RAM_CYCLEZ0\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3265\,
            I => \U400_SDRAM.RAM_CYCLEZ0\
        );

    \I__464\ : InMux
    port map (
            O => \N__3260\,
            I => \N__3251\
        );

    \I__463\ : InMux
    port map (
            O => \N__3259\,
            I => \N__3251\
        );

    \I__462\ : InMux
    port map (
            O => \N__3258\,
            I => \N__3251\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__3251\,
            I => \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3Z0Z_0\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__3248\,
            I => \U400_SDRAM.N_230_cascade_\
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__3245\,
            I => \N__3242\
        );

    \I__458\ : InMux
    port map (
            O => \N__3242\,
            I => \N__3239\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3239\,
            I => \N__3236\
        );

    \I__456\ : Sp12to4
    port map (
            O => \N__3236\,
            I => \N__3233\
        );

    \I__455\ : Span12Mux_s10_v
    port map (
            O => \N__3233\,
            I => \N__3230\
        );

    \I__454\ : Odrv12
    port map (
            O => \N__3230\,
            I => \A_c_19\
        );

    \I__453\ : IoInMux
    port map (
            O => \N__3227\,
            I => \N__3224\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3224\,
            I => \N__3221\
        );

    \I__451\ : Odrv12
    port map (
            O => \N__3221\,
            I => \MA_c_9\
        );

    \I__450\ : InMux
    port map (
            O => \N__3218\,
            I => \N__3215\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3215\,
            I => \A_c_30\
        );

    \I__448\ : InMux
    port map (
            O => \N__3212\,
            I => \N__3209\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3209\,
            I => \N__3206\
        );

    \I__446\ : Span12Mux_s10_h
    port map (
            O => \N__3206\,
            I => \N__3203\
        );

    \I__445\ : Odrv12
    port map (
            O => \N__3203\,
            I => \A_c_29\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__3200\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_\
        );

    \I__443\ : InMux
    port map (
            O => \N__3197\,
            I => \N__3194\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__3194\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en\
        );

    \I__441\ : CEMux
    port map (
            O => \N__3191\,
            I => \N__3188\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3188\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__3185\,
            I => \U400_SDRAM.CS0_EN_0_cascade_\
        );

    \I__438\ : InMux
    port map (
            O => \N__3182\,
            I => \N__3178\
        );

    \I__437\ : InMux
    port map (
            O => \N__3181\,
            I => \N__3175\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3178\,
            I => \U400_SDRAM.CS0_ENZ0\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__3175\,
            I => \U400_SDRAM.CS0_ENZ0\
        );

    \I__434\ : CascadeMux
    port map (
            O => \N__3170\,
            I => \N__3166\
        );

    \I__433\ : CascadeMux
    port map (
            O => \N__3169\,
            I => \N__3163\
        );

    \I__432\ : InMux
    port map (
            O => \N__3166\,
            I => \N__3158\
        );

    \I__431\ : InMux
    port map (
            O => \N__3163\,
            I => \N__3158\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3158\,
            I => \N__3155\
        );

    \I__429\ : Span4Mux_v
    port map (
            O => \N__3155\,
            I => \N__3152\
        );

    \I__428\ : Odrv4
    port map (
            O => \N__3152\,
            I => \A_c_23\
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__3149\,
            I => \U400_SDRAM.CS1_EN_0_cascade_\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__3146\,
            I => \U400_SDRAM.N_114_cascade_\
        );

    \I__425\ : InMux
    port map (
            O => \N__3143\,
            I => \N__3140\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3140\,
            I => \U400_SDRAM.N_220\
        );

    \I__423\ : InMux
    port map (
            O => \N__3137\,
            I => \N__3134\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3134\,
            I => \U400_SDRAM.N_258\
        );

    \I__421\ : InMux
    port map (
            O => \N__3131\,
            I => \N__3128\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3128\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_0_1\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__3125\,
            I => \U400_SDRAM.N_258_cascade_\
        );

    \I__418\ : InMux
    port map (
            O => \N__3122\,
            I => \N__3119\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3119\,
            I => \N__3116\
        );

    \I__416\ : Span4Mux_h
    port map (
            O => \N__3116\,
            I => \N__3113\
        );

    \I__415\ : Odrv4
    port map (
            O => \N__3113\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_0_0\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__3110\,
            I => \U400_SDRAM.N_240_cascade_\
        );

    \I__413\ : InMux
    port map (
            O => \N__3107\,
            I => \N__3103\
        );

    \I__412\ : InMux
    port map (
            O => \N__3106\,
            I => \N__3100\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3103\,
            I => \N__3097\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3100\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__409\ : Odrv4
    port map (
            O => \N__3097\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__408\ : InMux
    port map (
            O => \N__3092\,
            I => \N__3088\
        );

    \I__407\ : InMux
    port map (
            O => \N__3091\,
            I => \N__3085\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3088\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__3085\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__404\ : CascadeMux
    port map (
            O => \N__3080\,
            I => \N__3076\
        );

    \I__403\ : InMux
    port map (
            O => \N__3079\,
            I => \N__3073\
        );

    \I__402\ : InMux
    port map (
            O => \N__3076\,
            I => \N__3070\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__3073\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3070\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__399\ : InMux
    port map (
            O => \N__3065\,
            I => \N__3060\
        );

    \I__398\ : InMux
    port map (
            O => \N__3064\,
            I => \N__3055\
        );

    \I__397\ : InMux
    port map (
            O => \N__3063\,
            I => \N__3055\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3060\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__3055\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__394\ : InMux
    port map (
            O => \N__3050\,
            I => \N__3046\
        );

    \I__393\ : InMux
    port map (
            O => \N__3049\,
            I => \N__3043\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__3046\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__3043\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__390\ : InMux
    port map (
            O => \N__3038\,
            I => \N__3034\
        );

    \I__389\ : InMux
    port map (
            O => \N__3037\,
            I => \N__3031\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3034\,
            I => \N__3028\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3031\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__386\ : Odrv4
    port map (
            O => \N__3028\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__385\ : CascadeMux
    port map (
            O => \N__3023\,
            I => \N__3019\
        );

    \I__384\ : InMux
    port map (
            O => \N__3022\,
            I => \N__3016\
        );

    \I__383\ : InMux
    port map (
            O => \N__3019\,
            I => \N__3013\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3016\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__3013\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__380\ : CascadeMux
    port map (
            O => \N__3008\,
            I => \N__3004\
        );

    \I__379\ : CascadeMux
    port map (
            O => \N__3007\,
            I => \N__3001\
        );

    \I__378\ : InMux
    port map (
            O => \N__3004\,
            I => \N__2996\
        );

    \I__377\ : InMux
    port map (
            O => \N__3001\,
            I => \N__2989\
        );

    \I__376\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2989\
        );

    \I__375\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2989\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__2996\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2989\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__372\ : SRMux
    port map (
            O => \N__2984\,
            I => \N__2981\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2981\,
            I => \N__2977\
        );

    \I__370\ : SRMux
    port map (
            O => \N__2980\,
            I => \N__2974\
        );

    \I__369\ : Span4Mux_h
    port map (
            O => \N__2977\,
            I => \N__2971\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2974\,
            I => \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2\
        );

    \I__367\ : Odrv4
    port map (
            O => \N__2971\,
            I => \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2\
        );

    \I__366\ : InMux
    port map (
            O => \N__2966\,
            I => \N__2963\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2963\,
            I => \N__2960\
        );

    \I__364\ : Odrv12
    port map (
            O => \N__2960\,
            I => \A_c_8\
        );

    \I__363\ : CascadeMux
    port map (
            O => \N__2957\,
            I => \N__2954\
        );

    \I__362\ : InMux
    port map (
            O => \N__2954\,
            I => \N__2951\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2951\,
            I => \N__2948\
        );

    \I__360\ : Span4Mux_v
    port map (
            O => \N__2948\,
            I => \N__2945\
        );

    \I__359\ : Span4Mux_v
    port map (
            O => \N__2945\,
            I => \N__2942\
        );

    \I__358\ : Odrv4
    port map (
            O => \N__2942\,
            I => \A_c_16\
        );

    \I__357\ : IoInMux
    port map (
            O => \N__2939\,
            I => \N__2936\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2936\,
            I => \N__2933\
        );

    \I__355\ : Odrv4
    port map (
            O => \N__2933\,
            I => \MA_c_6\
        );

    \I__354\ : InMux
    port map (
            O => \N__2930\,
            I => \N__2927\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__2927\,
            I => \U400_SDRAM.N_216\
        );

    \I__352\ : InMux
    port map (
            O => \N__2924\,
            I => \N__2921\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2921\,
            I => \N__2917\
        );

    \I__350\ : InMux
    port map (
            O => \N__2920\,
            I => \N__2914\
        );

    \I__349\ : Odrv4
    port map (
            O => \N__2917\,
            I => \U400_SDRAM.N_187\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2914\,
            I => \U400_SDRAM.N_187\
        );

    \I__347\ : InMux
    port map (
            O => \N__2909\,
            I => \N__2906\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2906\,
            I => \N__2903\
        );

    \I__345\ : Odrv4
    port map (
            O => \N__2903\,
            I => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_2_0\
        );

    \I__344\ : CascadeMux
    port map (
            O => \N__2900\,
            I => \N__2897\
        );

    \I__343\ : InMux
    port map (
            O => \N__2897\,
            I => \N__2894\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2894\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_0\
        );

    \I__341\ : InMux
    port map (
            O => \N__2891\,
            I => \N__2888\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2888\,
            I => \U400_SDRAM.TACK_7_iv_i_i_2\
        );

    \I__339\ : CascadeMux
    port map (
            O => \N__2885\,
            I => \U400_SDRAM.TACK_7_iv_i_i_1_0_cascade_\
        );

    \I__338\ : IoInMux
    port map (
            O => \N__2882\,
            I => \N__2879\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2879\,
            I => \N__2876\
        );

    \I__336\ : Span4Mux_s3_h
    port map (
            O => \N__2876\,
            I => \N__2873\
        );

    \I__335\ : Odrv4
    port map (
            O => \N__2873\,
            I => \CS0n_c\
        );

    \I__334\ : IoInMux
    port map (
            O => \N__2870\,
            I => \N__2867\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2867\,
            I => \N__2864\
        );

    \I__332\ : Odrv12
    port map (
            O => \N__2864\,
            I => \CASn_c\
        );

    \I__331\ : IoInMux
    port map (
            O => \N__2861\,
            I => \N__2858\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2858\,
            I => \N__2855\
        );

    \I__329\ : Odrv12
    port map (
            O => \N__2855\,
            I => \WEn_c\
        );

    \I__328\ : IoInMux
    port map (
            O => \N__2852\,
            I => \N__2849\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2849\,
            I => \N__2846\
        );

    \I__326\ : Odrv12
    port map (
            O => \N__2846\,
            I => \RASn_c\
        );

    \I__325\ : InMux
    port map (
            O => \N__2843\,
            I => \N__2840\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2840\,
            I => \N__2837\
        );

    \I__323\ : Span4Mux_h
    port map (
            O => \N__2837\,
            I => \N__2834\
        );

    \I__322\ : Sp12to4
    port map (
            O => \N__2834\,
            I => \N__2831\
        );

    \I__321\ : Span12Mux_v
    port map (
            O => \N__2831\,
            I => \N__2828\
        );

    \I__320\ : Odrv12
    port map (
            O => \N__2828\,
            I => \A_c_24\
        );

    \I__319\ : CascadeMux
    port map (
            O => \N__2825\,
            I => \N__2822\
        );

    \I__318\ : InMux
    port map (
            O => \N__2822\,
            I => \N__2819\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2819\,
            I => \N__2816\
        );

    \I__316\ : Span12Mux_s10_v
    port map (
            O => \N__2816\,
            I => \N__2813\
        );

    \I__315\ : Odrv12
    port map (
            O => \N__2813\,
            I => \A_c_18\
        );

    \I__314\ : IoInMux
    port map (
            O => \N__2810\,
            I => \N__2807\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2807\,
            I => \N__2804\
        );

    \I__312\ : Span4Mux_s1_v
    port map (
            O => \N__2804\,
            I => \N__2801\
        );

    \I__311\ : Odrv4
    port map (
            O => \N__2801\,
            I => \MA_c_8\
        );

    \I__310\ : InMux
    port map (
            O => \N__2798\,
            I => \N__2795\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2795\,
            I => \N__2792\
        );

    \I__308\ : Odrv12
    port map (
            O => \N__2792\,
            I => \A_c_9\
        );

    \I__307\ : CascadeMux
    port map (
            O => \N__2789\,
            I => \N__2786\
        );

    \I__306\ : InMux
    port map (
            O => \N__2786\,
            I => \N__2783\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2783\,
            I => \N__2780\
        );

    \I__304\ : Span4Mux_v
    port map (
            O => \N__2780\,
            I => \N__2777\
        );

    \I__303\ : Odrv4
    port map (
            O => \N__2777\,
            I => \A_c_17\
        );

    \I__302\ : IoInMux
    port map (
            O => \N__2774\,
            I => \N__2771\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2771\,
            I => \N__2768\
        );

    \I__300\ : Span4Mux_s1_v
    port map (
            O => \N__2768\,
            I => \N__2765\
        );

    \I__299\ : Odrv4
    port map (
            O => \N__2765\,
            I => \MA_c_7\
        );

    \I__298\ : InMux
    port map (
            O => \N__2762\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_4\
        );

    \I__297\ : InMux
    port map (
            O => \N__2759\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_5\
        );

    \I__296\ : InMux
    port map (
            O => \N__2756\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_6\
        );

    \I__295\ : InMux
    port map (
            O => \N__2753\,
            I => \N__2750\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2750\,
            I => \N__2747\
        );

    \I__293\ : Odrv4
    port map (
            O => \N__2747\,
            I => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_0_0\
        );

    \I__292\ : CascadeMux
    port map (
            O => \N__2744\,
            I => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a2_1_0_cascade_\
        );

    \I__291\ : InMux
    port map (
            O => \N__2741\,
            I => \N__2737\
        );

    \I__290\ : InMux
    port map (
            O => \N__2740\,
            I => \N__2734\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2737\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2734\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__287\ : InMux
    port map (
            O => \N__2729\,
            I => \N__2725\
        );

    \I__286\ : InMux
    port map (
            O => \N__2728\,
            I => \N__2722\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2725\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2722\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__283\ : CascadeMux
    port map (
            O => \N__2717\,
            I => \N__2713\
        );

    \I__282\ : InMux
    port map (
            O => \N__2716\,
            I => \N__2710\
        );

    \I__281\ : InMux
    port map (
            O => \N__2713\,
            I => \N__2707\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2710\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2707\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__278\ : InMux
    port map (
            O => \N__2702\,
            I => \N__2698\
        );

    \I__277\ : InMux
    port map (
            O => \N__2701\,
            I => \N__2695\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2698\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2695\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__274\ : CascadeMux
    port map (
            O => \N__2690\,
            I => \U400_SDRAM.N_97_cascade_\
        );

    \I__273\ : CascadeMux
    port map (
            O => \N__2687\,
            I => \U400_SDRAM.N_256_cascade_\
        );

    \I__272\ : InMux
    port map (
            O => \N__2684\,
            I => \N__2681\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2681\,
            I => \N__2677\
        );

    \I__270\ : InMux
    port map (
            O => \N__2680\,
            I => \N__2674\
        );

    \I__269\ : Odrv4
    port map (
            O => \N__2677\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2674\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__267\ : InMux
    port map (
            O => \N__2669\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_4\
        );

    \I__266\ : InMux
    port map (
            O => \N__2666\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_5\
        );

    \I__265\ : InMux
    port map (
            O => \N__2663\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_6\
        );

    \I__264\ : InMux
    port map (
            O => \N__2660\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_7\
        );

    \I__263\ : InMux
    port map (
            O => \N__2657\,
            I => \bfn_4_6_0_\
        );

    \I__262\ : InMux
    port map (
            O => \N__2654\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_0\
        );

    \I__261\ : InMux
    port map (
            O => \N__2651\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_1\
        );

    \I__260\ : InMux
    port map (
            O => \N__2648\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_2\
        );

    \I__259\ : InMux
    port map (
            O => \N__2645\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_3\
        );

    \I__258\ : IoInMux
    port map (
            O => \N__2642\,
            I => \N__2639\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2639\,
            I => \RESETn_c_i\
        );

    \I__256\ : IoInMux
    port map (
            O => \N__2636\,
            I => \N__2633\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2633\,
            I => \CONSTANT_ONE_NET\
        );

    \I__254\ : InMux
    port map (
            O => \N__2630\,
            I => \N__2627\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2627\,
            I => \N__2624\
        );

    \I__252\ : Odrv12
    port map (
            O => \N__2624\,
            I => \A_c_27\
        );

    \I__251\ : InMux
    port map (
            O => \N__2621\,
            I => \N__2618\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2618\,
            I => \N__2615\
        );

    \I__249\ : Odrv4
    port map (
            O => \N__2615\,
            I => \A_c_28\
        );

    \I__248\ : CascadeMux
    port map (
            O => \N__2612\,
            I => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a2_1_0_0_cascade_\
        );

    \I__247\ : InMux
    port map (
            O => \N__2609\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_1\
        );

    \I__246\ : InMux
    port map (
            O => \N__2606\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_2\
        );

    \I__245\ : InMux
    port map (
            O => \N__2603\,
            I => \U400_SDRAM.un2_REFRESH_COUNTER_cry_3\
        );

    \I__244\ : IoInMux
    port map (
            O => \N__2600\,
            I => \N__2597\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__2597\,
            I => \N__2594\
        );

    \I__242\ : IoSpan4Mux
    port map (
            O => \N__2594\,
            I => \N__2591\
        );

    \I__241\ : IoSpan4Mux
    port map (
            O => \N__2591\,
            I => \N__2588\
        );

    \I__240\ : Span4Mux_s2_h
    port map (
            O => \N__2588\,
            I => \N__2585\
        );

    \I__239\ : Sp12to4
    port map (
            O => \N__2585\,
            I => \N__2582\
        );

    \I__238\ : Odrv12
    port map (
            O => \N__2582\,
            I => \CLK40_ibuf_gb_io_gb_input\
        );

    \INVU400_SDRAM.MA_nesr_2C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_2C_net\,
            I => \N__4076\
        );

    \INVU400_SDRAM.MA_nesr_3C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_3C_net\,
            I => \N__4075\
        );

    \INVU400_SDRAM.MA_nesr_10C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_10C_net\,
            I => \N__4072\
        );

    \INVU400_SDRAM.MA_nesr_5C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_5C_net\,
            I => \N__4073\
        );

    \INVU400_SDRAM.MA_nesr_11C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_11C_net\,
            I => \N__4069\
        );

    \INVU400_SDRAM.SDRAM_CMD_ne_0C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_ne_0C_net\,
            I => \N__4062\
        );

    \INVU400_SDRAM.MA_nesr_12C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_12C_net\,
            I => \N__4066\
        );

    \INVU400_SDRAM.CS1nC\ : INV
    port map (
            O => \INVU400_SDRAM.CS1nC_net\,
            I => \N__4053\
        );

    \INVU400_SDRAM.SDRAM_CMD_1C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_1C_net\,
            I => \N__4057\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_1C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_1C_net\,
            I => \N__4061\
        );

    \INVU400_SDRAM.BANK0C\ : INV
    port map (
            O => \INVU400_SDRAM.BANK0C_net\,
            I => \N__4068\
        );

    \INVU400_SDRAM.MA_nesr_9C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_9C_net\,
            I => \N__4059\
        );

    \INVU400_SDRAM.CS0_ENC\ : INV
    port map (
            O => \INVU400_SDRAM.CS0_ENC_net\,
            I => \N__4056\
        );

    \INVU400_SDRAM.REFRESH_COUNTER_1C\ : INV
    port map (
            O => \INVU400_SDRAM.REFRESH_COUNTER_1C_net\,
            I => \N__4060\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_0C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            I => \N__4065\
        );

    \INVU400_SDRAM.MA_nesr_6C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_6C_net\,
            I => \N__4063\
        );

    \INVU400_SDRAM.MA_nesr_8C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_8C_net\,
            I => \N__4054\
        );

    \INVU400_SDRAM.RASnC\ : INV
    port map (
            O => \INVU400_SDRAM.RASnC_net\,
            I => \N__4051\
        );

    \INVU400_SDRAM.CASnC\ : INV
    port map (
            O => \INVU400_SDRAM.CASnC_net\,
            I => \N__4050\
        );

    \INVU400_SDRAM.CS0nC\ : INV
    port map (
            O => \INVU400_SDRAM.CS0nC_net\,
            I => \N__4052\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_2C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            I => \N__4055\
        );

    \INVU400_SDRAM.REFRESH_COUNTER_2C\ : INV
    port map (
            O => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            I => \N__4058\
        );

    \INVU400_SDRAM.SDRAM_CONFIGUREDC\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CONFIGUREDC_net\,
            I => \N__4064\
        );

    \IN_MUX_bfv_4_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_5_0_\
        );

    \IN_MUX_bfv_4_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_6_0_\
        );

    \CLK40_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2600\,
            GLOBALBUFFEROUTPUT => \CLK40_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2642\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3980\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2_2_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__2630\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2621\,
            lcout => \U400_ADDRESS_DECODE_RAM_SPACE_i_o3_0_o2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5457\,
            in2 => \_gnd_net_\,
            in3 => \N__2684\,
            lcout => \U400_SDRAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CONFIGUREDC_net\,
            ce => 'H',
            sr => \N__6163\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_5_0_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4817\,
            in1 => \N__4617\,
            in2 => \_gnd_net_\,
            in3 => \N__4898\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a2_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111010101"
        )
    port map (
            in0 => \N__3931\,
            in1 => \N__5456\,
            in2 => \N__2612\,
            in3 => \N__4349\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.un2_REFRESH_COUNTER_cry_1_c_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3065\,
            in2 => \N__3008\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_5_0_\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_2_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3092\,
            in2 => \_gnd_net_\,
            in3 => \N__2609\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un2_REFRESH_COUNTER_cry_1\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_2\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__2984\
        );

    \U400_SDRAM.REFRESH_COUNTER_3_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3106\,
            in2 => \_gnd_net_\,
            in3 => \N__2606\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un2_REFRESH_COUNTER_cry_2\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_3\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__2984\
        );

    \U400_SDRAM.REFRESH_COUNTER_4_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3079\,
            in2 => \_gnd_net_\,
            in3 => \N__2603\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un2_REFRESH_COUNTER_cry_3\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_4\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__2984\
        );

    \U400_SDRAM.REFRESH_COUNTER_5_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3050\,
            in2 => \_gnd_net_\,
            in3 => \N__2669\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un2_REFRESH_COUNTER_cry_4\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_5\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__2984\
        );

    \U400_SDRAM.REFRESH_COUNTER_6_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3037\,
            in2 => \_gnd_net_\,
            in3 => \N__2666\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un2_REFRESH_COUNTER_cry_5\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_6\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__2984\
        );

    \U400_SDRAM.REFRESH_COUNTER_7_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3022\,
            in2 => \_gnd_net_\,
            in3 => \N__2663\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un2_REFRESH_COUNTER_cry_6\,
            carryout => \U400_SDRAM.un2_REFRESH_COUNTER_cry_7\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__2984\
        );

    \U400_SDRAM.REFRESH_COUNTER_8_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3792\,
            in2 => \_gnd_net_\,
            in3 => \N__2660\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__2984\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4907\,
            in2 => \_gnd_net_\,
            in3 => \N__2657\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \bfn_4_6_0_\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4819\,
            in2 => \_gnd_net_\,
            in3 => \N__2654\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_1\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_0\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_2_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3496\,
            in1 => \N__4462\,
            in2 => \_gnd_net_\,
            in3 => \N__2651\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_1\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_2\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4618\,
            in2 => \_gnd_net_\,
            in3 => \N__2648\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_3\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_2\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_4_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3497\,
            in1 => \N__2702\,
            in2 => \_gnd_net_\,
            in3 => \N__2645\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_3\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_4\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_5_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3490\,
            in1 => \N__2729\,
            in2 => \_gnd_net_\,
            in3 => \N__2762\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_4\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_5\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_6_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3498\,
            in1 => \N__2741\,
            in2 => \_gnd_net_\,
            in3 => \N__2759\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_5\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_6\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_7_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3491\,
            in1 => \N__2716\,
            in2 => \_gnd_net_\,
            in3 => \N__2756\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__3444\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5516\,
            in1 => \N__2924\,
            in2 => \_gnd_net_\,
            in3 => \N__4444\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_a2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__2753\,
            in1 => \N__3420\,
            in2 => \N__2744\,
            in3 => \N__2680\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2740\,
            in1 => \N__2728\,
            in2 => \N__2717\,
            in3 => \N__2701\,
            lcout => \U400_SDRAM.N_97\,
            ltout => \U400_SDRAM.N_97_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_0_2_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__4442\,
            in1 => \N__4598\,
            in2 => \N__2690\,
            in3 => \N__4926\,
            lcout => \U400_SDRAM.N_256\,
            ltout => \U400_SDRAM.N_256_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5523\,
            in2 => \N__2687\,
            in3 => \N__4808\,
            lcout => \U400_SDRAM.SDRAM_CMD_3_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCA2_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110110011"
        )
    port map (
            in0 => \N__4809\,
            in1 => \N__3930\,
            in2 => \N__5547\,
            in3 => \N__5396\,
            lcout => \U400_SDRAM.SDRAM_CONFIGURED_RNIJKCAZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_2_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__4337\,
            in1 => \N__5522\,
            in2 => \N__4616\,
            in3 => \N__4443\,
            lcout => \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIE9F21_1_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4807\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4336\,
            lcout => \U400_SDRAM.N_239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS0n_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000000011111111"
        )
    port map (
            in0 => \N__6450\,
            in1 => \N__6067\,
            in2 => \N__5969\,
            in3 => \N__3182\,
            lcout => \CS0n_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0nC_net\,
            ce => 'H',
            sr => \N__6157\
        );

    \U400_SDRAM.CASn_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6069\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CASnC_net\,
            ce => 'H',
            sr => \N__6158\
        );

    \U400_SDRAM.WEn_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5967\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CASnC_net\,
            ce => 'H',
            sr => \N__6158\
        );

    \U400_SDRAM.RASn_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6489\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RASnC_net\,
            ce => 'H',
            sr => \N__6159\
        );

    \U400_SDRAM.MA_nesr_8_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__6491\,
            in1 => \N__2843\,
            in2 => \N__2825\,
            in3 => \N__6332\,
            lcout => \MA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_8C_net\,
            ce => \N__6268\,
            sr => \N__6162\
        );

    \U400_SDRAM.MA_nesr_7_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__6490\,
            in1 => \N__2798\,
            in2 => \N__2789\,
            in3 => \N__6331\,
            lcout => \MA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_8C_net\,
            ce => \N__6268\,
            sr => \N__6162\
        );

    \U400_SDRAM.MA_nesr_6_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__2966\,
            in1 => \N__6503\,
            in2 => \N__2957\,
            in3 => \N__6338\,
            lcout => \MA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_6C_net\,
            ce => \N__6269\,
            sr => \N__6169\
        );

    \U400_SDRAM.TACK_RNO_3_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__2930\,
            in1 => \N__2920\,
            in2 => \_gnd_net_\,
            in3 => \N__4488\,
            lcout => \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6187\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3197\,
            lcout => \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_6_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__4818\,
            in1 => \N__4900\,
            in2 => \N__4678\,
            in3 => \N__4609\,
            lcout => \U400_SDRAM.N_216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_RNI07LH_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__4659\,
            in1 => \N__4899\,
            in2 => \_gnd_net_\,
            in3 => \N__4608\,
            lcout => \U400_SDRAM.N_187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_0_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__3278\,
            in1 => \N__2909\,
            in2 => \N__2900\,
            in3 => \N__3499\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            ce => \N__3445\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_5_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100010"
        )
    port map (
            in0 => \N__4908\,
            in1 => \N__4664\,
            in2 => \N__4619\,
            in3 => \N__4461\,
            lcout => \U400_SDRAM.TACK_7_iv_i_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_4_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010101001110"
        )
    port map (
            in0 => \N__4820\,
            in1 => \N__4611\,
            in2 => \N__4679\,
            in3 => \N__4909\,
            lcout => OPEN,
            ltout => \U400_SDRAM.TACK_7_iv_i_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_1_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__2891\,
            in1 => \N__3137\,
            in2 => \N__2885\,
            in3 => \N__4356\,
            lcout => \U400_SDRAM.N_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_RNI18LH_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4663\,
            in1 => \N__4806\,
            in2 => \_gnd_net_\,
            in3 => \N__4610\,
            lcout => \U400_SDRAM.N_258\,
            ltout => \U400_SDRAM.N_258_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_0_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110011"
        )
    port map (
            in0 => \N__4910\,
            in1 => \N__3131\,
            in2 => \N__3125\,
            in3 => \N__3122\,
            lcout => \U400_SDRAM.N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNISAQQ4_1_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__4795\,
            in1 => \N__5039\,
            in2 => \_gnd_net_\,
            in3 => \N__5395\,
            lcout => \U400_SDRAM.N_240\,
            ltout => \U400_SDRAM.N_240_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3982\,
            in2 => \N__3110\,
            in3 => \N__5001\,
            lcout => \U400_SDRAM.N_219_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNIMIPA1_1_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3107\,
            in1 => \N__3091\,
            in2 => \N__3080\,
            in3 => \N__3063\,
            lcout => \U400_SDRAM.un1_REFRESH_COUNTERlto7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_1_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3064\,
            in1 => \_gnd_net_\,
            in2 => \N__3007\,
            in3 => \_gnd_net_\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__2980\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNIUQPA1_5_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3049\,
            in1 => \N__3038\,
            in2 => \N__3023\,
            in3 => \N__2999\,
            lcout => \U400_SDRAM.un1_REFRESH_COUNTERlto7_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_0_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3000\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__2980\
        );

    \U400_SDRAM.CS0_EN_RNO_0_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__3181\,
            in1 => \N__3259\,
            in2 => \N__3169\,
            in3 => \N__3550\,
            lcout => OPEN,
            ltout => \U400_SDRAM.CS0_EN_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS0_EN_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__4798\,
            in1 => \N__5045\,
            in2 => \N__3185\,
            in3 => \N__5397\,
            lcout => \U400_SDRAM.CS0_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0_ENC_net\,
            ce => 'H',
            sr => \N__6160\
        );

    \U400_SDRAM.CS1_EN_RNO_0_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000101110"
        )
    port map (
            in0 => \N__3631\,
            in1 => \N__3260\,
            in2 => \N__3170\,
            in3 => \N__3551\,
            lcout => OPEN,
            ltout => \U400_SDRAM.CS1_EN_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS1_EN_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__4799\,
            in1 => \N__5046\,
            in2 => \N__3149\,
            in3 => \N__5398\,
            lcout => \U400_SDRAM.CS1_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0_ENC_net\,
            ce => 'H',
            sr => \N__6160\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_2_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4441\,
            in1 => \N__4925\,
            in2 => \N__4597\,
            in3 => \N__4331\,
            lcout => \U400_SDRAM.N_114\,
            ltout => \U400_SDRAM.N_114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000001000"
        )
    port map (
            in0 => \N__5527\,
            in1 => \N__4789\,
            in2 => \N__3146\,
            in3 => \N__4380\,
            lcout => \U400_SDRAM.N_242\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIVG1P5_2_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__3143\,
            in1 => \N__3941\,
            in2 => \_gnd_net_\,
            in3 => \N__3258\,
            lcout => \U400_SDRAM.N_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI4ECU1_2_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__4333\,
            in1 => \N__4468\,
            in2 => \N__3530\,
            in3 => \N__5520\,
            lcout => \U400_SDRAM.N_220\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIRRB91_0_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4930\,
            in1 => \N__4589\,
            in2 => \_gnd_net_\,
            in3 => \N__4335\,
            lcout => \U400_SDRAM.N_261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI7D8G1_0_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__4931\,
            in1 => \N__4588\,
            in2 => \N__4813\,
            in3 => \N__4332\,
            lcout => \U400_SDRAM.N_140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__4590\,
            in1 => \N__3421\,
            in2 => \_gnd_net_\,
            in3 => \N__5047\,
            lcout => \U400_SDRAM.N_207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3_0_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100110001"
        )
    port map (
            in0 => \N__4785\,
            in1 => \N__5391\,
            in2 => \N__5546\,
            in3 => \N__4381\,
            lcout => \U400_SDRAM.SDRAM_CONFIGURED_RNI5POA3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI36NC1_2_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101111"
        )
    port map (
            in0 => \N__4334\,
            in1 => \N__4469\,
            in2 => \N__4949\,
            in3 => \N__5521\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI2LE84_2_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__3952\,
            in1 => \N__3661\,
            in2 => \N__3248\,
            in3 => \N__3419\,
            lcout => \U400_SDRAM.N_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_9_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6502\,
            in1 => \N__6068\,
            in2 => \N__3245\,
            in3 => \N__5968\,
            lcout => \MA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_9C_net\,
            ce => \N__6267\,
            sr => \N__6164\
        );

    \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2_1_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__3218\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3212\,
            lcout => \U400_ADDRESS_DECODE_RAM_SPACE_i_o3_0_o2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.BURST_RNISKH51_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4217\,
            in1 => \N__4106\,
            in2 => \N__4256\,
            in3 => \N__3738\,
            lcout => \U400_SDRAM.TA_COUNTER_0_sqmuxa\,
            ltout => \U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__4171\,
            in1 => \N__3706\,
            in2 => \N__3200\,
            in3 => \N__4146\,
            lcout => \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_EN_i_ess_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__4147\,
            in1 => \N__3983\,
            in2 => \_gnd_net_\,
            in3 => \N__4172\,
            lcout => \TA_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4070\,
            ce => \N__3191\,
            sr => \N__6171\
        );

    \U400_SDRAM.BANK0_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__3367\,
            in1 => \N__3340\,
            in2 => \N__3398\,
            in3 => \N__5002\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK0C_net\,
            ce => 'H',
            sr => \N__6165\
        );

    \U400_SDRAM.BANK1_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__5003\,
            in1 => \N__3316\,
            in2 => \N__3356\,
            in3 => \N__3341\,
            lcout => \BANK1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK0C_net\,
            ce => 'H',
            sr => \N__6165\
        );

    \U400_SDRAM.RAM_CYCLE_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__3272\,
            in1 => \N__3572\,
            in2 => \N__3981\,
            in3 => \N__5150\,
            lcout => \U400_SDRAM.RAM_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK0C_net\,
            ce => 'H',
            sr => \N__6165\
        );

    \U400_SDRAM.WRITE_CYCLE_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__3570\,
            in1 => \N__3305\,
            in2 => \_gnd_net_\,
            in3 => \N__4671\,
            lcout => \U400_SDRAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK0C_net\,
            ce => 'H',
            sr => \N__6165\
        );

    \U400_SDRAM.TACK_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__3293\,
            in1 => \N__3287\,
            in2 => \_gnd_net_\,
            in3 => \N__4151\,
            lcout => \U400_SDRAM.TACKZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK0C_net\,
            ce => 'H',
            sr => \N__6165\
        );

    \U400_SDRAM.BURST_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__5757\,
            in1 => \N__3571\,
            in2 => \N__3743\,
            in3 => \N__5824\,
            lcout => \U400_SDRAM.BURSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK0C_net\,
            ce => 'H',
            sr => \N__6165\
        );

    \U400_SDRAM.BURST8_i_0_i_i_o2_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5756\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5823\,
            lcout => \U400_SDRAM.N_118\,
            ltout => \U400_SDRAM.N_118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5394\,
            in1 => \N__5043\,
            in2 => \N__3281\,
            in3 => \N__4998\,
            lcout => \U400_SDRAM.N_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__4999\,
            in1 => \N__5054\,
            in2 => \N__3966\,
            in3 => \N__3271\,
            lcout => \U400_SDRAM.RAM_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4067\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_RNO_3_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110101010"
        )
    port map (
            in0 => \N__4774\,
            in1 => \N__4587\,
            in2 => \_gnd_net_\,
            in3 => \N__4901\,
            lcout => \U400_SDRAM.N_189\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNI8BL33_8_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__3799\,
            in1 => \N__3829\,
            in2 => \N__5544\,
            in3 => \N__3814\,
            lcout => \U400_SDRAM.N_236\,
            ltout => \U400_SDRAM.N_236_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNI58I35_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5393\,
            in1 => \N__4794\,
            in2 => \N__3575\,
            in3 => \N__4996\,
            lcout => \U400_SDRAM.N_23_i\,
            ltout => \U400_SDRAM.N_23_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNIRHEJ5_0_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__3940\,
            in1 => \_gnd_net_\,
            in2 => \N__3560\,
            in3 => \_gnd_net_\,
            lcout => \U400_SDRAM.N_259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNIUFE78_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__5392\,
            in1 => \N__3557\,
            in2 => \N__5048\,
            in3 => \N__4997\,
            lcout => \U400_SDRAM.N_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_1_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__3542\,
            in1 => \N__3492\,
            in2 => \N__3512\,
            in3 => \N__3520\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_1C_net\,
            ce => \N__3446\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001100110"
        )
    port map (
            in0 => \N__4773\,
            in1 => \N__4574\,
            in2 => \N__4687\,
            in3 => \N__4940\,
            lcout => \U400_SDRAM.N_198\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_3_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__3521\,
            in1 => \N__3511\,
            in2 => \N__3500\,
            in3 => \N__3458\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_1C_net\,
            ce => \N__3446\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__3428\,
            in1 => \N__4826\,
            in2 => \N__3677\,
            in3 => \N__3641\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_1_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101010"
        )
    port map (
            in0 => \N__6040\,
            in1 => \N__3689\,
            in2 => \N__3680\,
            in3 => \N__5349\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5549\,
            in1 => \N__4592\,
            in2 => \_gnd_net_\,
            in3 => \N__4946\,
            lcout => \U400_SDRAM.N_250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111101010"
        )
    port map (
            in0 => \N__4947\,
            in1 => \N__5550\,
            in2 => \N__4615\,
            in3 => \N__4492\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_31_i_i_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__3650\,
            in1 => \N__3932\,
            in2 => \N__3668\,
            in3 => \N__5552\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_31_i_i_i_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_2_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__6425\,
            in1 => \N__5350\,
            in2 => \N__3665\,
            in3 => \N__4961\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_ne_RNO_0_0_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101011111111"
        )
    port map (
            in0 => \N__3662\,
            in1 => \N__4796\,
            in2 => \N__4688\,
            in3 => \N__3936\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001111"
        )
    port map (
            in0 => \N__5551\,
            in1 => \N__3649\,
            in2 => \N__3965\,
            in3 => \N__4393\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS1n_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__6426\,
            in1 => \N__6031\,
            in2 => \N__3635\,
            in3 => \N__5924\,
            lcout => \CS1n_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS1nC_net\,
            ce => 'H',
            sr => \N__6161\
        );

    \U400_SDRAM.MA_nesr_12_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6462\,
            in1 => \N__6074\,
            in2 => \N__3605\,
            in3 => \N__5960\,
            lcout => \MA_c_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_12C_net\,
            ce => \N__6258\,
            sr => \N__6170\
        );

    \U400_SDRAM.TA_OUT_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__4288\,
            in1 => \N__3713\,
            in2 => \N__3769\,
            in3 => \N__3722\,
            lcout => \TA_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4074\,
            ce => 'H',
            sr => \N__6173\
        );

    \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4279\,
            in1 => \N__4213\,
            in2 => \N__4255\,
            in3 => \N__4102\,
            lcout => \U400_SDRAM.TA_COUNTER27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_UUBEn_i_0_0_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__5857\,
            in1 => \N__5246\,
            in2 => \N__5195\,
            in3 => \N__5267\,
            lcout => \N_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4278\,
            in1 => \N__4212\,
            in2 => \N__4254\,
            in3 => \N__4103\,
            lcout => \U400_SDRAM.TA_COUNTER23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_OUT_RNO_0_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4105\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3739\,
            lcout => \U400_SDRAM.TA_EN11_m\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_OUT_RNO_2_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__4104\,
            in1 => \N__4249\,
            in2 => \N__4222\,
            in3 => \N__4280\,
            lcout => OPEN,
            ltout => \U400_SDRAM.un1_TA_COUNTER26_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_OUT_RNO_1_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4177\,
            in2 => \N__3716\,
            in3 => \N__4148\,
            lcout => \U400_SDRAM.un1_TA_COUNTER26_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_1_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__4109\,
            in1 => \N__3968\,
            in2 => \N__4223\,
            in3 => \N__3695\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNI0LUG4_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__4149\,
            in1 => \N__3707\,
            in2 => \N__4178\,
            in3 => \N__4117\,
            lcout => \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0\,
            ltout => \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_2_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__4284\,
            in1 => \N__4189\,
            in2 => \N__4292\,
            in3 => \N__3969\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_3_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110010000000"
        )
    port map (
            in0 => \N__4190\,
            in1 => \N__3970\,
            in2 => \N__4289\,
            in3 => \N__4253\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4218\,
            in2 => \_gnd_net_\,
            in3 => \N__4107\,
            lcout => \U400_SDRAM.CO1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__4108\,
            in1 => \N__4173\,
            in2 => \_gnd_net_\,
            in3 => \N__4150\,
            lcout => OPEN,
            ltout => \U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_0_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__3967\,
            in1 => \_gnd_net_\,
            in2 => \N__4121\,
            in3 => \N__4118\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4071\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_RNO_2_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__3989\,
            in1 => \N__4473\,
            in2 => \N__5545\,
            in3 => \N__4357\,
            lcout => \U400_SDRAM.un1_SDRAM_COUNTER52_2_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.RAM_SPACE_i_o3_0_o2dup_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__5083\,
            in1 => \N__5120\,
            in2 => \N__5144\,
            in3 => \N__3942\,
            lcout => \RAM_SPACE_i_o3_0_o2dup\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_RNO_1_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__3833\,
            in1 => \N__3818\,
            in2 => \N__3803\,
            in3 => \N__4995\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_195_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_RNO_0_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__5159\,
            in1 => \N__4596\,
            in2 => \N__5153\,
            in3 => \N__4948\,
            lcout => \U400_SDRAM.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5143\,
            in1 => \N__5116\,
            in2 => \N__5090\,
            in3 => \N__5063\,
            lcout => \U400_SDRAM.N_225\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__4491\,
            in1 => \N__5044\,
            in2 => \_gnd_net_\,
            in3 => \N__5000\,
            lcout => \U400_SDRAM.N_228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_6_1_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4790\,
            in1 => \N__4572\,
            in2 => \_gnd_net_\,
            in3 => \N__4941\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_a2_2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_5_1_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110000"
        )
    port map (
            in0 => \N__4573\,
            in1 => \N__5528\,
            in2 => \N__4955\,
            in3 => \N__4489\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111111010"
        )
    port map (
            in0 => \N__4490\,
            in1 => \N__5529\,
            in2 => \N__4952\,
            in3 => \N__4942\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_ne_RNO_2_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__4797\,
            in1 => \N__4680\,
            in2 => \N__5548\,
            in3 => \N__4591\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_a2_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_ne_RNO_1_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__4493\,
            in1 => \N__4394\,
            in2 => \N__4364\,
            in3 => \N__4361\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_ne_0_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__5533\,
            in1 => \N__5414\,
            in2 => \N__5408\,
            in3 => \N__5405\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_ne_0C_net\,
            ce => \N__5354\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_11_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6485\,
            in1 => \N__6075\,
            in2 => \N__5336\,
            in3 => \N__5959\,
            lcout => \MA_c_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_11C_net\,
            ce => \N__6254\,
            sr => \N__6172\
        );

    \U400_SDRAM.MA_nesr_RNO_0_5_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001110"
        )
    port map (
            in0 => \N__6499\,
            in1 => \N__6070\,
            in2 => \N__5312\,
            in3 => \N__5958\,
            lcout => \U400_SDRAM.MA_5_iv_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_5_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__5300\,
            in1 => \N__5288\,
            in2 => \_gnd_net_\,
            in3 => \N__6337\,
            lcout => \MA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_5C_net\,
            ce => \N__6265\,
            sr => \N__6178\
        );

    \U400_BYTE_ENABLE.un1_UUBEn_i_0_0_x2_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5822\,
            in2 => \_gnd_net_\,
            in3 => \N__5755\,
            lcout => \U400_BYTE_ENABLE.N_101_i\,
            ltout => \U400_BYTE_ENABLE.N_101_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_LMBEn_i_0_0_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010000"
        )
    port map (
            in0 => \N__5853\,
            in1 => \N__5245\,
            in2 => \N__5261\,
            in3 => \N__5193\,
            lcout => \un1_LMBEn_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_UMBEn_i_0_0_o2_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__5759\,
            in1 => \N__5238\,
            in2 => \N__5825\,
            in3 => \N__5183\,
            lcout => \U400_BYTE_ENABLE.N_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_ne_RNIIMNC_0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6474\,
            in1 => \N__6062\,
            in2 => \_gnd_net_\,
            in3 => \N__5954\,
            lcout => \U400_SDRAM.MA19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_ne_RNI80KS_0_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011110111"
        )
    port map (
            in0 => \N__6475\,
            in1 => \N__6063\,
            in2 => \N__6191\,
            in3 => \N__5955\,
            lcout => \U400_SDRAM.un1_MA20_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_10_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001000100"
        )
    port map (
            in0 => \N__6501\,
            in1 => \N__6076\,
            in2 => \N__6110\,
            in3 => \N__5956\,
            lcout => \MA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_10C_net\,
            ce => \N__6237\,
            sr => \N__6177\
        );

    \U400_SDRAM.MA_nesr_RNO_0_1_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001110"
        )
    port map (
            in0 => \N__6500\,
            in1 => \N__6077\,
            in2 => \N__5984\,
            in3 => \N__5957\,
            lcout => \U400_SDRAM.MA_5_iv_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_UMBEn_i_0_0_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001000"
        )
    port map (
            in0 => \N__5812\,
            in1 => \N__5867\,
            in2 => \N__5758\,
            in3 => \N__5770\,
            lcout => \N_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_LLBEn_i_0_0_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110100"
        )
    port map (
            in0 => \N__5866\,
            in1 => \N__5811\,
            in2 => \N__5771\,
            in3 => \N__5748\,
            lcout => \un1_LLBEn_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TAn_obuft_RNO_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5684\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_526_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_3_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__5663\,
            in1 => \N__6495\,
            in2 => \N__5654\,
            in3 => \N__6310\,
            lcout => \MA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_3C_net\,
            ce => \N__6241\,
            sr => \N__6179\
        );

    \U400_SDRAM.MA_nesr_2_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__6335\,
            in1 => \N__5621\,
            in2 => \N__5609\,
            in3 => \N__6497\,
            lcout => \MA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_2C_net\,
            ce => \N__6266\,
            sr => \N__6180\
        );

    \U400_SDRAM.MA_nesr_0_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__5588\,
            in1 => \N__6496\,
            in2 => \N__5576\,
            in3 => \N__6334\,
            lcout => \MA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_2C_net\,
            ce => \N__6266\,
            sr => \N__6180\
        );

    \U400_SDRAM.MA_nesr_4_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__6336\,
            in1 => \N__6530\,
            in2 => \N__6518\,
            in3 => \N__6498\,
            lcout => \MA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_2C_net\,
            ce => \N__6266\,
            sr => \N__6180\
        );

    \U400_SDRAM.MA_nesr_1_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__6353\,
            in1 => \N__6347\,
            in2 => \_gnd_net_\,
            in3 => \N__6333\,
            lcout => \MA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_2C_net\,
            ce => \N__6266\,
            sr => \N__6180\
        );
end \INTERFACE\;

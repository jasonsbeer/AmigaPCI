// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Feb 8 2025 11:10:31

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    DRA,
    CMA,
    A,
    RAMENn,
    TSn,
    DMA_LATCH,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    LDSn,
    LATCH_CLK,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    DBRn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    input [9:0] DRA;
    output [10:0] CMA;
    input [20:0] A;
    output RAMENn;
    input TSn;
    output DMA_LATCH;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    input DBRn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__11113;
    wire N__11112;
    wire N__11111;
    wire N__11104;
    wire N__11103;
    wire N__11102;
    wire N__11095;
    wire N__11094;
    wire N__11093;
    wire N__11086;
    wire N__11085;
    wire N__11084;
    wire N__11077;
    wire N__11076;
    wire N__11075;
    wire N__11068;
    wire N__11067;
    wire N__11066;
    wire N__11059;
    wire N__11058;
    wire N__11057;
    wire N__11050;
    wire N__11049;
    wire N__11048;
    wire N__11041;
    wire N__11040;
    wire N__11039;
    wire N__11032;
    wire N__11031;
    wire N__11030;
    wire N__11023;
    wire N__11022;
    wire N__11021;
    wire N__11014;
    wire N__11013;
    wire N__11012;
    wire N__11005;
    wire N__11004;
    wire N__11003;
    wire N__10996;
    wire N__10995;
    wire N__10994;
    wire N__10987;
    wire N__10986;
    wire N__10985;
    wire N__10978;
    wire N__10977;
    wire N__10976;
    wire N__10969;
    wire N__10968;
    wire N__10967;
    wire N__10960;
    wire N__10959;
    wire N__10958;
    wire N__10951;
    wire N__10950;
    wire N__10949;
    wire N__10942;
    wire N__10941;
    wire N__10940;
    wire N__10933;
    wire N__10932;
    wire N__10931;
    wire N__10924;
    wire N__10923;
    wire N__10922;
    wire N__10915;
    wire N__10914;
    wire N__10913;
    wire N__10906;
    wire N__10905;
    wire N__10904;
    wire N__10897;
    wire N__10896;
    wire N__10895;
    wire N__10888;
    wire N__10887;
    wire N__10886;
    wire N__10879;
    wire N__10878;
    wire N__10877;
    wire N__10870;
    wire N__10869;
    wire N__10868;
    wire N__10861;
    wire N__10860;
    wire N__10859;
    wire N__10852;
    wire N__10851;
    wire N__10850;
    wire N__10843;
    wire N__10842;
    wire N__10841;
    wire N__10834;
    wire N__10833;
    wire N__10832;
    wire N__10825;
    wire N__10824;
    wire N__10823;
    wire N__10816;
    wire N__10815;
    wire N__10814;
    wire N__10807;
    wire N__10806;
    wire N__10805;
    wire N__10798;
    wire N__10797;
    wire N__10796;
    wire N__10789;
    wire N__10788;
    wire N__10787;
    wire N__10780;
    wire N__10779;
    wire N__10778;
    wire N__10771;
    wire N__10770;
    wire N__10769;
    wire N__10762;
    wire N__10761;
    wire N__10760;
    wire N__10753;
    wire N__10752;
    wire N__10751;
    wire N__10744;
    wire N__10743;
    wire N__10742;
    wire N__10735;
    wire N__10734;
    wire N__10733;
    wire N__10726;
    wire N__10725;
    wire N__10724;
    wire N__10717;
    wire N__10716;
    wire N__10715;
    wire N__10708;
    wire N__10707;
    wire N__10706;
    wire N__10699;
    wire N__10698;
    wire N__10697;
    wire N__10690;
    wire N__10689;
    wire N__10688;
    wire N__10681;
    wire N__10680;
    wire N__10679;
    wire N__10672;
    wire N__10671;
    wire N__10670;
    wire N__10663;
    wire N__10662;
    wire N__10661;
    wire N__10654;
    wire N__10653;
    wire N__10652;
    wire N__10645;
    wire N__10644;
    wire N__10643;
    wire N__10636;
    wire N__10635;
    wire N__10634;
    wire N__10627;
    wire N__10626;
    wire N__10625;
    wire N__10618;
    wire N__10617;
    wire N__10616;
    wire N__10609;
    wire N__10608;
    wire N__10607;
    wire N__10600;
    wire N__10599;
    wire N__10598;
    wire N__10591;
    wire N__10590;
    wire N__10589;
    wire N__10582;
    wire N__10581;
    wire N__10580;
    wire N__10573;
    wire N__10572;
    wire N__10571;
    wire N__10564;
    wire N__10563;
    wire N__10562;
    wire N__10555;
    wire N__10554;
    wire N__10553;
    wire N__10546;
    wire N__10545;
    wire N__10544;
    wire N__10537;
    wire N__10536;
    wire N__10535;
    wire N__10528;
    wire N__10527;
    wire N__10526;
    wire N__10519;
    wire N__10518;
    wire N__10517;
    wire N__10510;
    wire N__10509;
    wire N__10508;
    wire N__10501;
    wire N__10500;
    wire N__10499;
    wire N__10492;
    wire N__10491;
    wire N__10490;
    wire N__10483;
    wire N__10482;
    wire N__10481;
    wire N__10474;
    wire N__10473;
    wire N__10472;
    wire N__10465;
    wire N__10464;
    wire N__10463;
    wire N__10456;
    wire N__10455;
    wire N__10454;
    wire N__10447;
    wire N__10446;
    wire N__10445;
    wire N__10438;
    wire N__10437;
    wire N__10436;
    wire N__10429;
    wire N__10428;
    wire N__10427;
    wire N__10420;
    wire N__10419;
    wire N__10418;
    wire N__10411;
    wire N__10410;
    wire N__10409;
    wire N__10402;
    wire N__10401;
    wire N__10400;
    wire N__10393;
    wire N__10392;
    wire N__10391;
    wire N__10384;
    wire N__10383;
    wire N__10382;
    wire N__10375;
    wire N__10374;
    wire N__10373;
    wire N__10366;
    wire N__10365;
    wire N__10364;
    wire N__10357;
    wire N__10356;
    wire N__10355;
    wire N__10348;
    wire N__10347;
    wire N__10346;
    wire N__10339;
    wire N__10338;
    wire N__10337;
    wire N__10320;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10308;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10296;
    wire N__10293;
    wire N__10292;
    wire N__10291;
    wire N__10288;
    wire N__10287;
    wire N__10286;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10254;
    wire N__10249;
    wire N__10246;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10232;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10222;
    wire N__10217;
    wire N__10216;
    wire N__10211;
    wire N__10208;
    wire N__10207;
    wire N__10204;
    wire N__10201;
    wire N__10200;
    wire N__10197;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10170;
    wire N__10165;
    wire N__10162;
    wire N__10157;
    wire N__10152;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10139;
    wire N__10138;
    wire N__10137;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10120;
    wire N__10119;
    wire N__10118;
    wire N__10117;
    wire N__10116;
    wire N__10115;
    wire N__10112;
    wire N__10111;
    wire N__10110;
    wire N__10109;
    wire N__10108;
    wire N__10105;
    wire N__10102;
    wire N__10101;
    wire N__10100;
    wire N__10099;
    wire N__10098;
    wire N__10097;
    wire N__10096;
    wire N__10095;
    wire N__10094;
    wire N__10093;
    wire N__10092;
    wire N__10091;
    wire N__10090;
    wire N__10089;
    wire N__10088;
    wire N__10087;
    wire N__10086;
    wire N__10085;
    wire N__10084;
    wire N__10083;
    wire N__10082;
    wire N__10081;
    wire N__10080;
    wire N__10079;
    wire N__10078;
    wire N__10075;
    wire N__10072;
    wire N__9993;
    wire N__9990;
    wire N__9987;
    wire N__9986;
    wire N__9983;
    wire N__9982;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9954;
    wire N__9951;
    wire N__9948;
    wire N__9945;
    wire N__9942;
    wire N__9939;
    wire N__9936;
    wire N__9933;
    wire N__9930;
    wire N__9927;
    wire N__9924;
    wire N__9921;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9909;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9882;
    wire N__9879;
    wire N__9878;
    wire N__9877;
    wire N__9876;
    wire N__9875;
    wire N__9872;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9860;
    wire N__9855;
    wire N__9852;
    wire N__9849;
    wire N__9846;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9774;
    wire N__9771;
    wire N__9770;
    wire N__9767;
    wire N__9766;
    wire N__9763;
    wire N__9762;
    wire N__9759;
    wire N__9756;
    wire N__9751;
    wire N__9748;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9732;
    wire N__9729;
    wire N__9726;
    wire N__9725;
    wire N__9724;
    wire N__9723;
    wire N__9722;
    wire N__9719;
    wire N__9718;
    wire N__9713;
    wire N__9710;
    wire N__9709;
    wire N__9706;
    wire N__9705;
    wire N__9702;
    wire N__9699;
    wire N__9698;
    wire N__9697;
    wire N__9696;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9688;
    wire N__9685;
    wire N__9684;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9664;
    wire N__9661;
    wire N__9660;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9648;
    wire N__9647;
    wire N__9646;
    wire N__9643;
    wire N__9642;
    wire N__9641;
    wire N__9640;
    wire N__9639;
    wire N__9636;
    wire N__9631;
    wire N__9622;
    wire N__9621;
    wire N__9620;
    wire N__9619;
    wire N__9616;
    wire N__9615;
    wire N__9610;
    wire N__9607;
    wire N__9602;
    wire N__9599;
    wire N__9594;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9578;
    wire N__9573;
    wire N__9570;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9550;
    wire N__9543;
    wire N__9528;
    wire N__9525;
    wire N__9524;
    wire N__9523;
    wire N__9522;
    wire N__9519;
    wire N__9518;
    wire N__9515;
    wire N__9514;
    wire N__9513;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9495;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9477;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9450;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9442;
    wire N__9439;
    wire N__9436;
    wire N__9433;
    wire N__9430;
    wire N__9427;
    wire N__9424;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9399;
    wire N__9396;
    wire N__9393;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9375;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9358;
    wire N__9355;
    wire N__9346;
    wire N__9343;
    wire N__9336;
    wire N__9333;
    wire N__9330;
    wire N__9329;
    wire N__9328;
    wire N__9325;
    wire N__9324;
    wire N__9319;
    wire N__9316;
    wire N__9313;
    wire N__9310;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9276;
    wire N__9273;
    wire N__9272;
    wire N__9271;
    wire N__9268;
    wire N__9263;
    wire N__9258;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9221;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9210;
    wire N__9207;
    wire N__9202;
    wire N__9199;
    wire N__9196;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9129;
    wire N__9126;
    wire N__9125;
    wire N__9124;
    wire N__9123;
    wire N__9122;
    wire N__9121;
    wire N__9120;
    wire N__9119;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9111;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9101;
    wire N__9100;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9092;
    wire N__9089;
    wire N__9088;
    wire N__9085;
    wire N__9084;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9076;
    wire N__9063;
    wire N__9060;
    wire N__9045;
    wire N__9042;
    wire N__9041;
    wire N__9040;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9018;
    wire N__9015;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9003;
    wire N__9000;
    wire N__8995;
    wire N__8992;
    wire N__8983;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8961;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8947;
    wire N__8946;
    wire N__8941;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8927;
    wire N__8922;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8898;
    wire N__8897;
    wire N__8896;
    wire N__8895;
    wire N__8894;
    wire N__8893;
    wire N__8890;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8870;
    wire N__8867;
    wire N__8866;
    wire N__8863;
    wire N__8860;
    wire N__8857;
    wire N__8856;
    wire N__8849;
    wire N__8846;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8814;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8787;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8772;
    wire N__8769;
    wire N__8766;
    wire N__8763;
    wire N__8760;
    wire N__8757;
    wire N__8754;
    wire N__8751;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8732;
    wire N__8731;
    wire N__8730;
    wire N__8729;
    wire N__8728;
    wire N__8727;
    wire N__8726;
    wire N__8725;
    wire N__8724;
    wire N__8723;
    wire N__8722;
    wire N__8721;
    wire N__8720;
    wire N__8719;
    wire N__8718;
    wire N__8717;
    wire N__8716;
    wire N__8715;
    wire N__8714;
    wire N__8713;
    wire N__8712;
    wire N__8711;
    wire N__8710;
    wire N__8707;
    wire N__8706;
    wire N__8705;
    wire N__8704;
    wire N__8703;
    wire N__8702;
    wire N__8701;
    wire N__8700;
    wire N__8699;
    wire N__8698;
    wire N__8697;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8619;
    wire N__8616;
    wire N__8613;
    wire N__8610;
    wire N__8609;
    wire N__8608;
    wire N__8607;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8589;
    wire N__8586;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8574;
    wire N__8571;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8561;
    wire N__8558;
    wire N__8557;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8538;
    wire N__8535;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8523;
    wire N__8520;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8503;
    wire N__8500;
    wire N__8497;
    wire N__8494;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8463;
    wire N__8462;
    wire N__8461;
    wire N__8460;
    wire N__8459;
    wire N__8458;
    wire N__8457;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8431;
    wire N__8430;
    wire N__8427;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8407;
    wire N__8406;
    wire N__8405;
    wire N__8404;
    wire N__8403;
    wire N__8400;
    wire N__8399;
    wire N__8398;
    wire N__8397;
    wire N__8396;
    wire N__8393;
    wire N__8386;
    wire N__8379;
    wire N__8370;
    wire N__8369;
    wire N__8368;
    wire N__8365;
    wire N__8364;
    wire N__8361;
    wire N__8360;
    wire N__8357;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8328;
    wire N__8325;
    wire N__8320;
    wire N__8317;
    wire N__8298;
    wire N__8295;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8272;
    wire N__8271;
    wire N__8270;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8256;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8244;
    wire N__8241;
    wire N__8238;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8220;
    wire N__8217;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire N__8207;
    wire N__8206;
    wire N__8205;
    wire N__8202;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8184;
    wire N__8181;
    wire N__8178;
    wire N__8175;
    wire N__8172;
    wire N__8169;
    wire N__8168;
    wire N__8167;
    wire N__8166;
    wire N__8163;
    wire N__8160;
    wire N__8157;
    wire N__8154;
    wire N__8147;
    wire N__8142;
    wire N__8139;
    wire N__8136;
    wire N__8133;
    wire N__8132;
    wire N__8127;
    wire N__8124;
    wire N__8121;
    wire N__8118;
    wire N__8115;
    wire N__8112;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8094;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8082;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8066;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8040;
    wire N__8037;
    wire N__8034;
    wire N__8031;
    wire N__8028;
    wire N__8027;
    wire N__8022;
    wire N__8021;
    wire N__8020;
    wire N__8017;
    wire N__8012;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7982;
    wire N__7981;
    wire N__7980;
    wire N__7975;
    wire N__7970;
    wire N__7965;
    wire N__7962;
    wire N__7959;
    wire N__7956;
    wire N__7953;
    wire N__7950;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7917;
    wire N__7914;
    wire N__7913;
    wire N__7912;
    wire N__7909;
    wire N__7908;
    wire N__7905;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7881;
    wire N__7878;
    wire N__7875;
    wire N__7872;
    wire N__7871;
    wire N__7870;
    wire N__7867;
    wire N__7864;
    wire N__7861;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7849;
    wire N__7846;
    wire N__7843;
    wire N__7840;
    wire N__7837;
    wire N__7834;
    wire N__7831;
    wire N__7828;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7812;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7804;
    wire N__7801;
    wire N__7798;
    wire N__7795;
    wire N__7790;
    wire N__7789;
    wire N__7786;
    wire N__7783;
    wire N__7780;
    wire N__7777;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7749;
    wire N__7748;
    wire N__7747;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7735;
    wire N__7734;
    wire N__7733;
    wire N__7732;
    wire N__7731;
    wire N__7730;
    wire N__7727;
    wire N__7724;
    wire N__7721;
    wire N__7704;
    wire N__7701;
    wire N__7698;
    wire N__7697;
    wire N__7696;
    wire N__7695;
    wire N__7694;
    wire N__7693;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7685;
    wire N__7682;
    wire N__7677;
    wire N__7672;
    wire N__7667;
    wire N__7664;
    wire N__7663;
    wire N__7662;
    wire N__7661;
    wire N__7658;
    wire N__7657;
    wire N__7654;
    wire N__7647;
    wire N__7644;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7632;
    wire N__7629;
    wire N__7624;
    wire N__7621;
    wire N__7618;
    wire N__7617;
    wire N__7616;
    wire N__7615;
    wire N__7614;
    wire N__7613;
    wire N__7612;
    wire N__7607;
    wire N__7602;
    wire N__7597;
    wire N__7588;
    wire N__7583;
    wire N__7578;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7551;
    wire N__7550;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7533;
    wire N__7532;
    wire N__7531;
    wire N__7530;
    wire N__7527;
    wire N__7522;
    wire N__7517;
    wire N__7514;
    wire N__7511;
    wire N__7500;
    wire N__7497;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7485;
    wire N__7482;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7468;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7456;
    wire N__7449;
    wire N__7446;
    wire N__7443;
    wire N__7440;
    wire N__7437;
    wire N__7434;
    wire N__7431;
    wire N__7428;
    wire N__7425;
    wire N__7422;
    wire N__7419;
    wire N__7416;
    wire N__7413;
    wire N__7410;
    wire N__7407;
    wire N__7404;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7396;
    wire N__7391;
    wire N__7388;
    wire N__7387;
    wire N__7386;
    wire N__7385;
    wire N__7382;
    wire N__7379;
    wire N__7376;
    wire N__7373;
    wire N__7370;
    wire N__7359;
    wire N__7358;
    wire N__7357;
    wire N__7356;
    wire N__7353;
    wire N__7350;
    wire N__7349;
    wire N__7348;
    wire N__7347;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7322;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7306;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7281;
    wire N__7278;
    wire N__7275;
    wire N__7272;
    wire N__7269;
    wire N__7266;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7254;
    wire N__7251;
    wire N__7248;
    wire N__7245;
    wire N__7242;
    wire N__7239;
    wire N__7236;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7206;
    wire N__7205;
    wire N__7204;
    wire N__7203;
    wire N__7196;
    wire N__7193;
    wire N__7192;
    wire N__7191;
    wire N__7188;
    wire N__7185;
    wire N__7180;
    wire N__7173;
    wire N__7170;
    wire N__7167;
    wire N__7164;
    wire N__7161;
    wire N__7158;
    wire N__7155;
    wire N__7152;
    wire N__7149;
    wire N__7146;
    wire N__7143;
    wire N__7140;
    wire N__7137;
    wire N__7134;
    wire N__7133;
    wire N__7130;
    wire N__7127;
    wire N__7124;
    wire N__7119;
    wire N__7116;
    wire N__7113;
    wire N__7110;
    wire N__7107;
    wire N__7104;
    wire N__7101;
    wire N__7098;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7086;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7035;
    wire N__7032;
    wire N__7029;
    wire N__7026;
    wire N__7023;
    wire N__7020;
    wire N__7017;
    wire N__7014;
    wire N__7011;
    wire N__7008;
    wire N__7005;
    wire N__7002;
    wire N__6999;
    wire N__6996;
    wire N__6993;
    wire N__6990;
    wire N__6987;
    wire N__6984;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6957;
    wire N__6954;
    wire N__6951;
    wire N__6948;
    wire N__6945;
    wire N__6942;
    wire N__6939;
    wire N__6936;
    wire N__6933;
    wire N__6930;
    wire N__6927;
    wire N__6924;
    wire N__6921;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6882;
    wire N__6879;
    wire N__6876;
    wire N__6873;
    wire N__6870;
    wire N__6867;
    wire N__6864;
    wire N__6861;
    wire N__6858;
    wire N__6855;
    wire N__6852;
    wire N__6849;
    wire N__6846;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6819;
    wire N__6816;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6804;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6780;
    wire N__6777;
    wire N__6774;
    wire N__6771;
    wire N__6768;
    wire N__6767;
    wire N__6762;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6737;
    wire N__6736;
    wire N__6733;
    wire N__6728;
    wire N__6725;
    wire N__6720;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6710;
    wire N__6705;
    wire N__6702;
    wire N__6699;
    wire N__6696;
    wire N__6695;
    wire N__6694;
    wire N__6693;
    wire N__6692;
    wire N__6691;
    wire N__6690;
    wire N__6687;
    wire N__6680;
    wire N__6677;
    wire N__6672;
    wire N__6663;
    wire N__6662;
    wire N__6659;
    wire N__6658;
    wire N__6657;
    wire N__6654;
    wire N__6653;
    wire N__6648;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6636;
    wire N__6627;
    wire N__6626;
    wire N__6625;
    wire N__6624;
    wire N__6623;
    wire N__6622;
    wire N__6619;
    wire N__6616;
    wire N__6613;
    wire N__6608;
    wire N__6605;
    wire N__6600;
    wire N__6591;
    wire N__6590;
    wire N__6589;
    wire N__6588;
    wire N__6587;
    wire N__6586;
    wire N__6585;
    wire N__6584;
    wire N__6581;
    wire N__6576;
    wire N__6573;
    wire N__6564;
    wire N__6555;
    wire N__6554;
    wire N__6551;
    wire N__6550;
    wire N__6549;
    wire N__6548;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6536;
    wire N__6531;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6497;
    wire N__6494;
    wire N__6491;
    wire N__6486;
    wire N__6483;
    wire N__6480;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6468;
    wire N__6465;
    wire N__6464;
    wire N__6461;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6420;
    wire N__6417;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6375;
    wire N__6372;
    wire N__6371;
    wire N__6370;
    wire N__6369;
    wire N__6368;
    wire N__6367;
    wire N__6366;
    wire N__6359;
    wire N__6356;
    wire N__6349;
    wire N__6342;
    wire N__6339;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6327;
    wire N__6324;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6297;
    wire N__6294;
    wire N__6291;
    wire N__6290;
    wire N__6289;
    wire N__6288;
    wire N__6285;
    wire N__6282;
    wire N__6277;
    wire N__6276;
    wire N__6271;
    wire N__6268;
    wire N__6265;
    wire N__6258;
    wire N__6257;
    wire N__6256;
    wire N__6253;
    wire N__6252;
    wire N__6251;
    wire N__6250;
    wire N__6243;
    wire N__6242;
    wire N__6241;
    wire N__6238;
    wire N__6233;
    wire N__6230;
    wire N__6227;
    wire N__6226;
    wire N__6221;
    wire N__6218;
    wire N__6215;
    wire N__6210;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6188;
    wire N__6185;
    wire N__6182;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6170;
    wire N__6169;
    wire N__6168;
    wire N__6165;
    wire N__6162;
    wire N__6157;
    wire N__6150;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6142;
    wire N__6137;
    wire N__6136;
    wire N__6135;
    wire N__6134;
    wire N__6133;
    wire N__6132;
    wire N__6129;
    wire N__6126;
    wire N__6123;
    wire N__6122;
    wire N__6119;
    wire N__6118;
    wire N__6117;
    wire N__6114;
    wire N__6111;
    wire N__6110;
    wire N__6109;
    wire N__6108;
    wire N__6107;
    wire N__6106;
    wire N__6103;
    wire N__6096;
    wire N__6095;
    wire N__6092;
    wire N__6091;
    wire N__6090;
    wire N__6087;
    wire N__6084;
    wire N__6083;
    wire N__6078;
    wire N__6075;
    wire N__6070;
    wire N__6063;
    wire N__6060;
    wire N__6057;
    wire N__6048;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6030;
    wire N__6015;
    wire N__6014;
    wire N__6013;
    wire N__6012;
    wire N__6011;
    wire N__6008;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__6000;
    wire N__5999;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5981;
    wire N__5980;
    wire N__5979;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5971;
    wire N__5970;
    wire N__5963;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5951;
    wire N__5948;
    wire N__5941;
    wire N__5936;
    wire N__5933;
    wire N__5916;
    wire N__5915;
    wire N__5914;
    wire N__5913;
    wire N__5908;
    wire N__5907;
    wire N__5906;
    wire N__5905;
    wire N__5904;
    wire N__5903;
    wire N__5900;
    wire N__5899;
    wire N__5898;
    wire N__5895;
    wire N__5894;
    wire N__5891;
    wire N__5890;
    wire N__5887;
    wire N__5886;
    wire N__5883;
    wire N__5878;
    wire N__5873;
    wire N__5870;
    wire N__5869;
    wire N__5868;
    wire N__5865;
    wire N__5862;
    wire N__5859;
    wire N__5856;
    wire N__5849;
    wire N__5842;
    wire N__5835;
    wire N__5830;
    wire N__5817;
    wire N__5816;
    wire N__5815;
    wire N__5814;
    wire N__5813;
    wire N__5812;
    wire N__5811;
    wire N__5806;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5794;
    wire N__5793;
    wire N__5792;
    wire N__5791;
    wire N__5790;
    wire N__5789;
    wire N__5788;
    wire N__5787;
    wire N__5784;
    wire N__5783;
    wire N__5782;
    wire N__5781;
    wire N__5778;
    wire N__5775;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5758;
    wire N__5753;
    wire N__5748;
    wire N__5745;
    wire N__5738;
    wire N__5733;
    wire N__5730;
    wire N__5709;
    wire N__5706;
    wire N__5705;
    wire N__5702;
    wire N__5701;
    wire N__5700;
    wire N__5699;
    wire N__5698;
    wire N__5697;
    wire N__5696;
    wire N__5695;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5682;
    wire N__5677;
    wire N__5672;
    wire N__5671;
    wire N__5670;
    wire N__5669;
    wire N__5668;
    wire N__5667;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5655;
    wire N__5652;
    wire N__5645;
    wire N__5638;
    wire N__5633;
    wire N__5630;
    wire N__5613;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5598;
    wire N__5597;
    wire N__5596;
    wire N__5593;
    wire N__5588;
    wire N__5583;
    wire N__5582;
    wire N__5581;
    wire N__5580;
    wire N__5577;
    wire N__5570;
    wire N__5565;
    wire N__5562;
    wire N__5561;
    wire N__5560;
    wire N__5559;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5544;
    wire N__5535;
    wire N__5532;
    wire N__5529;
    wire N__5526;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5502;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5487;
    wire N__5484;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5472;
    wire N__5469;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5457;
    wire N__5454;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5432;
    wire N__5431;
    wire N__5426;
    wire N__5423;
    wire N__5418;
    wire N__5415;
    wire N__5414;
    wire N__5411;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5396;
    wire N__5391;
    wire N__5388;
    wire N__5387;
    wire N__5386;
    wire N__5383;
    wire N__5382;
    wire N__5379;
    wire N__5378;
    wire N__5377;
    wire N__5376;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5358;
    wire N__5355;
    wire N__5352;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5321;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5307;
    wire N__5304;
    wire N__5301;
    wire N__5298;
    wire N__5295;
    wire N__5292;
    wire N__5289;
    wire N__5286;
    wire N__5283;
    wire N__5280;
    wire N__5277;
    wire N__5274;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5262;
    wire N__5259;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5192;
    wire N__5191;
    wire N__5186;
    wire N__5183;
    wire N__5178;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5166;
    wire N__5163;
    wire N__5160;
    wire N__5157;
    wire N__5154;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5130;
    wire N__5127;
    wire N__5124;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5070;
    wire N__5069;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4977;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4965;
    wire N__4962;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4919;
    wire N__4918;
    wire N__4917;
    wire N__4916;
    wire N__4915;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4893;
    wire N__4888;
    wire N__4885;
    wire N__4882;
    wire N__4869;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4857;
    wire N__4856;
    wire N__4855;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4839;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4823;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4784;
    wire N__4783;
    wire N__4782;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4767;
    wire N__4766;
    wire N__4763;
    wire N__4756;
    wire N__4753;
    wire N__4746;
    wire N__4743;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4728;
    wire N__4725;
    wire N__4722;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4710;
    wire N__4707;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4695;
    wire N__4692;
    wire N__4689;
    wire N__4686;
    wire N__4683;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4647;
    wire N__4644;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4619;
    wire N__4618;
    wire N__4617;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4601;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4590;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4512;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4500;
    wire N__4499;
    wire N__4498;
    wire N__4497;
    wire N__4488;
    wire N__4485;
    wire N__4482;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4467;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4442;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4422;
    wire N__4419;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4395;
    wire N__4392;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4287;
    wire N__4284;
    wire N__4281;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4260;
    wire N__4257;
    wire N__4254;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4242;
    wire N__4241;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4221;
    wire N__4220;
    wire N__4217;
    wire N__4214;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4197;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4161;
    wire N__4158;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4122;
    wire N__4119;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4107;
    wire N__4104;
    wire N__4101;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4047;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4039;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3972;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3960;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3950;
    wire N__3945;
    wire N__3944;
    wire N__3941;
    wire N__3938;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3914;
    wire N__3911;
    wire N__3908;
    wire N__3903;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3891;
    wire N__3888;
    wire N__3887;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3875;
    wire N__3870;
    wire N__3867;
    wire N__3866;
    wire N__3865;
    wire N__3862;
    wire N__3857;
    wire N__3854;
    wire N__3849;
    wire N__3846;
    wire N__3843;
    wire N__3840;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3828;
    wire N__3825;
    wire N__3822;
    wire N__3819;
    wire N__3816;
    wire N__3813;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3795;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_PLL_i_i;
    wire N_1012_i;
    wire bfn_7_5_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire DBDIR_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_a3_0_0 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0_cascade_ ;
    wire \U712_CYCLE_TERM.N_223_i_0_en_cascade_ ;
    wire TACK_EN_i_ess;
    wire \U712_CYCLE_TERM.N_223_i_0_en_0 ;
    wire AWEn_c;
    wire N_242;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH5lto1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire \U712_CHIP_RAM.N_381_cascade_ ;
    wire VBENn_c;
    wire A_c_13;
    wire A_c_6;
    wire A_c_18;
    wire A_c_16;
    wire N_187_i;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_0_a3_0_cascade_ ;
    wire \U712_CHIP_RAM.N_273 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.N_328_cascade_ ;
    wire \U712_CHIP_RAM.N_332_cascade_ ;
    wire \U712_CHIP_RAM.A_m_2_20 ;
    wire A_c_20;
    wire \U712_CHIP_RAM.A_m_2_20_cascade_ ;
    wire \U712_CHIP_RAM.BANK0_esr_RNOZ0Z_1_cascade_ ;
    wire BANK0_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_10_0_0 ;
    wire \U712_CHIP_RAM.CPU_TACK_e_1 ;
    wire CPU_TACKm;
    wire TACK_OUTn;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CHIP_RAM.N_243 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire RAMENn_c;
    wire REG_TACK;
    wire \U712_REG_SM.N_225 ;
    wire \U712_REG_SM.N_225_cascade_ ;
    wire \U712_REG_SM.N_292 ;
    wire \U712_REG_SM.REG_TACK_RNOZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNT_srsts_i_i_0_3_cascade_ ;
    wire \U712_REG_SM.N_289 ;
    wire \U712_REG_SM.N_289_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire RnW_c;
    wire \U712_CHIP_RAM.N_261_cascade_ ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.N_260 ;
    wire \U712_CHIP_RAM.N_342_cascade_ ;
    wire \U712_CHIP_RAM.N_381 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_1_cascade_ ;
    wire A_c_8;
    wire A_c_15;
    wire \U712_CHIP_RAM.N_270_4 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_0_0_i_1 ;
    wire \U712_CHIP_RAM.N_211_cascade_ ;
    wire \U712_CHIP_RAM.N_87 ;
    wire \U712_CHIP_RAM.N_266 ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a3_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_264 ;
    wire \U712_CHIP_RAM.N_264_cascade_ ;
    wire \U712_CHIP_RAM.N_36_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_209 ;
    wire \U712_CHIP_RAM.N_209_cascade_ ;
    wire \U712_CHIP_RAM.N_263 ;
    wire \U712_CHIP_RAM.N_246 ;
    wire \U712_CHIP_RAM.N_332 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_203 ;
    wire \U712_CHIP_RAM.N_203_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_3_0 ;
    wire \U712_CHIP_RAM.N_341 ;
    wire \U712_CHIP_RAM.REFRESH_SYNCZ0Z_1 ;
    wire RAS1n_c;
    wire \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0 ;
    wire TSn_c;
    wire REGSPACEn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_2 ;
    wire DBR_SYNCZ0Z_1;
    wire DBR_SYNCZ0Z_0;
    wire \U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_1_2_cascade_ ;
    wire \U712_REG_SM.N_245 ;
    wire \U712_REG_SM.N_215 ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.N_215_cascade_ ;
    wire \U712_REG_SM.N_228_cascade_ ;
    wire \U712_REG_SM.STATE_COUNT_srsts_i_i_0_1_cascade_ ;
    wire C1_c;
    wire C3_c;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire A_c_5;
    wire A_c_12;
    wire A_c_7;
    wire \U712_CHIP_RAM.N_347_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_284 ;
    wire \U712_CHIP_RAM.N_211 ;
    wire \U712_CHIP_RAM.N_64_1 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_64_1_cascade_ ;
    wire \U712_CHIP_RAM.N_340 ;
    wire \U712_CHIP_RAM.N_340_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7 ;
    wire \U712_CHIP_RAM.N_267 ;
    wire \U712_CHIP_RAM.N_281_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_0_i_0 ;
    wire \U712_CHIP_RAM.N_207_i ;
    wire A_c_11;
    wire A_c_4;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_1_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire bfn_10_8_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_36 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.N_285 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_a3_0_a3_0 ;
    wire \U712_CHIP_RAM.N_342 ;
    wire \U712_CHIP_RAM.N_328 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_2_i_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_2_i_2 ;
    wire \U712_REG_SM.N_210 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_248_cascade_ ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0 ;
    wire \U712_REG_SM.DS_EN_RNOZ0Z_0 ;
    wire \U712_REG_SM.N_300 ;
    wire \U712_REG_SM.N_228 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire REGENn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.un1_CMA28_0_i ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire CMA_c_5;
    wire A_c_9;
    wire A_c_2;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire A_c_10;
    wire A_c_3;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire A_c_14;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ;
    wire \U712_REG_SM.ASn_0_sqmuxa_1 ;
    wire \U712_REG_SM.N_226 ;
    wire ASn_c;
    wire CONSTANT_ONE_NET;
    wire CMA_c_10;
    wire CMA_c_0;
    wire A_c_17;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_ ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire \U712_CHIP_RAM.un5_DMA_CYCLE_START_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10_cascade_ ;
    wire CLK40_PLL_i;
    wire CLK40_PLL_i_i;
    wire DBRn_c;
    wire C1_c_g;
    wire RESETn_c;
    wire RESETn_c_i;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire WEn_c;
    wire DRA_c_5;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire DRA_c_4;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire RAS0n_c;
    wire AGNUS_REV_c;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire C3_c_g;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire \U712_BYTE_ENABLE.N_315_cascade_ ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_iZ0Z_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire CLK80_PLL;
    wire RESETn_c_i_g;
    wire CASLn_c;
    wire \U712_BYTE_ENABLE.N_311 ;
    wire \U712_BYTE_ENABLE.N_313 ;
    wire N_170;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_iZ0Z_0 ;
    wire N_174_i;
    wire N_172_i;
    wire SIZ_c_1;
    wire \U712_BYTE_ENABLE.un1_CLMBEn_iZ0Z_0 ;
    wire N_176_i;
    wire A_c_1;
    wire CPU_CYCLEm;
    wire DMA_CYCLEm;
    wire CASUn_c;
    wire \U712_BYTE_ENABLE.N_309_cascade_ ;
    wire DBENn_c;
    wire \U712_BYTE_ENABLE.un1_CUUBEn_iZ0Z_0 ;
    wire DS_ENm;
    wire A_c_0;
    wire SIZ_c_0;
    wire N_168;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__3792),
            .RESETB(N__7044),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__11113),
            .DIN(N__11112),
            .DOUT(N__11111),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__11113),
            .PADOUT(N__11112),
            .PADIN(N__11111),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9396),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11104),
            .DIN(N__11103),
            .DOUT(N__11102),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11104),
            .PADOUT(N__11103),
            .PADIN(N__11102),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__11095),
            .DIN(N__11094),
            .DOUT(N__11093),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__11095),
            .PADOUT(N__11094),
            .PADIN(N__11093),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8298),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__11086),
            .DIN(N__11085),
            .DOUT(N__11084),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__11086),
            .PADOUT(N__11085),
            .PADIN(N__11084),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4008),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__11077),
            .DIN(N__11076),
            .DOUT(N__11075),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__11077),
            .PADOUT(N__11076),
            .PADIN(N__11075),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__11068),
            .DIN(N__11067),
            .DOUT(N__11066),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__11068),
            .PADOUT(N__11067),
            .PADIN(N__11066),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__11059),
            .DIN(N__11058),
            .DOUT(N__11057),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__11059),
            .PADOUT(N__11058),
            .PADIN(N__11057),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__11050),
            .DIN(N__11049),
            .DOUT(N__11048),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__11050),
            .PADOUT(N__11049),
            .PADIN(N__11048),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__11041),
            .DIN(N__11040),
            .DOUT(N__11039),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__11041),
            .PADOUT(N__11040),
            .PADIN(N__11039),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__11032),
            .DIN(N__11031),
            .DOUT(N__11030),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__11032),
            .PADOUT(N__11031),
            .PADIN(N__11030),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11023),
            .DIN(N__11022),
            .DOUT(N__11021),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11023),
            .PADOUT(N__11022),
            .PADIN(N__11021),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__11014),
            .DIN(N__11013),
            .DOUT(N__11012),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__11014),
            .PADOUT(N__11013),
            .PADIN(N__11012),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7167),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__11005),
            .DIN(N__11004),
            .DOUT(N__11003),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__11005),
            .PADOUT(N__11004),
            .PADIN(N__11003),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__10996),
            .DIN(N__10995),
            .DOUT(N__10994),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__10996),
            .PADOUT(N__10995),
            .PADIN(N__10994),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4418),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__10987),
            .DIN(N__10986),
            .DOUT(N__10985),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__10987),
            .PADOUT(N__10986),
            .PADIN(N__10985),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__10978),
            .DIN(N__10977),
            .DOUT(N__10976),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__10978),
            .PADOUT(N__10977),
            .PADIN(N__10976),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__10969),
            .DIN(N__10968),
            .DOUT(N__10967),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__10969),
            .PADOUT(N__10968),
            .PADIN(N__10967),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3930),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__10960),
            .DIN(N__10959),
            .DOUT(N__10958),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__10960),
            .PADOUT(N__10959),
            .PADIN(N__10958),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__10951),
            .DIN(N__10950),
            .DOUT(N__10949),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__10951),
            .PADOUT(N__10950),
            .PADIN(N__10949),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__10942),
            .DIN(N__10941),
            .DOUT(N__10940),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__10942),
            .PADOUT(N__10941),
            .PADIN(N__10940),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7017),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__10933),
            .DIN(N__10932),
            .DOUT(N__10931),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__10933),
            .PADOUT(N__10932),
            .PADIN(N__10931),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__10924),
            .DIN(N__10923),
            .DOUT(N__10922),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__10924),
            .PADOUT(N__10923),
            .PADIN(N__10922),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8787),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__10915),
            .DIN(N__10914),
            .DOUT(N__10913),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__10915),
            .PADOUT(N__10914),
            .PADIN(N__10913),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__10906),
            .DIN(N__10905),
            .DOUT(N__10904),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__10906),
            .PADOUT(N__10905),
            .PADIN(N__10904),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__10897),
            .DIN(N__10896),
            .DOUT(N__10895),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__10897),
            .PADOUT(N__10896),
            .PADIN(N__10895),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__10888),
            .DIN(N__10887),
            .DOUT(N__10886),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__10888),
            .PADOUT(N__10887),
            .PADIN(N__10886),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__10879),
            .DIN(N__10878),
            .DOUT(N__10877),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__10879),
            .PADOUT(N__10878),
            .PADIN(N__10877),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__10870),
            .DIN(N__10869),
            .DOUT(N__10868),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__10870),
            .PADOUT(N__10869),
            .PADIN(N__10868),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__10861),
            .DIN(N__10860),
            .DOUT(N__10859),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__10861),
            .PADOUT(N__10860),
            .PADIN(N__10859),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__10852),
            .DIN(N__10851),
            .DOUT(N__10850),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__10852),
            .PADOUT(N__10851),
            .PADIN(N__10850),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__10843),
            .DIN(N__10842),
            .DOUT(N__10841),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__10843),
            .PADOUT(N__10842),
            .PADIN(N__10841),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__10834),
            .DIN(N__10833),
            .DOUT(N__10832),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__10834),
            .PADOUT(N__10833),
            .PADIN(N__10832),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__10825),
            .DIN(N__10824),
            .DOUT(N__10823),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__10825),
            .PADOUT(N__10824),
            .PADIN(N__10823),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__10816),
            .DIN(N__10815),
            .DOUT(N__10814),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__10816),
            .PADOUT(N__10815),
            .PADIN(N__10814),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__10807),
            .DIN(N__10806),
            .DOUT(N__10805),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__10807),
            .PADOUT(N__10806),
            .PADIN(N__10805),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__10798),
            .DIN(N__10797),
            .DOUT(N__10796),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__10798),
            .PADOUT(N__10797),
            .PADIN(N__10796),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9933),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__10789),
            .DIN(N__10788),
            .DOUT(N__10787),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__10789),
            .PADOUT(N__10788),
            .PADIN(N__10787),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7870),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__10780),
            .DIN(N__10779),
            .DOUT(N__10778),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__10780),
            .PADOUT(N__10779),
            .PADIN(N__10778),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__10771),
            .DIN(N__10770),
            .DOUT(N__10769),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__10771),
            .PADOUT(N__10770),
            .PADIN(N__10769),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7500),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__10762),
            .DIN(N__10761),
            .DOUT(N__10760),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__10762),
            .PADOUT(N__10761),
            .PADIN(N__10760),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__10753),
            .DIN(N__10752),
            .DOUT(N__10751),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__10753),
            .PADOUT(N__10752),
            .PADIN(N__10751),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4320),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__10744),
            .DIN(N__10743),
            .DOUT(N__10742),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__10744),
            .PADOUT(N__10743),
            .PADIN(N__10742),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7872),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__10735),
            .DIN(N__10734),
            .DOUT(N__10733),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__10735),
            .PADOUT(N__10734),
            .PADIN(N__10733),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3849),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__10726),
            .DIN(N__10725),
            .DOUT(N__10724),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__10726),
            .PADOUT(N__10725),
            .PADIN(N__10724),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__10717),
            .DIN(N__10716),
            .DOUT(N__10715),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__10717),
            .PADOUT(N__10716),
            .PADIN(N__10715),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7074),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__10708),
            .DIN(N__10707),
            .DOUT(N__10706),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__10708),
            .PADOUT(N__10707),
            .PADIN(N__10706),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6954),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__10699),
            .DIN(N__10698),
            .DOUT(N__10697),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__10699),
            .PADOUT(N__10698),
            .PADIN(N__10697),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__10690),
            .DIN(N__10689),
            .DOUT(N__10688),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__10690),
            .PADOUT(N__10689),
            .PADIN(N__10688),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__10681),
            .DIN(N__10680),
            .DOUT(N__10679),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__10681),
            .PADOUT(N__10680),
            .PADIN(N__10679),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_0_iopad (
            .OE(N__10672),
            .DIN(N__10671),
            .DOUT(N__10670),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__10672),
            .PADOUT(N__10671),
            .PADIN(N__10670),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__10663),
            .DIN(N__10662),
            .DOUT(N__10661),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__10663),
            .PADOUT(N__10662),
            .PADIN(N__10661),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7029),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__10654),
            .DIN(N__10653),
            .DOUT(N__10652),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__10654),
            .PADOUT(N__10653),
            .PADIN(N__10652),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__10645),
            .DIN(N__10644),
            .DOUT(N__10643),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__10645),
            .PADOUT(N__10644),
            .PADIN(N__10643),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7871),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__10636),
            .DIN(N__10635),
            .DOUT(N__10634),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__10636),
            .PADOUT(N__10635),
            .PADIN(N__10634),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7224),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__10627),
            .DIN(N__10626),
            .DOUT(N__10625),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__10627),
            .PADOUT(N__10626),
            .PADIN(N__10625),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8487),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__10618),
            .DIN(N__10617),
            .DOUT(N__10616),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__10618),
            .PADOUT(N__10617),
            .PADIN(N__10616),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4122),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__10609),
            .DIN(N__10608),
            .DOUT(N__10607),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__10609),
            .PADOUT(N__10608),
            .PADIN(N__10607),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7428),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__10600),
            .DIN(N__10599),
            .DOUT(N__10598),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__10600),
            .PADOUT(N__10599),
            .PADIN(N__10598),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6468),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__10591),
            .DIN(N__10590),
            .DOUT(N__10589),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__10591),
            .PADOUT(N__10590),
            .PADIN(N__10589),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__10582),
            .DIN(N__10581),
            .DOUT(N__10580),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__10582),
            .PADOUT(N__10581),
            .PADIN(N__10580),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__10573),
            .DIN(N__10572),
            .DOUT(N__10571),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__10573),
            .PADOUT(N__10572),
            .PADIN(N__10571),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9795),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__10564),
            .DIN(N__10563),
            .DOUT(N__10562),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__10564),
            .PADOUT(N__10563),
            .PADIN(N__10562),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8229),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__10555),
            .DIN(N__10554),
            .DOUT(N__10553),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__10555),
            .PADOUT(N__10554),
            .PADIN(N__10553),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3891),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__10546),
            .DIN(N__10545),
            .DOUT(N__10544),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__10546),
            .PADOUT(N__10545),
            .PADIN(N__10544),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9909),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_obuf_iopad (
            .OE(N__10537),
            .DIN(N__10536),
            .DOUT(N__10535),
            .PACKAGEPIN(DMA_LATCH));
    defparam DMA_LATCH_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_obuf_preio (
            .PADOEN(N__10537),
            .PADOUT(N__10536),
            .PADIN(N__10535),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__10528),
            .DIN(N__10527),
            .DOUT(N__10526),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__10528),
            .PADOUT(N__10527),
            .PADIN(N__10526),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__10519),
            .DIN(N__10518),
            .DOUT(N__10517),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__10519),
            .PADOUT(N__10518),
            .PADIN(N__10517),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__10510),
            .DIN(N__10509),
            .DOUT(N__10508),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__10510),
            .PADOUT(N__10509),
            .PADIN(N__10508),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__10501),
            .DIN(N__10500),
            .DOUT(N__10499),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__10501),
            .PADOUT(N__10500),
            .PADIN(N__10499),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__10492),
            .DIN(N__10491),
            .DOUT(N__10490),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__10492),
            .PADOUT(N__10491),
            .PADIN(N__10490),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6387),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__10483),
            .DIN(N__10482),
            .DOUT(N__10481),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__10483),
            .PADOUT(N__10482),
            .PADIN(N__10481),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__10474),
            .DIN(N__10473),
            .DOUT(N__10472),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__10474),
            .PADOUT(N__10473),
            .PADIN(N__10472),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9897),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__10465),
            .DIN(N__10464),
            .DOUT(N__10463),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__10465),
            .PADOUT(N__10464),
            .PADIN(N__10463),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__3831),
            .DIN0(),
            .DOUT0(N__4269),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__10456),
            .DIN(N__10455),
            .DOUT(N__10454),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__10456),
            .PADOUT(N__10455),
            .PADIN(N__10454),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6423),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__10447),
            .DIN(N__10446),
            .DOUT(N__10445),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__10447),
            .PADOUT(N__10446),
            .PADIN(N__10445),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__10438),
            .DIN(N__10437),
            .DOUT(N__10436),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__10438),
            .PADOUT(N__10437),
            .PADIN(N__10436),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__10429),
            .DIN(N__10428),
            .DOUT(N__10427),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__10429),
            .PADOUT(N__10428),
            .PADIN(N__10427),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6981),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__10420),
            .DIN(N__10419),
            .DOUT(N__10418),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__10420),
            .PADOUT(N__10419),
            .PADIN(N__10418),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__10411),
            .DIN(N__10410),
            .DOUT(N__10409),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__10411),
            .PADOUT(N__10410),
            .PADIN(N__10409),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__10402),
            .DIN(N__10401),
            .DOUT(N__10400),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__10402),
            .PADOUT(N__10401),
            .PADIN(N__10400),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__10393),
            .DIN(N__10392),
            .DOUT(N__10391),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__10393),
            .PADOUT(N__10392),
            .PADIN(N__10391),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__10384),
            .DIN(N__10383),
            .DOUT(N__10382),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__10384),
            .PADOUT(N__10383),
            .PADIN(N__10382),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6879),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__10375),
            .DIN(N__10374),
            .DOUT(N__10373),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__10375),
            .PADOUT(N__10374),
            .PADIN(N__10373),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10152),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__10366),
            .DIN(N__10365),
            .DOUT(N__10364),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__10366),
            .PADOUT(N__10365),
            .PADIN(N__10364),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4548),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__10357),
            .DIN(N__10356),
            .DOUT(N__10355),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__10357),
            .PADOUT(N__10356),
            .PADIN(N__10355),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__10348),
            .DIN(N__10347),
            .DOUT(N__10346),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__10348),
            .PADOUT(N__10347),
            .PADIN(N__10346),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__10339),
            .DIN(N__10338),
            .DOUT(N__10337),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__10339),
            .PADOUT(N__10338),
            .PADIN(N__10337),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6930),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2505 (
            .O(N__10320),
            .I(N__10316));
    InMux I__2504 (
            .O(N__10319),
            .I(N__10313));
    LocalMux I__2503 (
            .O(N__10316),
            .I(N__10308));
    LocalMux I__2502 (
            .O(N__10313),
            .I(N__10308));
    Span12Mux_h I__2501 (
            .O(N__10308),
            .I(N__10304));
    InMux I__2500 (
            .O(N__10307),
            .I(N__10301));
    Odrv12 I__2499 (
            .O(N__10304),
            .I(DS_ENm));
    LocalMux I__2498 (
            .O(N__10301),
            .I(DS_ENm));
    InMux I__2497 (
            .O(N__10296),
            .I(N__10293));
    LocalMux I__2496 (
            .O(N__10293),
            .I(N__10288));
    InMux I__2495 (
            .O(N__10292),
            .I(N__10281));
    InMux I__2494 (
            .O(N__10291),
            .I(N__10281));
    Span4Mux_h I__2493 (
            .O(N__10288),
            .I(N__10278));
    InMux I__2492 (
            .O(N__10287),
            .I(N__10275));
    InMux I__2491 (
            .O(N__10286),
            .I(N__10271));
    LocalMux I__2490 (
            .O(N__10281),
            .I(N__10268));
    Span4Mux_v I__2489 (
            .O(N__10278),
            .I(N__10265));
    LocalMux I__2488 (
            .O(N__10275),
            .I(N__10262));
    InMux I__2487 (
            .O(N__10274),
            .I(N__10259));
    LocalMux I__2486 (
            .O(N__10271),
            .I(N__10254));
    Sp12to4 I__2485 (
            .O(N__10268),
            .I(N__10254));
    Span4Mux_v I__2484 (
            .O(N__10265),
            .I(N__10249));
    Span4Mux_v I__2483 (
            .O(N__10262),
            .I(N__10249));
    LocalMux I__2482 (
            .O(N__10259),
            .I(N__10246));
    Span12Mux_v I__2481 (
            .O(N__10254),
            .I(N__10239));
    Sp12to4 I__2480 (
            .O(N__10249),
            .I(N__10239));
    Span12Mux_s10_v I__2479 (
            .O(N__10246),
            .I(N__10239));
    Span12Mux_h I__2478 (
            .O(N__10239),
            .I(N__10236));
    Odrv12 I__2477 (
            .O(N__10236),
            .I(A_c_0));
    CascadeMux I__2476 (
            .O(N__10233),
            .I(N__10228));
    CascadeMux I__2475 (
            .O(N__10232),
            .I(N__10225));
    InMux I__2474 (
            .O(N__10231),
            .I(N__10222));
    InMux I__2473 (
            .O(N__10228),
            .I(N__10217));
    InMux I__2472 (
            .O(N__10225),
            .I(N__10217));
    LocalMux I__2471 (
            .O(N__10222),
            .I(N__10211));
    LocalMux I__2470 (
            .O(N__10217),
            .I(N__10211));
    InMux I__2469 (
            .O(N__10216),
            .I(N__10208));
    Span4Mux_v I__2468 (
            .O(N__10211),
            .I(N__10204));
    LocalMux I__2467 (
            .O(N__10208),
            .I(N__10201));
    InMux I__2466 (
            .O(N__10207),
            .I(N__10197));
    Span4Mux_v I__2465 (
            .O(N__10204),
            .I(N__10194));
    Span4Mux_h I__2464 (
            .O(N__10201),
            .I(N__10191));
    InMux I__2463 (
            .O(N__10200),
            .I(N__10188));
    LocalMux I__2462 (
            .O(N__10197),
            .I(N__10185));
    Sp12to4 I__2461 (
            .O(N__10194),
            .I(N__10182));
    Span4Mux_v I__2460 (
            .O(N__10191),
            .I(N__10179));
    LocalMux I__2459 (
            .O(N__10188),
            .I(N__10176));
    Span12Mux_v I__2458 (
            .O(N__10185),
            .I(N__10173));
    Span12Mux_h I__2457 (
            .O(N__10182),
            .I(N__10170));
    Sp12to4 I__2456 (
            .O(N__10179),
            .I(N__10165));
    Span12Mux_v I__2455 (
            .O(N__10176),
            .I(N__10165));
    Span12Mux_v I__2454 (
            .O(N__10173),
            .I(N__10162));
    Span12Mux_v I__2453 (
            .O(N__10170),
            .I(N__10157));
    Span12Mux_h I__2452 (
            .O(N__10165),
            .I(N__10157));
    Odrv12 I__2451 (
            .O(N__10162),
            .I(SIZ_c_0));
    Odrv12 I__2450 (
            .O(N__10157),
            .I(SIZ_c_0));
    IoInMux I__2449 (
            .O(N__10152),
            .I(N__10149));
    LocalMux I__2448 (
            .O(N__10149),
            .I(N__10146));
    Span12Mux_s6_v I__2447 (
            .O(N__10146),
            .I(N__10143));
    Odrv12 I__2446 (
            .O(N__10143),
            .I(N_168));
    InMux I__2445 (
            .O(N__10140),
            .I(N__10133));
    InMux I__2444 (
            .O(N__10139),
            .I(N__10130));
    InMux I__2443 (
            .O(N__10138),
            .I(N__10127));
    InMux I__2442 (
            .O(N__10137),
            .I(N__10124));
    InMux I__2441 (
            .O(N__10136),
            .I(N__10121));
    LocalMux I__2440 (
            .O(N__10133),
            .I(N__10112));
    LocalMux I__2439 (
            .O(N__10130),
            .I(N__10105));
    LocalMux I__2438 (
            .O(N__10127),
            .I(N__10102));
    LocalMux I__2437 (
            .O(N__10124),
            .I(N__10075));
    LocalMux I__2436 (
            .O(N__10121),
            .I(N__10072));
    SRMux I__2435 (
            .O(N__10120),
            .I(N__9993));
    SRMux I__2434 (
            .O(N__10119),
            .I(N__9993));
    SRMux I__2433 (
            .O(N__10118),
            .I(N__9993));
    SRMux I__2432 (
            .O(N__10117),
            .I(N__9993));
    SRMux I__2431 (
            .O(N__10116),
            .I(N__9993));
    SRMux I__2430 (
            .O(N__10115),
            .I(N__9993));
    Glb2LocalMux I__2429 (
            .O(N__10112),
            .I(N__9993));
    SRMux I__2428 (
            .O(N__10111),
            .I(N__9993));
    SRMux I__2427 (
            .O(N__10110),
            .I(N__9993));
    SRMux I__2426 (
            .O(N__10109),
            .I(N__9993));
    SRMux I__2425 (
            .O(N__10108),
            .I(N__9993));
    Glb2LocalMux I__2424 (
            .O(N__10105),
            .I(N__9993));
    Glb2LocalMux I__2423 (
            .O(N__10102),
            .I(N__9993));
    SRMux I__2422 (
            .O(N__10101),
            .I(N__9993));
    SRMux I__2421 (
            .O(N__10100),
            .I(N__9993));
    SRMux I__2420 (
            .O(N__10099),
            .I(N__9993));
    SRMux I__2419 (
            .O(N__10098),
            .I(N__9993));
    SRMux I__2418 (
            .O(N__10097),
            .I(N__9993));
    SRMux I__2417 (
            .O(N__10096),
            .I(N__9993));
    SRMux I__2416 (
            .O(N__10095),
            .I(N__9993));
    SRMux I__2415 (
            .O(N__10094),
            .I(N__9993));
    SRMux I__2414 (
            .O(N__10093),
            .I(N__9993));
    SRMux I__2413 (
            .O(N__10092),
            .I(N__9993));
    SRMux I__2412 (
            .O(N__10091),
            .I(N__9993));
    SRMux I__2411 (
            .O(N__10090),
            .I(N__9993));
    SRMux I__2410 (
            .O(N__10089),
            .I(N__9993));
    SRMux I__2409 (
            .O(N__10088),
            .I(N__9993));
    SRMux I__2408 (
            .O(N__10087),
            .I(N__9993));
    SRMux I__2407 (
            .O(N__10086),
            .I(N__9993));
    SRMux I__2406 (
            .O(N__10085),
            .I(N__9993));
    SRMux I__2405 (
            .O(N__10084),
            .I(N__9993));
    SRMux I__2404 (
            .O(N__10083),
            .I(N__9993));
    SRMux I__2403 (
            .O(N__10082),
            .I(N__9993));
    SRMux I__2402 (
            .O(N__10081),
            .I(N__9993));
    SRMux I__2401 (
            .O(N__10080),
            .I(N__9993));
    SRMux I__2400 (
            .O(N__10079),
            .I(N__9993));
    SRMux I__2399 (
            .O(N__10078),
            .I(N__9993));
    Glb2LocalMux I__2398 (
            .O(N__10075),
            .I(N__9993));
    Glb2LocalMux I__2397 (
            .O(N__10072),
            .I(N__9993));
    GlobalMux I__2396 (
            .O(N__9993),
            .I(N__9990));
    gio2CtrlBuf I__2395 (
            .O(N__9990),
            .I(RESETn_c_i_g));
    InMux I__2394 (
            .O(N__9987),
            .I(N__9983));
    CascadeMux I__2393 (
            .O(N__9986),
            .I(N__9979));
    LocalMux I__2392 (
            .O(N__9983),
            .I(N__9976));
    InMux I__2391 (
            .O(N__9982),
            .I(N__9973));
    InMux I__2390 (
            .O(N__9979),
            .I(N__9970));
    Span4Mux_h I__2389 (
            .O(N__9976),
            .I(N__9965));
    LocalMux I__2388 (
            .O(N__9973),
            .I(N__9965));
    LocalMux I__2387 (
            .O(N__9970),
            .I(N__9962));
    Span4Mux_v I__2386 (
            .O(N__9965),
            .I(N__9959));
    Span12Mux_v I__2385 (
            .O(N__9962),
            .I(N__9954));
    Sp12to4 I__2384 (
            .O(N__9959),
            .I(N__9954));
    Span12Mux_h I__2383 (
            .O(N__9954),
            .I(N__9951));
    Span12Mux_v I__2382 (
            .O(N__9951),
            .I(N__9948));
    Odrv12 I__2381 (
            .O(N__9948),
            .I(CASLn_c));
    InMux I__2380 (
            .O(N__9945),
            .I(N__9942));
    LocalMux I__2379 (
            .O(N__9942),
            .I(\U712_BYTE_ENABLE.N_311 ));
    InMux I__2378 (
            .O(N__9939),
            .I(N__9936));
    LocalMux I__2377 (
            .O(N__9936),
            .I(\U712_BYTE_ENABLE.N_313 ));
    IoInMux I__2376 (
            .O(N__9933),
            .I(N__9930));
    LocalMux I__2375 (
            .O(N__9930),
            .I(N__9927));
    Span4Mux_s2_v I__2374 (
            .O(N__9927),
            .I(N__9924));
    Span4Mux_h I__2373 (
            .O(N__9924),
            .I(N__9921));
    Span4Mux_v I__2372 (
            .O(N__9921),
            .I(N__9918));
    Odrv4 I__2371 (
            .O(N__9918),
            .I(N_170));
    InMux I__2370 (
            .O(N__9915),
            .I(N__9912));
    LocalMux I__2369 (
            .O(N__9912),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_iZ0Z_0 ));
    IoInMux I__2368 (
            .O(N__9909),
            .I(N__9906));
    LocalMux I__2367 (
            .O(N__9906),
            .I(N__9903));
    Span12Mux_s11_h I__2366 (
            .O(N__9903),
            .I(N__9900));
    Odrv12 I__2365 (
            .O(N__9900),
            .I(N_174_i));
    IoInMux I__2364 (
            .O(N__9897),
            .I(N__9894));
    LocalMux I__2363 (
            .O(N__9894),
            .I(N__9891));
    IoSpan4Mux I__2362 (
            .O(N__9891),
            .I(N__9888));
    Span4Mux_s3_h I__2361 (
            .O(N__9888),
            .I(N__9885));
    Span4Mux_h I__2360 (
            .O(N__9885),
            .I(N__9882));
    Odrv4 I__2359 (
            .O(N__9882),
            .I(N_172_i));
    InMux I__2358 (
            .O(N__9879),
            .I(N__9872));
    InMux I__2357 (
            .O(N__9878),
            .I(N__9867));
    InMux I__2356 (
            .O(N__9877),
            .I(N__9867));
    CascadeMux I__2355 (
            .O(N__9876),
            .I(N__9864));
    CascadeMux I__2354 (
            .O(N__9875),
            .I(N__9861));
    LocalMux I__2353 (
            .O(N__9872),
            .I(N__9855));
    LocalMux I__2352 (
            .O(N__9867),
            .I(N__9855));
    InMux I__2351 (
            .O(N__9864),
            .I(N__9852));
    InMux I__2350 (
            .O(N__9861),
            .I(N__9849));
    CascadeMux I__2349 (
            .O(N__9860),
            .I(N__9846));
    Span4Mux_v I__2348 (
            .O(N__9855),
            .I(N__9839));
    LocalMux I__2347 (
            .O(N__9852),
            .I(N__9839));
    LocalMux I__2346 (
            .O(N__9849),
            .I(N__9839));
    InMux I__2345 (
            .O(N__9846),
            .I(N__9836));
    Span4Mux_h I__2344 (
            .O(N__9839),
            .I(N__9833));
    LocalMux I__2343 (
            .O(N__9836),
            .I(N__9830));
    Span4Mux_v I__2342 (
            .O(N__9833),
            .I(N__9827));
    Span4Mux_h I__2341 (
            .O(N__9830),
            .I(N__9824));
    Sp12to4 I__2340 (
            .O(N__9827),
            .I(N__9821));
    Span4Mux_v I__2339 (
            .O(N__9824),
            .I(N__9818));
    Span12Mux_h I__2338 (
            .O(N__9821),
            .I(N__9815));
    Sp12to4 I__2337 (
            .O(N__9818),
            .I(N__9812));
    Span12Mux_v I__2336 (
            .O(N__9815),
            .I(N__9809));
    Span12Mux_v I__2335 (
            .O(N__9812),
            .I(N__9806));
    Odrv12 I__2334 (
            .O(N__9809),
            .I(SIZ_c_1));
    Odrv12 I__2333 (
            .O(N__9806),
            .I(SIZ_c_1));
    InMux I__2332 (
            .O(N__9801),
            .I(N__9798));
    LocalMux I__2331 (
            .O(N__9798),
            .I(\U712_BYTE_ENABLE.un1_CLMBEn_iZ0Z_0 ));
    IoInMux I__2330 (
            .O(N__9795),
            .I(N__9792));
    LocalMux I__2329 (
            .O(N__9792),
            .I(N__9789));
    IoSpan4Mux I__2328 (
            .O(N__9789),
            .I(N__9786));
    Span4Mux_s1_h I__2327 (
            .O(N__9786),
            .I(N__9783));
    Sp12to4 I__2326 (
            .O(N__9783),
            .I(N__9780));
    Span12Mux_v I__2325 (
            .O(N__9780),
            .I(N__9777));
    Odrv12 I__2324 (
            .O(N__9777),
            .I(N_176_i));
    InMux I__2323 (
            .O(N__9774),
            .I(N__9771));
    LocalMux I__2322 (
            .O(N__9771),
            .I(N__9767));
    CascadeMux I__2321 (
            .O(N__9770),
            .I(N__9763));
    Span4Mux_v I__2320 (
            .O(N__9767),
            .I(N__9759));
    InMux I__2319 (
            .O(N__9766),
            .I(N__9756));
    InMux I__2318 (
            .O(N__9763),
            .I(N__9751));
    InMux I__2317 (
            .O(N__9762),
            .I(N__9751));
    Span4Mux_v I__2316 (
            .O(N__9759),
            .I(N__9748));
    LocalMux I__2315 (
            .O(N__9756),
            .I(N__9743));
    LocalMux I__2314 (
            .O(N__9751),
            .I(N__9743));
    Span4Mux_v I__2313 (
            .O(N__9748),
            .I(N__9740));
    Sp12to4 I__2312 (
            .O(N__9743),
            .I(N__9737));
    Sp12to4 I__2311 (
            .O(N__9740),
            .I(N__9732));
    Span12Mux_v I__2310 (
            .O(N__9737),
            .I(N__9732));
    Span12Mux_h I__2309 (
            .O(N__9732),
            .I(N__9729));
    Odrv12 I__2308 (
            .O(N__9729),
            .I(A_c_1));
    CascadeMux I__2307 (
            .O(N__9726),
            .I(N__9719));
    InMux I__2306 (
            .O(N__9725),
            .I(N__9713));
    InMux I__2305 (
            .O(N__9724),
            .I(N__9713));
    CascadeMux I__2304 (
            .O(N__9723),
            .I(N__9710));
    CascadeMux I__2303 (
            .O(N__9722),
            .I(N__9706));
    InMux I__2302 (
            .O(N__9719),
            .I(N__9702));
    InMux I__2301 (
            .O(N__9718),
            .I(N__9699));
    LocalMux I__2300 (
            .O(N__9713),
            .I(N__9692));
    InMux I__2299 (
            .O(N__9710),
            .I(N__9689));
    InMux I__2298 (
            .O(N__9709),
            .I(N__9685));
    InMux I__2297 (
            .O(N__9706),
            .I(N__9680));
    InMux I__2296 (
            .O(N__9705),
            .I(N__9677));
    LocalMux I__2295 (
            .O(N__9702),
            .I(N__9674));
    LocalMux I__2294 (
            .O(N__9699),
            .I(N__9671));
    InMux I__2293 (
            .O(N__9698),
            .I(N__9664));
    InMux I__2292 (
            .O(N__9697),
            .I(N__9664));
    InMux I__2291 (
            .O(N__9696),
            .I(N__9664));
    InMux I__2290 (
            .O(N__9695),
            .I(N__9661));
    Span4Mux_v I__2289 (
            .O(N__9692),
            .I(N__9655));
    LocalMux I__2288 (
            .O(N__9689),
            .I(N__9655));
    InMux I__2287 (
            .O(N__9688),
            .I(N__9652));
    LocalMux I__2286 (
            .O(N__9685),
            .I(N__9649));
    CascadeMux I__2285 (
            .O(N__9684),
            .I(N__9643));
    InMux I__2284 (
            .O(N__9683),
            .I(N__9636));
    LocalMux I__2283 (
            .O(N__9680),
            .I(N__9631));
    LocalMux I__2282 (
            .O(N__9677),
            .I(N__9631));
    Span4Mux_h I__2281 (
            .O(N__9674),
            .I(N__9622));
    Span4Mux_v I__2280 (
            .O(N__9671),
            .I(N__9622));
    LocalMux I__2279 (
            .O(N__9664),
            .I(N__9622));
    LocalMux I__2278 (
            .O(N__9661),
            .I(N__9622));
    CascadeMux I__2277 (
            .O(N__9660),
            .I(N__9616));
    Span4Mux_h I__2276 (
            .O(N__9655),
            .I(N__9610));
    LocalMux I__2275 (
            .O(N__9652),
            .I(N__9610));
    Span4Mux_v I__2274 (
            .O(N__9649),
            .I(N__9607));
    InMux I__2273 (
            .O(N__9648),
            .I(N__9602));
    InMux I__2272 (
            .O(N__9647),
            .I(N__9602));
    InMux I__2271 (
            .O(N__9646),
            .I(N__9599));
    InMux I__2270 (
            .O(N__9643),
            .I(N__9594));
    InMux I__2269 (
            .O(N__9642),
            .I(N__9594));
    InMux I__2268 (
            .O(N__9641),
            .I(N__9589));
    InMux I__2267 (
            .O(N__9640),
            .I(N__9589));
    InMux I__2266 (
            .O(N__9639),
            .I(N__9586));
    LocalMux I__2265 (
            .O(N__9636),
            .I(N__9583));
    Span4Mux_v I__2264 (
            .O(N__9631),
            .I(N__9578));
    Span4Mux_h I__2263 (
            .O(N__9622),
            .I(N__9578));
    InMux I__2262 (
            .O(N__9621),
            .I(N__9573));
    InMux I__2261 (
            .O(N__9620),
            .I(N__9573));
    InMux I__2260 (
            .O(N__9619),
            .I(N__9570));
    InMux I__2259 (
            .O(N__9616),
            .I(N__9567));
    InMux I__2258 (
            .O(N__9615),
            .I(N__9564));
    Span4Mux_h I__2257 (
            .O(N__9610),
            .I(N__9561));
    Sp12to4 I__2256 (
            .O(N__9607),
            .I(N__9550));
    LocalMux I__2255 (
            .O(N__9602),
            .I(N__9550));
    LocalMux I__2254 (
            .O(N__9599),
            .I(N__9550));
    LocalMux I__2253 (
            .O(N__9594),
            .I(N__9550));
    LocalMux I__2252 (
            .O(N__9589),
            .I(N__9550));
    LocalMux I__2251 (
            .O(N__9586),
            .I(N__9543));
    Span4Mux_h I__2250 (
            .O(N__9583),
            .I(N__9543));
    Span4Mux_h I__2249 (
            .O(N__9578),
            .I(N__9543));
    LocalMux I__2248 (
            .O(N__9573),
            .I(CPU_CYCLEm));
    LocalMux I__2247 (
            .O(N__9570),
            .I(CPU_CYCLEm));
    LocalMux I__2246 (
            .O(N__9567),
            .I(CPU_CYCLEm));
    LocalMux I__2245 (
            .O(N__9564),
            .I(CPU_CYCLEm));
    Odrv4 I__2244 (
            .O(N__9561),
            .I(CPU_CYCLEm));
    Odrv12 I__2243 (
            .O(N__9550),
            .I(CPU_CYCLEm));
    Odrv4 I__2242 (
            .O(N__9543),
            .I(CPU_CYCLEm));
    InMux I__2241 (
            .O(N__9528),
            .I(N__9525));
    LocalMux I__2240 (
            .O(N__9525),
            .I(N__9519));
    CascadeMux I__2239 (
            .O(N__9524),
            .I(N__9515));
    InMux I__2238 (
            .O(N__9523),
            .I(N__9510));
    InMux I__2237 (
            .O(N__9522),
            .I(N__9507));
    Span4Mux_v I__2236 (
            .O(N__9519),
            .I(N__9504));
    InMux I__2235 (
            .O(N__9518),
            .I(N__9501));
    InMux I__2234 (
            .O(N__9515),
            .I(N__9498));
    InMux I__2233 (
            .O(N__9514),
            .I(N__9495));
    InMux I__2232 (
            .O(N__9513),
            .I(N__9492));
    LocalMux I__2231 (
            .O(N__9510),
            .I(N__9489));
    LocalMux I__2230 (
            .O(N__9507),
            .I(N__9486));
    Sp12to4 I__2229 (
            .O(N__9504),
            .I(N__9477));
    LocalMux I__2228 (
            .O(N__9501),
            .I(N__9477));
    LocalMux I__2227 (
            .O(N__9498),
            .I(N__9477));
    LocalMux I__2226 (
            .O(N__9495),
            .I(N__9477));
    LocalMux I__2225 (
            .O(N__9492),
            .I(N__9473));
    Span12Mux_s8_v I__2224 (
            .O(N__9489),
            .I(N__9470));
    Span12Mux_v I__2223 (
            .O(N__9486),
            .I(N__9465));
    Span12Mux_h I__2222 (
            .O(N__9477),
            .I(N__9465));
    InMux I__2221 (
            .O(N__9476),
            .I(N__9462));
    Span4Mux_h I__2220 (
            .O(N__9473),
            .I(N__9459));
    Odrv12 I__2219 (
            .O(N__9470),
            .I(DMA_CYCLEm));
    Odrv12 I__2218 (
            .O(N__9465),
            .I(DMA_CYCLEm));
    LocalMux I__2217 (
            .O(N__9462),
            .I(DMA_CYCLEm));
    Odrv4 I__2216 (
            .O(N__9459),
            .I(DMA_CYCLEm));
    InMux I__2215 (
            .O(N__9450),
            .I(N__9446));
    InMux I__2214 (
            .O(N__9449),
            .I(N__9443));
    LocalMux I__2213 (
            .O(N__9446),
            .I(N__9439));
    LocalMux I__2212 (
            .O(N__9443),
            .I(N__9436));
    InMux I__2211 (
            .O(N__9442),
            .I(N__9433));
    Span4Mux_v I__2210 (
            .O(N__9439),
            .I(N__9430));
    Span4Mux_v I__2209 (
            .O(N__9436),
            .I(N__9427));
    LocalMux I__2208 (
            .O(N__9433),
            .I(N__9424));
    Sp12to4 I__2207 (
            .O(N__9430),
            .I(N__9419));
    Sp12to4 I__2206 (
            .O(N__9427),
            .I(N__9419));
    Span4Mux_v I__2205 (
            .O(N__9424),
            .I(N__9416));
    Span12Mux_h I__2204 (
            .O(N__9419),
            .I(N__9413));
    Sp12to4 I__2203 (
            .O(N__9416),
            .I(N__9410));
    Span12Mux_v I__2202 (
            .O(N__9413),
            .I(N__9407));
    Span12Mux_v I__2201 (
            .O(N__9410),
            .I(N__9404));
    Odrv12 I__2200 (
            .O(N__9407),
            .I(CASUn_c));
    Odrv12 I__2199 (
            .O(N__9404),
            .I(CASUn_c));
    CascadeMux I__2198 (
            .O(N__9399),
            .I(\U712_BYTE_ENABLE.N_309_cascade_ ));
    IoInMux I__2197 (
            .O(N__9396),
            .I(N__9393));
    LocalMux I__2196 (
            .O(N__9393),
            .I(N__9389));
    InMux I__2195 (
            .O(N__9392),
            .I(N__9386));
    IoSpan4Mux I__2194 (
            .O(N__9389),
            .I(N__9382));
    LocalMux I__2193 (
            .O(N__9386),
            .I(N__9379));
    InMux I__2192 (
            .O(N__9385),
            .I(N__9376));
    Sp12to4 I__2191 (
            .O(N__9382),
            .I(N__9371));
    Span4Mux_v I__2190 (
            .O(N__9379),
            .I(N__9368));
    LocalMux I__2189 (
            .O(N__9376),
            .I(N__9365));
    InMux I__2188 (
            .O(N__9375),
            .I(N__9362));
    InMux I__2187 (
            .O(N__9374),
            .I(N__9359));
    Span12Mux_s7_v I__2186 (
            .O(N__9371),
            .I(N__9355));
    Sp12to4 I__2185 (
            .O(N__9368),
            .I(N__9346));
    Sp12to4 I__2184 (
            .O(N__9365),
            .I(N__9346));
    LocalMux I__2183 (
            .O(N__9362),
            .I(N__9346));
    LocalMux I__2182 (
            .O(N__9359),
            .I(N__9346));
    InMux I__2181 (
            .O(N__9358),
            .I(N__9343));
    Odrv12 I__2180 (
            .O(N__9355),
            .I(DBENn_c));
    Odrv12 I__2179 (
            .O(N__9346),
            .I(DBENn_c));
    LocalMux I__2178 (
            .O(N__9343),
            .I(DBENn_c));
    InMux I__2177 (
            .O(N__9336),
            .I(N__9333));
    LocalMux I__2176 (
            .O(N__9333),
            .I(\U712_BYTE_ENABLE.un1_CUUBEn_iZ0Z_0 ));
    InMux I__2175 (
            .O(N__9330),
            .I(N__9325));
    InMux I__2174 (
            .O(N__9329),
            .I(N__9319));
    InMux I__2173 (
            .O(N__9328),
            .I(N__9319));
    LocalMux I__2172 (
            .O(N__9325),
            .I(N__9316));
    InMux I__2171 (
            .O(N__9324),
            .I(N__9313));
    LocalMux I__2170 (
            .O(N__9319),
            .I(N__9310));
    Span4Mux_h I__2169 (
            .O(N__9316),
            .I(N__9305));
    LocalMux I__2168 (
            .O(N__9313),
            .I(N__9305));
    Span4Mux_v I__2167 (
            .O(N__9310),
            .I(N__9302));
    Span4Mux_v I__2166 (
            .O(N__9305),
            .I(N__9299));
    Span4Mux_v I__2165 (
            .O(N__9302),
            .I(N__9296));
    Span4Mux_v I__2164 (
            .O(N__9299),
            .I(N__9293));
    Sp12to4 I__2163 (
            .O(N__9296),
            .I(N__9290));
    Sp12to4 I__2162 (
            .O(N__9293),
            .I(N__9287));
    Span12Mux_h I__2161 (
            .O(N__9290),
            .I(N__9284));
    Span12Mux_h I__2160 (
            .O(N__9287),
            .I(N__9281));
    Odrv12 I__2159 (
            .O(N__9284),
            .I(DRA_c_4));
    Odrv12 I__2158 (
            .O(N__9281),
            .I(DRA_c_4));
    InMux I__2157 (
            .O(N__9276),
            .I(N__9273));
    LocalMux I__2156 (
            .O(N__9273),
            .I(N__9268));
    InMux I__2155 (
            .O(N__9272),
            .I(N__9263));
    InMux I__2154 (
            .O(N__9271),
            .I(N__9263));
    Span4Mux_h I__2153 (
            .O(N__9268),
            .I(N__9258));
    LocalMux I__2152 (
            .O(N__9263),
            .I(N__9258));
    Span4Mux_v I__2151 (
            .O(N__9258),
            .I(N__9254));
    InMux I__2150 (
            .O(N__9257),
            .I(N__9251));
    Span4Mux_v I__2149 (
            .O(N__9254),
            .I(N__9248));
    LocalMux I__2148 (
            .O(N__9251),
            .I(N__9245));
    Sp12to4 I__2147 (
            .O(N__9248),
            .I(N__9240));
    Span12Mux_v I__2146 (
            .O(N__9245),
            .I(N__9240));
    Span12Mux_h I__2145 (
            .O(N__9240),
            .I(N__9237));
    Odrv12 I__2144 (
            .O(N__9237),
            .I(DRA_c_3));
    InMux I__2143 (
            .O(N__9234),
            .I(N__9231));
    LocalMux I__2142 (
            .O(N__9231),
            .I(N__9228));
    Span4Mux_h I__2141 (
            .O(N__9228),
            .I(N__9225));
    Odrv4 I__2140 (
            .O(N__9225),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2139 (
            .O(N__9222),
            .I(N__9217));
    InMux I__2138 (
            .O(N__9221),
            .I(N__9214));
    InMux I__2137 (
            .O(N__9220),
            .I(N__9211));
    LocalMux I__2136 (
            .O(N__9217),
            .I(N__9207));
    LocalMux I__2135 (
            .O(N__9214),
            .I(N__9202));
    LocalMux I__2134 (
            .O(N__9211),
            .I(N__9202));
    InMux I__2133 (
            .O(N__9210),
            .I(N__9199));
    Span4Mux_v I__2132 (
            .O(N__9207),
            .I(N__9196));
    Sp12to4 I__2131 (
            .O(N__9202),
            .I(N__9191));
    LocalMux I__2130 (
            .O(N__9199),
            .I(N__9191));
    Sp12to4 I__2129 (
            .O(N__9196),
            .I(N__9188));
    Span12Mux_v I__2128 (
            .O(N__9191),
            .I(N__9185));
    Span12Mux_h I__2127 (
            .O(N__9188),
            .I(N__9182));
    Span12Mux_h I__2126 (
            .O(N__9185),
            .I(N__9179));
    Odrv12 I__2125 (
            .O(N__9182),
            .I(DRA_c_8));
    Odrv12 I__2124 (
            .O(N__9179),
            .I(DRA_c_8));
    InMux I__2123 (
            .O(N__9174),
            .I(N__9171));
    LocalMux I__2122 (
            .O(N__9171),
            .I(N__9168));
    Span4Mux_h I__2121 (
            .O(N__9168),
            .I(N__9165));
    Odrv4 I__2120 (
            .O(N__9165),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2119 (
            .O(N__9162),
            .I(N__9159));
    LocalMux I__2118 (
            .O(N__9159),
            .I(N__9155));
    InMux I__2117 (
            .O(N__9158),
            .I(N__9152));
    Span4Mux_v I__2116 (
            .O(N__9155),
            .I(N__9149));
    LocalMux I__2115 (
            .O(N__9152),
            .I(N__9146));
    Sp12to4 I__2114 (
            .O(N__9149),
            .I(N__9143));
    Span12Mux_v I__2113 (
            .O(N__9146),
            .I(N__9140));
    Span12Mux_h I__2112 (
            .O(N__9143),
            .I(N__9137));
    Span12Mux_h I__2111 (
            .O(N__9140),
            .I(N__9134));
    Odrv12 I__2110 (
            .O(N__9137),
            .I(RAS0n_c));
    Odrv12 I__2109 (
            .O(N__9134),
            .I(RAS0n_c));
    InMux I__2108 (
            .O(N__9129),
            .I(N__9126));
    LocalMux I__2107 (
            .O(N__9126),
            .I(N__9115));
    InMux I__2106 (
            .O(N__9125),
            .I(N__9112));
    CascadeMux I__2105 (
            .O(N__9124),
            .I(N__9108));
    CascadeMux I__2104 (
            .O(N__9123),
            .I(N__9105));
    CascadeMux I__2103 (
            .O(N__9122),
            .I(N__9102));
    CascadeMux I__2102 (
            .O(N__9121),
            .I(N__9096));
    CascadeMux I__2101 (
            .O(N__9120),
            .I(N__9093));
    CascadeMux I__2100 (
            .O(N__9119),
            .I(N__9089));
    CascadeMux I__2099 (
            .O(N__9118),
            .I(N__9085));
    Span4Mux_h I__2098 (
            .O(N__9115),
            .I(N__9080));
    LocalMux I__2097 (
            .O(N__9112),
            .I(N__9077));
    InMux I__2096 (
            .O(N__9111),
            .I(N__9063));
    InMux I__2095 (
            .O(N__9108),
            .I(N__9063));
    InMux I__2094 (
            .O(N__9105),
            .I(N__9063));
    InMux I__2093 (
            .O(N__9102),
            .I(N__9063));
    InMux I__2092 (
            .O(N__9101),
            .I(N__9063));
    InMux I__2091 (
            .O(N__9100),
            .I(N__9063));
    InMux I__2090 (
            .O(N__9099),
            .I(N__9060));
    InMux I__2089 (
            .O(N__9096),
            .I(N__9045));
    InMux I__2088 (
            .O(N__9093),
            .I(N__9045));
    InMux I__2087 (
            .O(N__9092),
            .I(N__9045));
    InMux I__2086 (
            .O(N__9089),
            .I(N__9045));
    InMux I__2085 (
            .O(N__9088),
            .I(N__9045));
    InMux I__2084 (
            .O(N__9085),
            .I(N__9045));
    InMux I__2083 (
            .O(N__9084),
            .I(N__9045));
    CascadeMux I__2082 (
            .O(N__9083),
            .I(N__9042));
    Span4Mux_v I__2081 (
            .O(N__9080),
            .I(N__9035));
    Span4Mux_v I__2080 (
            .O(N__9077),
            .I(N__9035));
    InMux I__2079 (
            .O(N__9076),
            .I(N__9032));
    LocalMux I__2078 (
            .O(N__9063),
            .I(N__9029));
    LocalMux I__2077 (
            .O(N__9060),
            .I(N__9026));
    LocalMux I__2076 (
            .O(N__9045),
            .I(N__9023));
    InMux I__2075 (
            .O(N__9042),
            .I(N__9018));
    InMux I__2074 (
            .O(N__9041),
            .I(N__9018));
    InMux I__2073 (
            .O(N__9040),
            .I(N__9015));
    Sp12to4 I__2072 (
            .O(N__9035),
            .I(N__9011));
    LocalMux I__2071 (
            .O(N__9032),
            .I(N__9008));
    Span4Mux_v I__2070 (
            .O(N__9029),
            .I(N__9003));
    Span4Mux_h I__2069 (
            .O(N__9026),
            .I(N__9003));
    Span4Mux_v I__2068 (
            .O(N__9023),
            .I(N__9000));
    LocalMux I__2067 (
            .O(N__9018),
            .I(N__8995));
    LocalMux I__2066 (
            .O(N__9015),
            .I(N__8995));
    InMux I__2065 (
            .O(N__9014),
            .I(N__8992));
    Span12Mux_h I__2064 (
            .O(N__9011),
            .I(N__8983));
    Span12Mux_v I__2063 (
            .O(N__9008),
            .I(N__8983));
    Sp12to4 I__2062 (
            .O(N__9003),
            .I(N__8983));
    Sp12to4 I__2061 (
            .O(N__9000),
            .I(N__8983));
    Sp12to4 I__2060 (
            .O(N__8995),
            .I(N__8978));
    LocalMux I__2059 (
            .O(N__8992),
            .I(N__8978));
    Span12Mux_v I__2058 (
            .O(N__8983),
            .I(N__8975));
    Span12Mux_v I__2057 (
            .O(N__8978),
            .I(N__8972));
    Span12Mux_h I__2056 (
            .O(N__8975),
            .I(N__8969));
    Span12Mux_h I__2055 (
            .O(N__8972),
            .I(N__8966));
    Odrv12 I__2054 (
            .O(N__8969),
            .I(AGNUS_REV_c));
    Odrv12 I__2053 (
            .O(N__8966),
            .I(AGNUS_REV_c));
    InMux I__2052 (
            .O(N__8961),
            .I(N__8957));
    CascadeMux I__2051 (
            .O(N__8960),
            .I(N__8954));
    LocalMux I__2050 (
            .O(N__8957),
            .I(N__8951));
    InMux I__2049 (
            .O(N__8954),
            .I(N__8948));
    Span4Mux_h I__2048 (
            .O(N__8951),
            .I(N__8941));
    LocalMux I__2047 (
            .O(N__8948),
            .I(N__8941));
    InMux I__2046 (
            .O(N__8947),
            .I(N__8938));
    InMux I__2045 (
            .O(N__8946),
            .I(N__8935));
    Span4Mux_v I__2044 (
            .O(N__8941),
            .I(N__8932));
    LocalMux I__2043 (
            .O(N__8938),
            .I(N__8927));
    LocalMux I__2042 (
            .O(N__8935),
            .I(N__8927));
    Sp12to4 I__2041 (
            .O(N__8932),
            .I(N__8922));
    Span12Mux_v I__2040 (
            .O(N__8927),
            .I(N__8922));
    Span12Mux_h I__2039 (
            .O(N__8922),
            .I(N__8919));
    Span12Mux_v I__2038 (
            .O(N__8919),
            .I(N__8916));
    Odrv12 I__2037 (
            .O(N__8916),
            .I(DRA_c_9));
    InMux I__2036 (
            .O(N__8913),
            .I(N__8910));
    LocalMux I__2035 (
            .O(N__8910),
            .I(N__8907));
    Span4Mux_v I__2034 (
            .O(N__8907),
            .I(N__8904));
    Odrv4 I__2033 (
            .O(N__8904),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    InMux I__2032 (
            .O(N__8901),
            .I(N__8898));
    LocalMux I__2031 (
            .O(N__8898),
            .I(N__8890));
    ClkMux I__2030 (
            .O(N__8897),
            .I(N__8877));
    ClkMux I__2029 (
            .O(N__8896),
            .I(N__8877));
    ClkMux I__2028 (
            .O(N__8895),
            .I(N__8877));
    ClkMux I__2027 (
            .O(N__8894),
            .I(N__8877));
    ClkMux I__2026 (
            .O(N__8893),
            .I(N__8877));
    Glb2LocalMux I__2025 (
            .O(N__8890),
            .I(N__8877));
    GlobalMux I__2024 (
            .O(N__8877),
            .I(N__8874));
    gio2CtrlBuf I__2023 (
            .O(N__8874),
            .I(C3_c_g));
    CEMux I__2022 (
            .O(N__8871),
            .I(N__8867));
    CEMux I__2021 (
            .O(N__8870),
            .I(N__8863));
    LocalMux I__2020 (
            .O(N__8867),
            .I(N__8860));
    CEMux I__2019 (
            .O(N__8866),
            .I(N__8857));
    LocalMux I__2018 (
            .O(N__8863),
            .I(N__8849));
    Span4Mux_v I__2017 (
            .O(N__8860),
            .I(N__8849));
    LocalMux I__2016 (
            .O(N__8857),
            .I(N__8849));
    CEMux I__2015 (
            .O(N__8856),
            .I(N__8846));
    Span4Mux_v I__2014 (
            .O(N__8849),
            .I(N__8841));
    LocalMux I__2013 (
            .O(N__8846),
            .I(N__8841));
    Span4Mux_v I__2012 (
            .O(N__8841),
            .I(N__8838));
    Odrv4 I__2011 (
            .O(N__8838),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ));
    CascadeMux I__2010 (
            .O(N__8835),
            .I(N__8831));
    InMux I__2009 (
            .O(N__8834),
            .I(N__8828));
    InMux I__2008 (
            .O(N__8831),
            .I(N__8825));
    LocalMux I__2007 (
            .O(N__8828),
            .I(N__8822));
    LocalMux I__2006 (
            .O(N__8825),
            .I(N__8818));
    Span4Mux_v I__2005 (
            .O(N__8822),
            .I(N__8815));
    InMux I__2004 (
            .O(N__8821),
            .I(N__8810));
    Span4Mux_v I__2003 (
            .O(N__8818),
            .I(N__8807));
    Span4Mux_h I__2002 (
            .O(N__8815),
            .I(N__8804));
    InMux I__2001 (
            .O(N__8814),
            .I(N__8801));
    InMux I__2000 (
            .O(N__8813),
            .I(N__8798));
    LocalMux I__1999 (
            .O(N__8810),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1998 (
            .O(N__8807),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1997 (
            .O(N__8804),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1996 (
            .O(N__8801),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1995 (
            .O(N__8798),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1994 (
            .O(N__8787),
            .I(N__8784));
    LocalMux I__1993 (
            .O(N__8784),
            .I(N__8781));
    Span4Mux_s3_v I__1992 (
            .O(N__8781),
            .I(N__8778));
    Span4Mux_v I__1991 (
            .O(N__8778),
            .I(N__8775));
    Span4Mux_h I__1990 (
            .O(N__8775),
            .I(N__8772));
    Odrv4 I__1989 (
            .O(N__8772),
            .I(CRCSn_c));
    CascadeMux I__1988 (
            .O(N__8769),
            .I(\U712_BYTE_ENABLE.N_315_cascade_ ));
    InMux I__1987 (
            .O(N__8766),
            .I(N__8763));
    LocalMux I__1986 (
            .O(N__8763),
            .I(N__8760));
    Span4Mux_v I__1985 (
            .O(N__8760),
            .I(N__8757));
    Span4Mux_h I__1984 (
            .O(N__8757),
            .I(N__8754));
    Odrv4 I__1983 (
            .O(N__8754),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_iZ0Z_0 ));
    InMux I__1982 (
            .O(N__8751),
            .I(N__8747));
    InMux I__1981 (
            .O(N__8750),
            .I(N__8744));
    LocalMux I__1980 (
            .O(N__8747),
            .I(N__8739));
    LocalMux I__1979 (
            .O(N__8744),
            .I(N__8739));
    Odrv4 I__1978 (
            .O(N__8739),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__1977 (
            .O(N__8736),
            .I(N__8733));
    LocalMux I__1976 (
            .O(N__8733),
            .I(N__8707));
    ClkMux I__1975 (
            .O(N__8732),
            .I(N__8628));
    ClkMux I__1974 (
            .O(N__8731),
            .I(N__8628));
    ClkMux I__1973 (
            .O(N__8730),
            .I(N__8628));
    ClkMux I__1972 (
            .O(N__8729),
            .I(N__8628));
    ClkMux I__1971 (
            .O(N__8728),
            .I(N__8628));
    ClkMux I__1970 (
            .O(N__8727),
            .I(N__8628));
    ClkMux I__1969 (
            .O(N__8726),
            .I(N__8628));
    ClkMux I__1968 (
            .O(N__8725),
            .I(N__8628));
    ClkMux I__1967 (
            .O(N__8724),
            .I(N__8628));
    ClkMux I__1966 (
            .O(N__8723),
            .I(N__8628));
    ClkMux I__1965 (
            .O(N__8722),
            .I(N__8628));
    ClkMux I__1964 (
            .O(N__8721),
            .I(N__8628));
    ClkMux I__1963 (
            .O(N__8720),
            .I(N__8628));
    ClkMux I__1962 (
            .O(N__8719),
            .I(N__8628));
    ClkMux I__1961 (
            .O(N__8718),
            .I(N__8628));
    ClkMux I__1960 (
            .O(N__8717),
            .I(N__8628));
    ClkMux I__1959 (
            .O(N__8716),
            .I(N__8628));
    ClkMux I__1958 (
            .O(N__8715),
            .I(N__8628));
    ClkMux I__1957 (
            .O(N__8714),
            .I(N__8628));
    ClkMux I__1956 (
            .O(N__8713),
            .I(N__8628));
    ClkMux I__1955 (
            .O(N__8712),
            .I(N__8628));
    ClkMux I__1954 (
            .O(N__8711),
            .I(N__8628));
    ClkMux I__1953 (
            .O(N__8710),
            .I(N__8628));
    Glb2LocalMux I__1952 (
            .O(N__8707),
            .I(N__8628));
    ClkMux I__1951 (
            .O(N__8706),
            .I(N__8628));
    ClkMux I__1950 (
            .O(N__8705),
            .I(N__8628));
    ClkMux I__1949 (
            .O(N__8704),
            .I(N__8628));
    ClkMux I__1948 (
            .O(N__8703),
            .I(N__8628));
    ClkMux I__1947 (
            .O(N__8702),
            .I(N__8628));
    ClkMux I__1946 (
            .O(N__8701),
            .I(N__8628));
    ClkMux I__1945 (
            .O(N__8700),
            .I(N__8628));
    ClkMux I__1944 (
            .O(N__8699),
            .I(N__8628));
    ClkMux I__1943 (
            .O(N__8698),
            .I(N__8628));
    ClkMux I__1942 (
            .O(N__8697),
            .I(N__8628));
    GlobalMux I__1941 (
            .O(N__8628),
            .I(CLK80_PLL));
    InMux I__1940 (
            .O(N__8625),
            .I(N__8622));
    LocalMux I__1939 (
            .O(N__8622),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__1938 (
            .O(N__8619),
            .I(N__8616));
    LocalMux I__1937 (
            .O(N__8616),
            .I(N__8613));
    Odrv4 I__1936 (
            .O(N__8613),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__1935 (
            .O(N__8610),
            .I(N__8602));
    InMux I__1934 (
            .O(N__8609),
            .I(N__8602));
    InMux I__1933 (
            .O(N__8608),
            .I(N__8599));
    InMux I__1932 (
            .O(N__8607),
            .I(N__8596));
    LocalMux I__1931 (
            .O(N__8602),
            .I(N__8589));
    LocalMux I__1930 (
            .O(N__8599),
            .I(N__8589));
    LocalMux I__1929 (
            .O(N__8596),
            .I(N__8589));
    Span4Mux_v I__1928 (
            .O(N__8589),
            .I(N__8586));
    Sp12to4 I__1927 (
            .O(N__8586),
            .I(N__8583));
    Span12Mux_h I__1926 (
            .O(N__8583),
            .I(N__8580));
    Odrv12 I__1925 (
            .O(N__8580),
            .I(DRA_c_7));
    InMux I__1924 (
            .O(N__8577),
            .I(N__8574));
    LocalMux I__1923 (
            .O(N__8574),
            .I(N__8571));
    Span4Mux_h I__1922 (
            .O(N__8571),
            .I(N__8568));
    Odrv4 I__1921 (
            .O(N__8568),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    CEMux I__1920 (
            .O(N__8565),
            .I(N__8562));
    LocalMux I__1919 (
            .O(N__8562),
            .I(N__8558));
    CEMux I__1918 (
            .O(N__8561),
            .I(N__8554));
    Span4Mux_v I__1917 (
            .O(N__8558),
            .I(N__8551));
    CEMux I__1916 (
            .O(N__8557),
            .I(N__8548));
    LocalMux I__1915 (
            .O(N__8554),
            .I(N__8545));
    Odrv4 I__1914 (
            .O(N__8551),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ));
    LocalMux I__1913 (
            .O(N__8548),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ));
    Odrv12 I__1912 (
            .O(N__8545),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ));
    InMux I__1911 (
            .O(N__8538),
            .I(N__8535));
    LocalMux I__1910 (
            .O(N__8535),
            .I(N__8531));
    InMux I__1909 (
            .O(N__8534),
            .I(N__8528));
    Odrv12 I__1908 (
            .O(N__8531),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__1907 (
            .O(N__8528),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1906 (
            .O(N__8523),
            .I(N__8520));
    LocalMux I__1905 (
            .O(N__8520),
            .I(N__8516));
    InMux I__1904 (
            .O(N__8519),
            .I(N__8513));
    Sp12to4 I__1903 (
            .O(N__8516),
            .I(N__8509));
    LocalMux I__1902 (
            .O(N__8513),
            .I(N__8506));
    InMux I__1901 (
            .O(N__8512),
            .I(N__8503));
    Span12Mux_v I__1900 (
            .O(N__8509),
            .I(N__8500));
    Span4Mux_v I__1899 (
            .O(N__8506),
            .I(N__8497));
    LocalMux I__1898 (
            .O(N__8503),
            .I(N__8494));
    Odrv12 I__1897 (
            .O(N__8500),
            .I(REG_CYCLEm));
    Odrv4 I__1896 (
            .O(N__8497),
            .I(REG_CYCLEm));
    Odrv12 I__1895 (
            .O(N__8494),
            .I(REG_CYCLEm));
    IoInMux I__1894 (
            .O(N__8487),
            .I(N__8484));
    LocalMux I__1893 (
            .O(N__8484),
            .I(N__8481));
    IoSpan4Mux I__1892 (
            .O(N__8481),
            .I(N__8478));
    IoSpan4Mux I__1891 (
            .O(N__8478),
            .I(N__8475));
    Sp12to4 I__1890 (
            .O(N__8475),
            .I(N__8472));
    Span12Mux_s7_h I__1889 (
            .O(N__8472),
            .I(N__8469));
    Odrv12 I__1888 (
            .O(N__8469),
            .I(DRDENn_c));
    InMux I__1887 (
            .O(N__8466),
            .I(N__8463));
    LocalMux I__1886 (
            .O(N__8463),
            .I(N__8453));
    CascadeMux I__1885 (
            .O(N__8462),
            .I(N__8450));
    CascadeMux I__1884 (
            .O(N__8461),
            .I(N__8447));
    CascadeMux I__1883 (
            .O(N__8460),
            .I(N__8444));
    InMux I__1882 (
            .O(N__8459),
            .I(N__8440));
    CascadeMux I__1881 (
            .O(N__8458),
            .I(N__8437));
    CascadeMux I__1880 (
            .O(N__8457),
            .I(N__8434));
    CascadeMux I__1879 (
            .O(N__8456),
            .I(N__8431));
    Span4Mux_h I__1878 (
            .O(N__8453),
            .I(N__8427));
    InMux I__1877 (
            .O(N__8450),
            .I(N__8420));
    InMux I__1876 (
            .O(N__8447),
            .I(N__8420));
    InMux I__1875 (
            .O(N__8444),
            .I(N__8420));
    InMux I__1874 (
            .O(N__8443),
            .I(N__8417));
    LocalMux I__1873 (
            .O(N__8440),
            .I(N__8414));
    InMux I__1872 (
            .O(N__8437),
            .I(N__8411));
    InMux I__1871 (
            .O(N__8434),
            .I(N__8408));
    InMux I__1870 (
            .O(N__8431),
            .I(N__8400));
    CascadeMux I__1869 (
            .O(N__8430),
            .I(N__8393));
    Span4Mux_v I__1868 (
            .O(N__8427),
            .I(N__8386));
    LocalMux I__1867 (
            .O(N__8420),
            .I(N__8386));
    LocalMux I__1866 (
            .O(N__8417),
            .I(N__8386));
    Span4Mux_h I__1865 (
            .O(N__8414),
            .I(N__8379));
    LocalMux I__1864 (
            .O(N__8411),
            .I(N__8379));
    LocalMux I__1863 (
            .O(N__8408),
            .I(N__8379));
    InMux I__1862 (
            .O(N__8407),
            .I(N__8370));
    InMux I__1861 (
            .O(N__8406),
            .I(N__8370));
    InMux I__1860 (
            .O(N__8405),
            .I(N__8370));
    InMux I__1859 (
            .O(N__8404),
            .I(N__8370));
    CascadeMux I__1858 (
            .O(N__8403),
            .I(N__8365));
    LocalMux I__1857 (
            .O(N__8400),
            .I(N__8361));
    CascadeMux I__1856 (
            .O(N__8399),
            .I(N__8357));
    InMux I__1855 (
            .O(N__8398),
            .I(N__8350));
    InMux I__1854 (
            .O(N__8397),
            .I(N__8350));
    InMux I__1853 (
            .O(N__8396),
            .I(N__8350));
    InMux I__1852 (
            .O(N__8393),
            .I(N__8347));
    Span4Mux_h I__1851 (
            .O(N__8386),
            .I(N__8344));
    Span4Mux_v I__1850 (
            .O(N__8379),
            .I(N__8339));
    LocalMux I__1849 (
            .O(N__8370),
            .I(N__8339));
    InMux I__1848 (
            .O(N__8369),
            .I(N__8336));
    InMux I__1847 (
            .O(N__8368),
            .I(N__8333));
    InMux I__1846 (
            .O(N__8365),
            .I(N__8328));
    InMux I__1845 (
            .O(N__8364),
            .I(N__8328));
    Span4Mux_h I__1844 (
            .O(N__8361),
            .I(N__8325));
    InMux I__1843 (
            .O(N__8360),
            .I(N__8320));
    InMux I__1842 (
            .O(N__8357),
            .I(N__8320));
    LocalMux I__1841 (
            .O(N__8350),
            .I(N__8317));
    LocalMux I__1840 (
            .O(N__8347),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1839 (
            .O(N__8344),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1838 (
            .O(N__8339),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1837 (
            .O(N__8336),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1836 (
            .O(N__8333),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1835 (
            .O(N__8328),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1834 (
            .O(N__8325),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1833 (
            .O(N__8320),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1832 (
            .O(N__8317),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__1831 (
            .O(N__8298),
            .I(N__8295));
    LocalMux I__1830 (
            .O(N__8295),
            .I(N__8292));
    Span4Mux_s0_v I__1829 (
            .O(N__8292),
            .I(N__8289));
    Sp12to4 I__1828 (
            .O(N__8289),
            .I(N__8286));
    Span12Mux_h I__1827 (
            .O(N__8286),
            .I(N__8283));
    Odrv12 I__1826 (
            .O(N__8283),
            .I(CASn_c));
    InMux I__1825 (
            .O(N__8280),
            .I(N__8276));
    InMux I__1824 (
            .O(N__8279),
            .I(N__8273));
    LocalMux I__1823 (
            .O(N__8276),
            .I(N__8266));
    LocalMux I__1822 (
            .O(N__8273),
            .I(N__8263));
    InMux I__1821 (
            .O(N__8272),
            .I(N__8256));
    InMux I__1820 (
            .O(N__8271),
            .I(N__8256));
    InMux I__1819 (
            .O(N__8270),
            .I(N__8256));
    CascadeMux I__1818 (
            .O(N__8269),
            .I(N__8252));
    Span4Mux_v I__1817 (
            .O(N__8266),
            .I(N__8249));
    Span4Mux_v I__1816 (
            .O(N__8263),
            .I(N__8244));
    LocalMux I__1815 (
            .O(N__8256),
            .I(N__8244));
    InMux I__1814 (
            .O(N__8255),
            .I(N__8241));
    InMux I__1813 (
            .O(N__8252),
            .I(N__8238));
    Odrv4 I__1812 (
            .O(N__8249),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1811 (
            .O(N__8244),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1810 (
            .O(N__8241),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1809 (
            .O(N__8238),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1808 (
            .O(N__8229),
            .I(N__8226));
    LocalMux I__1807 (
            .O(N__8226),
            .I(N__8223));
    Span4Mux_s2_h I__1806 (
            .O(N__8223),
            .I(N__8220));
    Sp12to4 I__1805 (
            .O(N__8220),
            .I(N__8217));
    Span12Mux_s7_v I__1804 (
            .O(N__8217),
            .I(N__8214));
    Span12Mux_h I__1803 (
            .O(N__8214),
            .I(N__8211));
    Odrv12 I__1802 (
            .O(N__8211),
            .I(WEn_c));
    InMux I__1801 (
            .O(N__8208),
            .I(N__8202));
    InMux I__1800 (
            .O(N__8207),
            .I(N__8199));
    InMux I__1799 (
            .O(N__8206),
            .I(N__8196));
    InMux I__1798 (
            .O(N__8205),
            .I(N__8193));
    LocalMux I__1797 (
            .O(N__8202),
            .I(N__8184));
    LocalMux I__1796 (
            .O(N__8199),
            .I(N__8184));
    LocalMux I__1795 (
            .O(N__8196),
            .I(N__8184));
    LocalMux I__1794 (
            .O(N__8193),
            .I(N__8184));
    Sp12to4 I__1793 (
            .O(N__8184),
            .I(N__8181));
    Span12Mux_v I__1792 (
            .O(N__8181),
            .I(N__8178));
    Span12Mux_h I__1791 (
            .O(N__8178),
            .I(N__8175));
    Odrv12 I__1790 (
            .O(N__8175),
            .I(DRA_c_5));
    InMux I__1789 (
            .O(N__8172),
            .I(N__8169));
    LocalMux I__1788 (
            .O(N__8169),
            .I(N__8163));
    InMux I__1787 (
            .O(N__8168),
            .I(N__8160));
    InMux I__1786 (
            .O(N__8167),
            .I(N__8157));
    InMux I__1785 (
            .O(N__8166),
            .I(N__8154));
    Span4Mux_h I__1784 (
            .O(N__8163),
            .I(N__8147));
    LocalMux I__1783 (
            .O(N__8160),
            .I(N__8147));
    LocalMux I__1782 (
            .O(N__8157),
            .I(N__8147));
    LocalMux I__1781 (
            .O(N__8154),
            .I(N__8142));
    Sp12to4 I__1780 (
            .O(N__8147),
            .I(N__8142));
    Span12Mux_v I__1779 (
            .O(N__8142),
            .I(N__8139));
    Span12Mux_h I__1778 (
            .O(N__8139),
            .I(N__8136));
    Odrv12 I__1777 (
            .O(N__8136),
            .I(DRA_c_6));
    InMux I__1776 (
            .O(N__8133),
            .I(N__8127));
    InMux I__1775 (
            .O(N__8132),
            .I(N__8127));
    LocalMux I__1774 (
            .O(N__8127),
            .I(N__8124));
    Odrv4 I__1773 (
            .O(N__8124),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1772 (
            .O(N__8121),
            .I(N__8118));
    LocalMux I__1771 (
            .O(N__8118),
            .I(N__8115));
    Span4Mux_h I__1770 (
            .O(N__8115),
            .I(N__8112));
    Odrv4 I__1769 (
            .O(N__8112),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__1768 (
            .O(N__8109),
            .I(N__8106));
    LocalMux I__1767 (
            .O(N__8106),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__1766 (
            .O(N__8103),
            .I(N__8100));
    LocalMux I__1765 (
            .O(N__8100),
            .I(N__8097));
    Odrv4 I__1764 (
            .O(N__8097),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    CascadeMux I__1763 (
            .O(N__8094),
            .I(N__8091));
    InMux I__1762 (
            .O(N__8091),
            .I(N__8088));
    LocalMux I__1761 (
            .O(N__8088),
            .I(N__8085));
    Odrv4 I__1760 (
            .O(N__8085),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__1759 (
            .O(N__8082),
            .I(N__8078));
    InMux I__1758 (
            .O(N__8081),
            .I(N__8075));
    LocalMux I__1757 (
            .O(N__8078),
            .I(N__8072));
    LocalMux I__1756 (
            .O(N__8075),
            .I(N__8069));
    Span4Mux_v I__1755 (
            .O(N__8072),
            .I(N__8066));
    Span4Mux_h I__1754 (
            .O(N__8069),
            .I(N__8063));
    Sp12to4 I__1753 (
            .O(N__8066),
            .I(N__8060));
    Sp12to4 I__1752 (
            .O(N__8063),
            .I(N__8057));
    Span12Mux_h I__1751 (
            .O(N__8060),
            .I(N__8054));
    Span12Mux_v I__1750 (
            .O(N__8057),
            .I(N__8051));
    Span12Mux_v I__1749 (
            .O(N__8054),
            .I(N__8048));
    Span12Mux_h I__1748 (
            .O(N__8051),
            .I(N__8045));
    Odrv12 I__1747 (
            .O(N__8048),
            .I(DRA_c_0));
    Odrv12 I__1746 (
            .O(N__8045),
            .I(DRA_c_0));
    InMux I__1745 (
            .O(N__8040),
            .I(N__8037));
    LocalMux I__1744 (
            .O(N__8037),
            .I(N__8034));
    Span4Mux_h I__1743 (
            .O(N__8034),
            .I(N__8031));
    Odrv4 I__1742 (
            .O(N__8031),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__1741 (
            .O(N__8028),
            .I(N__8022));
    InMux I__1740 (
            .O(N__8027),
            .I(N__8022));
    LocalMux I__1739 (
            .O(N__8022),
            .I(N__8017));
    InMux I__1738 (
            .O(N__8021),
            .I(N__8012));
    InMux I__1737 (
            .O(N__8020),
            .I(N__8012));
    Span4Mux_h I__1736 (
            .O(N__8017),
            .I(N__8007));
    LocalMux I__1735 (
            .O(N__8012),
            .I(N__8007));
    Span4Mux_v I__1734 (
            .O(N__8007),
            .I(N__8004));
    Sp12to4 I__1733 (
            .O(N__8004),
            .I(N__8001));
    Span12Mux_v I__1732 (
            .O(N__8001),
            .I(N__7998));
    Span12Mux_h I__1731 (
            .O(N__7998),
            .I(N__7995));
    Odrv12 I__1730 (
            .O(N__7995),
            .I(DRA_c_1));
    InMux I__1729 (
            .O(N__7992),
            .I(N__7989));
    LocalMux I__1728 (
            .O(N__7989),
            .I(N__7986));
    Odrv4 I__1727 (
            .O(N__7986),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1726 (
            .O(N__7983),
            .I(N__7975));
    InMux I__1725 (
            .O(N__7982),
            .I(N__7975));
    InMux I__1724 (
            .O(N__7981),
            .I(N__7970));
    InMux I__1723 (
            .O(N__7980),
            .I(N__7970));
    LocalMux I__1722 (
            .O(N__7975),
            .I(N__7965));
    LocalMux I__1721 (
            .O(N__7970),
            .I(N__7965));
    Sp12to4 I__1720 (
            .O(N__7965),
            .I(N__7962));
    Span12Mux_v I__1719 (
            .O(N__7962),
            .I(N__7959));
    Span12Mux_h I__1718 (
            .O(N__7959),
            .I(N__7956));
    Odrv12 I__1717 (
            .O(N__7956),
            .I(DRA_c_2));
    InMux I__1716 (
            .O(N__7953),
            .I(N__7950));
    LocalMux I__1715 (
            .O(N__7950),
            .I(N__7947));
    Span4Mux_h I__1714 (
            .O(N__7947),
            .I(N__7944));
    Odrv4 I__1713 (
            .O(N__7944),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1712 (
            .O(N__7941),
            .I(N__7938));
    LocalMux I__1711 (
            .O(N__7938),
            .I(N__7935));
    Span4Mux_v I__1710 (
            .O(N__7935),
            .I(N__7932));
    Odrv4 I__1709 (
            .O(N__7932),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__1708 (
            .O(N__7929),
            .I(N__7926));
    LocalMux I__1707 (
            .O(N__7926),
            .I(N__7923));
    Span4Mux_v I__1706 (
            .O(N__7923),
            .I(N__7920));
    Odrv4 I__1705 (
            .O(N__7920),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    CascadeMux I__1704 (
            .O(N__7917),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10_cascade_ ));
    CascadeMux I__1703 (
            .O(N__7914),
            .I(N__7909));
    InMux I__1702 (
            .O(N__7913),
            .I(N__7905));
    InMux I__1701 (
            .O(N__7912),
            .I(N__7898));
    InMux I__1700 (
            .O(N__7909),
            .I(N__7898));
    InMux I__1699 (
            .O(N__7908),
            .I(N__7898));
    LocalMux I__1698 (
            .O(N__7905),
            .I(N__7895));
    LocalMux I__1697 (
            .O(N__7898),
            .I(N__7892));
    Span4Mux_v I__1696 (
            .O(N__7895),
            .I(N__7889));
    Span4Mux_v I__1695 (
            .O(N__7892),
            .I(N__7886));
    Span4Mux_v I__1694 (
            .O(N__7889),
            .I(N__7881));
    Span4Mux_h I__1693 (
            .O(N__7886),
            .I(N__7881));
    Span4Mux_v I__1692 (
            .O(N__7881),
            .I(N__7878));
    Span4Mux_v I__1691 (
            .O(N__7878),
            .I(N__7875));
    Odrv4 I__1690 (
            .O(N__7875),
            .I(CLK40_PLL_i));
    IoInMux I__1689 (
            .O(N__7872),
            .I(N__7867));
    IoInMux I__1688 (
            .O(N__7871),
            .I(N__7864));
    IoInMux I__1687 (
            .O(N__7870),
            .I(N__7861));
    LocalMux I__1686 (
            .O(N__7867),
            .I(N__7858));
    LocalMux I__1685 (
            .O(N__7864),
            .I(N__7855));
    LocalMux I__1684 (
            .O(N__7861),
            .I(N__7852));
    Span4Mux_s3_v I__1683 (
            .O(N__7858),
            .I(N__7849));
    Span4Mux_s3_h I__1682 (
            .O(N__7855),
            .I(N__7846));
    Span12Mux_s3_v I__1681 (
            .O(N__7852),
            .I(N__7843));
    Sp12to4 I__1680 (
            .O(N__7849),
            .I(N__7840));
    Span4Mux_h I__1679 (
            .O(N__7846),
            .I(N__7837));
    Span12Mux_v I__1678 (
            .O(N__7843),
            .I(N__7834));
    Span12Mux_h I__1677 (
            .O(N__7840),
            .I(N__7831));
    Span4Mux_h I__1676 (
            .O(N__7837),
            .I(N__7828));
    Span12Mux_h I__1675 (
            .O(N__7834),
            .I(N__7825));
    Span12Mux_v I__1674 (
            .O(N__7831),
            .I(N__7822));
    Span4Mux_h I__1673 (
            .O(N__7828),
            .I(N__7819));
    Odrv12 I__1672 (
            .O(N__7825),
            .I(CLK40_PLL_i_i));
    Odrv12 I__1671 (
            .O(N__7822),
            .I(CLK40_PLL_i_i));
    Odrv4 I__1670 (
            .O(N__7819),
            .I(CLK40_PLL_i_i));
    InMux I__1669 (
            .O(N__7812),
            .I(N__7808));
    InMux I__1668 (
            .O(N__7811),
            .I(N__7805));
    LocalMux I__1667 (
            .O(N__7808),
            .I(N__7801));
    LocalMux I__1666 (
            .O(N__7805),
            .I(N__7798));
    InMux I__1665 (
            .O(N__7804),
            .I(N__7795));
    Span4Mux_h I__1664 (
            .O(N__7801),
            .I(N__7790));
    Span4Mux_v I__1663 (
            .O(N__7798),
            .I(N__7790));
    LocalMux I__1662 (
            .O(N__7795),
            .I(N__7786));
    Span4Mux_v I__1661 (
            .O(N__7790),
            .I(N__7783));
    InMux I__1660 (
            .O(N__7789),
            .I(N__7780));
    Span4Mux_v I__1659 (
            .O(N__7786),
            .I(N__7777));
    Span4Mux_v I__1658 (
            .O(N__7783),
            .I(N__7772));
    LocalMux I__1657 (
            .O(N__7780),
            .I(N__7772));
    Sp12to4 I__1656 (
            .O(N__7777),
            .I(N__7769));
    Span4Mux_h I__1655 (
            .O(N__7772),
            .I(N__7766));
    Span12Mux_h I__1654 (
            .O(N__7769),
            .I(N__7763));
    Span4Mux_v I__1653 (
            .O(N__7766),
            .I(N__7760));
    Span12Mux_v I__1652 (
            .O(N__7763),
            .I(N__7757));
    Span4Mux_h I__1651 (
            .O(N__7760),
            .I(N__7754));
    Odrv12 I__1650 (
            .O(N__7757),
            .I(DBRn_c));
    Odrv4 I__1649 (
            .O(N__7754),
            .I(DBRn_c));
    InMux I__1648 (
            .O(N__7749),
            .I(N__7743));
    InMux I__1647 (
            .O(N__7748),
            .I(N__7740));
    InMux I__1646 (
            .O(N__7747),
            .I(N__7735));
    InMux I__1645 (
            .O(N__7746),
            .I(N__7735));
    LocalMux I__1644 (
            .O(N__7743),
            .I(N__7727));
    LocalMux I__1643 (
            .O(N__7740),
            .I(N__7724));
    LocalMux I__1642 (
            .O(N__7735),
            .I(N__7721));
    ClkMux I__1641 (
            .O(N__7734),
            .I(N__7704));
    ClkMux I__1640 (
            .O(N__7733),
            .I(N__7704));
    ClkMux I__1639 (
            .O(N__7732),
            .I(N__7704));
    ClkMux I__1638 (
            .O(N__7731),
            .I(N__7704));
    ClkMux I__1637 (
            .O(N__7730),
            .I(N__7704));
    Glb2LocalMux I__1636 (
            .O(N__7727),
            .I(N__7704));
    Glb2LocalMux I__1635 (
            .O(N__7724),
            .I(N__7704));
    Glb2LocalMux I__1634 (
            .O(N__7721),
            .I(N__7704));
    GlobalMux I__1633 (
            .O(N__7704),
            .I(N__7701));
    gio2CtrlBuf I__1632 (
            .O(N__7701),
            .I(C1_c_g));
    InMux I__1631 (
            .O(N__7698),
            .I(N__7689));
    InMux I__1630 (
            .O(N__7697),
            .I(N__7686));
    InMux I__1629 (
            .O(N__7696),
            .I(N__7682));
    InMux I__1628 (
            .O(N__7695),
            .I(N__7677));
    InMux I__1627 (
            .O(N__7694),
            .I(N__7677));
    InMux I__1626 (
            .O(N__7693),
            .I(N__7672));
    InMux I__1625 (
            .O(N__7692),
            .I(N__7672));
    LocalMux I__1624 (
            .O(N__7689),
            .I(N__7667));
    LocalMux I__1623 (
            .O(N__7686),
            .I(N__7667));
    InMux I__1622 (
            .O(N__7685),
            .I(N__7664));
    LocalMux I__1621 (
            .O(N__7682),
            .I(N__7658));
    LocalMux I__1620 (
            .O(N__7677),
            .I(N__7654));
    LocalMux I__1619 (
            .O(N__7672),
            .I(N__7647));
    Span4Mux_v I__1618 (
            .O(N__7667),
            .I(N__7647));
    LocalMux I__1617 (
            .O(N__7664),
            .I(N__7647));
    InMux I__1616 (
            .O(N__7663),
            .I(N__7644));
    InMux I__1615 (
            .O(N__7662),
            .I(N__7641));
    InMux I__1614 (
            .O(N__7661),
            .I(N__7638));
    Span4Mux_h I__1613 (
            .O(N__7658),
            .I(N__7635));
    InMux I__1612 (
            .O(N__7657),
            .I(N__7632));
    Span4Mux_v I__1611 (
            .O(N__7654),
            .I(N__7629));
    Span4Mux_h I__1610 (
            .O(N__7647),
            .I(N__7624));
    LocalMux I__1609 (
            .O(N__7644),
            .I(N__7624));
    LocalMux I__1608 (
            .O(N__7641),
            .I(N__7621));
    LocalMux I__1607 (
            .O(N__7638),
            .I(N__7618));
    Sp12to4 I__1606 (
            .O(N__7635),
            .I(N__7607));
    LocalMux I__1605 (
            .O(N__7632),
            .I(N__7607));
    Span4Mux_v I__1604 (
            .O(N__7629),
            .I(N__7602));
    Span4Mux_v I__1603 (
            .O(N__7624),
            .I(N__7602));
    Span4Mux_v I__1602 (
            .O(N__7621),
            .I(N__7597));
    Span4Mux_v I__1601 (
            .O(N__7618),
            .I(N__7597));
    InMux I__1600 (
            .O(N__7617),
            .I(N__7588));
    InMux I__1599 (
            .O(N__7616),
            .I(N__7588));
    InMux I__1598 (
            .O(N__7615),
            .I(N__7588));
    InMux I__1597 (
            .O(N__7614),
            .I(N__7588));
    InMux I__1596 (
            .O(N__7613),
            .I(N__7583));
    InMux I__1595 (
            .O(N__7612),
            .I(N__7583));
    Span12Mux_v I__1594 (
            .O(N__7607),
            .I(N__7578));
    Sp12to4 I__1593 (
            .O(N__7602),
            .I(N__7578));
    Sp12to4 I__1592 (
            .O(N__7597),
            .I(N__7571));
    LocalMux I__1591 (
            .O(N__7588),
            .I(N__7571));
    LocalMux I__1590 (
            .O(N__7583),
            .I(N__7571));
    Span12Mux_h I__1589 (
            .O(N__7578),
            .I(N__7568));
    Span12Mux_h I__1588 (
            .O(N__7571),
            .I(N__7565));
    Odrv12 I__1587 (
            .O(N__7568),
            .I(RESETn_c));
    Odrv12 I__1586 (
            .O(N__7565),
            .I(RESETn_c));
    IoInMux I__1585 (
            .O(N__7560),
            .I(N__7557));
    LocalMux I__1584 (
            .O(N__7557),
            .I(N__7554));
    Odrv12 I__1583 (
            .O(N__7554),
            .I(RESETn_c_i));
    InMux I__1582 (
            .O(N__7551),
            .I(N__7547));
    InMux I__1581 (
            .O(N__7550),
            .I(N__7544));
    LocalMux I__1580 (
            .O(N__7547),
            .I(N__7541));
    LocalMux I__1579 (
            .O(N__7544),
            .I(N__7537));
    Span4Mux_h I__1578 (
            .O(N__7541),
            .I(N__7534));
    InMux I__1577 (
            .O(N__7540),
            .I(N__7527));
    Span4Mux_v I__1576 (
            .O(N__7537),
            .I(N__7522));
    Span4Mux_v I__1575 (
            .O(N__7534),
            .I(N__7522));
    InMux I__1574 (
            .O(N__7533),
            .I(N__7517));
    InMux I__1573 (
            .O(N__7532),
            .I(N__7517));
    InMux I__1572 (
            .O(N__7531),
            .I(N__7514));
    InMux I__1571 (
            .O(N__7530),
            .I(N__7511));
    LocalMux I__1570 (
            .O(N__7527),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__1569 (
            .O(N__7522),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1568 (
            .O(N__7517),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1567 (
            .O(N__7514),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1566 (
            .O(N__7511),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__1565 (
            .O(N__7500),
            .I(N__7497));
    LocalMux I__1564 (
            .O(N__7497),
            .I(N__7494));
    IoSpan4Mux I__1563 (
            .O(N__7494),
            .I(N__7491));
    Sp12to4 I__1562 (
            .O(N__7491),
            .I(N__7488));
    Span12Mux_s7_v I__1561 (
            .O(N__7488),
            .I(N__7485));
    Odrv12 I__1560 (
            .O(N__7485),
            .I(RASn_c));
    InMux I__1559 (
            .O(N__7482),
            .I(N__7478));
    InMux I__1558 (
            .O(N__7481),
            .I(N__7475));
    LocalMux I__1557 (
            .O(N__7478),
            .I(N__7472));
    LocalMux I__1556 (
            .O(N__7475),
            .I(N__7469));
    Span4Mux_v I__1555 (
            .O(N__7472),
            .I(N__7464));
    Span4Mux_v I__1554 (
            .O(N__7469),
            .I(N__7461));
    InMux I__1553 (
            .O(N__7468),
            .I(N__7456));
    InMux I__1552 (
            .O(N__7467),
            .I(N__7456));
    Odrv4 I__1551 (
            .O(N__7464),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    Odrv4 I__1550 (
            .O(N__7461),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1549 (
            .O(N__7456),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    InMux I__1548 (
            .O(N__7449),
            .I(N__7446));
    LocalMux I__1547 (
            .O(N__7446),
            .I(N__7443));
    Span4Mux_v I__1546 (
            .O(N__7443),
            .I(N__7440));
    Span4Mux_v I__1545 (
            .O(N__7440),
            .I(N__7437));
    Sp12to4 I__1544 (
            .O(N__7437),
            .I(N__7434));
    Span12Mux_h I__1543 (
            .O(N__7434),
            .I(N__7431));
    Odrv12 I__1542 (
            .O(N__7431),
            .I(A_c_19));
    IoInMux I__1541 (
            .O(N__7428),
            .I(N__7425));
    LocalMux I__1540 (
            .O(N__7425),
            .I(N__7422));
    IoSpan4Mux I__1539 (
            .O(N__7422),
            .I(N__7419));
    IoSpan4Mux I__1538 (
            .O(N__7419),
            .I(N__7416));
    Span4Mux_s2_h I__1537 (
            .O(N__7416),
            .I(N__7413));
    Sp12to4 I__1536 (
            .O(N__7413),
            .I(N__7410));
    Odrv12 I__1535 (
            .O(N__7410),
            .I(CMA_c_9));
    CEMux I__1534 (
            .O(N__7407),
            .I(N__7404));
    LocalMux I__1533 (
            .O(N__7404),
            .I(N__7400));
    CEMux I__1532 (
            .O(N__7403),
            .I(N__7397));
    Span4Mux_v I__1531 (
            .O(N__7400),
            .I(N__7391));
    LocalMux I__1530 (
            .O(N__7397),
            .I(N__7391));
    CEMux I__1529 (
            .O(N__7396),
            .I(N__7388));
    Span4Mux_v I__1528 (
            .O(N__7391),
            .I(N__7382));
    LocalMux I__1527 (
            .O(N__7388),
            .I(N__7379));
    CEMux I__1526 (
            .O(N__7387),
            .I(N__7376));
    CEMux I__1525 (
            .O(N__7386),
            .I(N__7373));
    CEMux I__1524 (
            .O(N__7385),
            .I(N__7370));
    Odrv4 I__1523 (
            .O(N__7382),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv12 I__1522 (
            .O(N__7379),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__1521 (
            .O(N__7376),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__1520 (
            .O(N__7373),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    LocalMux I__1519 (
            .O(N__7370),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    CascadeMux I__1518 (
            .O(N__7359),
            .I(N__7353));
    CascadeMux I__1517 (
            .O(N__7358),
            .I(N__7350));
    CascadeMux I__1516 (
            .O(N__7357),
            .I(N__7343));
    CascadeMux I__1515 (
            .O(N__7356),
            .I(N__7340));
    InMux I__1514 (
            .O(N__7353),
            .I(N__7337));
    InMux I__1513 (
            .O(N__7350),
            .I(N__7333));
    InMux I__1512 (
            .O(N__7349),
            .I(N__7330));
    InMux I__1511 (
            .O(N__7348),
            .I(N__7327));
    InMux I__1510 (
            .O(N__7347),
            .I(N__7322));
    InMux I__1509 (
            .O(N__7346),
            .I(N__7322));
    InMux I__1508 (
            .O(N__7343),
            .I(N__7317));
    InMux I__1507 (
            .O(N__7340),
            .I(N__7317));
    LocalMux I__1506 (
            .O(N__7337),
            .I(N__7314));
    InMux I__1505 (
            .O(N__7336),
            .I(N__7311));
    LocalMux I__1504 (
            .O(N__7333),
            .I(N__7306));
    LocalMux I__1503 (
            .O(N__7330),
            .I(N__7306));
    LocalMux I__1502 (
            .O(N__7327),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1501 (
            .O(N__7322),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1500 (
            .O(N__7317),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__1499 (
            .O(N__7314),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__1498 (
            .O(N__7311),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv12 I__1497 (
            .O(N__7306),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    InMux I__1496 (
            .O(N__7293),
            .I(N__7290));
    LocalMux I__1495 (
            .O(N__7290),
            .I(N__7287));
    Odrv4 I__1494 (
            .O(N__7287),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    InMux I__1493 (
            .O(N__7284),
            .I(N__7281));
    LocalMux I__1492 (
            .O(N__7281),
            .I(N__7278));
    Odrv4 I__1491 (
            .O(N__7278),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__1490 (
            .O(N__7275),
            .I(N__7272));
    LocalMux I__1489 (
            .O(N__7272),
            .I(N__7269));
    Span4Mux_v I__1488 (
            .O(N__7269),
            .I(N__7266));
    Span4Mux_h I__1487 (
            .O(N__7266),
            .I(N__7262));
    InMux I__1486 (
            .O(N__7265),
            .I(N__7259));
    Odrv4 I__1485 (
            .O(N__7262),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    LocalMux I__1484 (
            .O(N__7259),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__1483 (
            .O(N__7254),
            .I(N__7251));
    LocalMux I__1482 (
            .O(N__7251),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    InMux I__1481 (
            .O(N__7248),
            .I(N__7245));
    LocalMux I__1480 (
            .O(N__7245),
            .I(N__7242));
    Odrv12 I__1479 (
            .O(N__7242),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__1478 (
            .O(N__7239),
            .I(N__7236));
    LocalMux I__1477 (
            .O(N__7236),
            .I(N__7233));
    Span4Mux_h I__1476 (
            .O(N__7233),
            .I(N__7230));
    Odrv4 I__1475 (
            .O(N__7230),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    CascadeMux I__1474 (
            .O(N__7227),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_ ));
    IoInMux I__1473 (
            .O(N__7224),
            .I(N__7221));
    LocalMux I__1472 (
            .O(N__7221),
            .I(N__7218));
    Span12Mux_s4_h I__1471 (
            .O(N__7218),
            .I(N__7215));
    Span12Mux_h I__1470 (
            .O(N__7215),
            .I(N__7212));
    Odrv12 I__1469 (
            .O(N__7212),
            .I(CMA_c_4));
    CascadeMux I__1468 (
            .O(N__7209),
            .I(N__7206));
    InMux I__1467 (
            .O(N__7206),
            .I(N__7196));
    InMux I__1466 (
            .O(N__7205),
            .I(N__7196));
    InMux I__1465 (
            .O(N__7204),
            .I(N__7196));
    InMux I__1464 (
            .O(N__7203),
            .I(N__7193));
    LocalMux I__1463 (
            .O(N__7196),
            .I(N__7188));
    LocalMux I__1462 (
            .O(N__7193),
            .I(N__7185));
    InMux I__1461 (
            .O(N__7192),
            .I(N__7180));
    InMux I__1460 (
            .O(N__7191),
            .I(N__7180));
    Odrv4 I__1459 (
            .O(N__7188),
            .I(\U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5Z0Z_1 ));
    Odrv4 I__1458 (
            .O(N__7185),
            .I(\U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5Z0Z_1 ));
    LocalMux I__1457 (
            .O(N__7180),
            .I(\U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5Z0Z_1 ));
    InMux I__1456 (
            .O(N__7173),
            .I(N__7170));
    LocalMux I__1455 (
            .O(N__7170),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1454 (
            .O(N__7167),
            .I(N__7164));
    LocalMux I__1453 (
            .O(N__7164),
            .I(N__7161));
    Span4Mux_s2_h I__1452 (
            .O(N__7161),
            .I(N__7158));
    Sp12to4 I__1451 (
            .O(N__7158),
            .I(N__7155));
    Span12Mux_v I__1450 (
            .O(N__7155),
            .I(N__7152));
    Span12Mux_h I__1449 (
            .O(N__7152),
            .I(N__7149));
    Odrv12 I__1448 (
            .O(N__7149),
            .I(CMA_c_7));
    InMux I__1447 (
            .O(N__7146),
            .I(N__7143));
    LocalMux I__1446 (
            .O(N__7143),
            .I(N__7140));
    Odrv4 I__1445 (
            .O(N__7140),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__1444 (
            .O(N__7137),
            .I(N__7134));
    LocalMux I__1443 (
            .O(N__7134),
            .I(N__7130));
    InMux I__1442 (
            .O(N__7133),
            .I(N__7127));
    Span4Mux_h I__1441 (
            .O(N__7130),
            .I(N__7124));
    LocalMux I__1440 (
            .O(N__7127),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    Odrv4 I__1439 (
            .O(N__7124),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    InMux I__1438 (
            .O(N__7119),
            .I(N__7116));
    LocalMux I__1437 (
            .O(N__7116),
            .I(N__7113));
    Span4Mux_v I__1436 (
            .O(N__7113),
            .I(N__7110));
    Span4Mux_h I__1435 (
            .O(N__7110),
            .I(N__7107));
    Odrv4 I__1434 (
            .O(N__7107),
            .I(\U712_CHIP_RAM.un5_DMA_CYCLE_START_0 ));
    InMux I__1433 (
            .O(N__7104),
            .I(N__7101));
    LocalMux I__1432 (
            .O(N__7101),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10 ));
    InMux I__1431 (
            .O(N__7098),
            .I(N__7094));
    InMux I__1430 (
            .O(N__7097),
            .I(N__7091));
    LocalMux I__1429 (
            .O(N__7094),
            .I(\U712_REG_SM.ASn_0_sqmuxa_1 ));
    LocalMux I__1428 (
            .O(N__7091),
            .I(\U712_REG_SM.ASn_0_sqmuxa_1 ));
    InMux I__1427 (
            .O(N__7086),
            .I(N__7082));
    InMux I__1426 (
            .O(N__7085),
            .I(N__7079));
    LocalMux I__1425 (
            .O(N__7082),
            .I(\U712_REG_SM.N_226 ));
    LocalMux I__1424 (
            .O(N__7079),
            .I(\U712_REG_SM.N_226 ));
    IoInMux I__1423 (
            .O(N__7074),
            .I(N__7071));
    LocalMux I__1422 (
            .O(N__7071),
            .I(N__7068));
    IoSpan4Mux I__1421 (
            .O(N__7068),
            .I(N__7065));
    Span4Mux_s1_v I__1420 (
            .O(N__7065),
            .I(N__7062));
    Span4Mux_v I__1419 (
            .O(N__7062),
            .I(N__7059));
    Sp12to4 I__1418 (
            .O(N__7059),
            .I(N__7056));
    Span12Mux_h I__1417 (
            .O(N__7056),
            .I(N__7052));
    InMux I__1416 (
            .O(N__7055),
            .I(N__7049));
    Odrv12 I__1415 (
            .O(N__7052),
            .I(ASn_c));
    LocalMux I__1414 (
            .O(N__7049),
            .I(ASn_c));
    IoInMux I__1413 (
            .O(N__7044),
            .I(N__7041));
    LocalMux I__1412 (
            .O(N__7041),
            .I(N__7038));
    Span4Mux_s2_v I__1411 (
            .O(N__7038),
            .I(N__7035));
    Span4Mux_v I__1410 (
            .O(N__7035),
            .I(N__7032));
    Odrv4 I__1409 (
            .O(N__7032),
            .I(CONSTANT_ONE_NET));
    IoInMux I__1408 (
            .O(N__7029),
            .I(N__7026));
    LocalMux I__1407 (
            .O(N__7026),
            .I(N__7023));
    Span12Mux_s8_v I__1406 (
            .O(N__7023),
            .I(N__7020));
    Odrv12 I__1405 (
            .O(N__7020),
            .I(CMA_c_10));
    IoInMux I__1404 (
            .O(N__7017),
            .I(N__7014));
    LocalMux I__1403 (
            .O(N__7014),
            .I(N__7011));
    IoSpan4Mux I__1402 (
            .O(N__7011),
            .I(N__7008));
    Span4Mux_s2_v I__1401 (
            .O(N__7008),
            .I(N__7005));
    Span4Mux_v I__1400 (
            .O(N__7005),
            .I(N__7002));
    Span4Mux_v I__1399 (
            .O(N__7002),
            .I(N__6999));
    Odrv4 I__1398 (
            .O(N__6999),
            .I(CMA_c_0));
    InMux I__1397 (
            .O(N__6996),
            .I(N__6993));
    LocalMux I__1396 (
            .O(N__6993),
            .I(N__6990));
    Span12Mux_v I__1395 (
            .O(N__6990),
            .I(N__6987));
    Span12Mux_h I__1394 (
            .O(N__6987),
            .I(N__6984));
    Odrv12 I__1393 (
            .O(N__6984),
            .I(A_c_17));
    IoInMux I__1392 (
            .O(N__6981),
            .I(N__6978));
    LocalMux I__1391 (
            .O(N__6978),
            .I(N__6975));
    IoSpan4Mux I__1390 (
            .O(N__6975),
            .I(N__6972));
    Span4Mux_s2_h I__1389 (
            .O(N__6972),
            .I(N__6969));
    Sp12to4 I__1388 (
            .O(N__6969),
            .I(N__6966));
    Span12Mux_h I__1387 (
            .O(N__6966),
            .I(N__6963));
    Odrv12 I__1386 (
            .O(N__6963),
            .I(CMA_c_8));
    InMux I__1385 (
            .O(N__6960),
            .I(N__6957));
    LocalMux I__1384 (
            .O(N__6957),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__1383 (
            .O(N__6954),
            .I(N__6951));
    LocalMux I__1382 (
            .O(N__6951),
            .I(N__6948));
    IoSpan4Mux I__1381 (
            .O(N__6948),
            .I(N__6945));
    Span4Mux_s3_h I__1380 (
            .O(N__6945),
            .I(N__6942));
    Span4Mux_h I__1379 (
            .O(N__6942),
            .I(N__6939));
    Sp12to4 I__1378 (
            .O(N__6939),
            .I(N__6936));
    Span12Mux_h I__1377 (
            .O(N__6936),
            .I(N__6933));
    Odrv12 I__1376 (
            .O(N__6933),
            .I(CMA_c_3));
    IoInMux I__1375 (
            .O(N__6930),
            .I(N__6927));
    LocalMux I__1374 (
            .O(N__6927),
            .I(N__6924));
    IoSpan4Mux I__1373 (
            .O(N__6924),
            .I(N__6921));
    Span4Mux_s3_h I__1372 (
            .O(N__6921),
            .I(N__6918));
    Span4Mux_v I__1371 (
            .O(N__6918),
            .I(N__6915));
    Span4Mux_h I__1370 (
            .O(N__6915),
            .I(N__6912));
    Sp12to4 I__1369 (
            .O(N__6912),
            .I(N__6909));
    Odrv12 I__1368 (
            .O(N__6909),
            .I(CMA_c_6));
    InMux I__1367 (
            .O(N__6906),
            .I(N__6903));
    LocalMux I__1366 (
            .O(N__6903),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__1365 (
            .O(N__6900),
            .I(N__6897));
    LocalMux I__1364 (
            .O(N__6897),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    InMux I__1363 (
            .O(N__6894),
            .I(N__6891));
    LocalMux I__1362 (
            .O(N__6891),
            .I(N__6888));
    Odrv4 I__1361 (
            .O(N__6888),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    InMux I__1360 (
            .O(N__6885),
            .I(N__6882));
    LocalMux I__1359 (
            .O(N__6882),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    IoInMux I__1358 (
            .O(N__6879),
            .I(N__6876));
    LocalMux I__1357 (
            .O(N__6876),
            .I(N__6873));
    IoSpan4Mux I__1356 (
            .O(N__6873),
            .I(N__6870));
    Span4Mux_s3_h I__1355 (
            .O(N__6870),
            .I(N__6867));
    Sp12to4 I__1354 (
            .O(N__6867),
            .I(N__6864));
    Span12Mux_h I__1353 (
            .O(N__6864),
            .I(N__6861));
    Odrv12 I__1352 (
            .O(N__6861),
            .I(CMA_c_5));
    InMux I__1351 (
            .O(N__6858),
            .I(N__6855));
    LocalMux I__1350 (
            .O(N__6855),
            .I(N__6852));
    Span4Mux_v I__1349 (
            .O(N__6852),
            .I(N__6849));
    Sp12to4 I__1348 (
            .O(N__6849),
            .I(N__6846));
    Span12Mux_h I__1347 (
            .O(N__6846),
            .I(N__6843));
    Odrv12 I__1346 (
            .O(N__6843),
            .I(A_c_9));
    InMux I__1345 (
            .O(N__6840),
            .I(N__6837));
    LocalMux I__1344 (
            .O(N__6837),
            .I(N__6834));
    Span4Mux_v I__1343 (
            .O(N__6834),
            .I(N__6831));
    Sp12to4 I__1342 (
            .O(N__6831),
            .I(N__6828));
    Span12Mux_v I__1341 (
            .O(N__6828),
            .I(N__6825));
    Span12Mux_h I__1340 (
            .O(N__6825),
            .I(N__6822));
    Odrv12 I__1339 (
            .O(N__6822),
            .I(A_c_2));
    InMux I__1338 (
            .O(N__6819),
            .I(N__6816));
    LocalMux I__1337 (
            .O(N__6816),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__1336 (
            .O(N__6813),
            .I(N__6810));
    LocalMux I__1335 (
            .O(N__6810),
            .I(N__6807));
    Span4Mux_v I__1334 (
            .O(N__6807),
            .I(N__6804));
    Sp12to4 I__1333 (
            .O(N__6804),
            .I(N__6801));
    Span12Mux_h I__1332 (
            .O(N__6801),
            .I(N__6798));
    Odrv12 I__1331 (
            .O(N__6798),
            .I(A_c_10));
    InMux I__1330 (
            .O(N__6795),
            .I(N__6792));
    LocalMux I__1329 (
            .O(N__6792),
            .I(N__6789));
    Span12Mux_h I__1328 (
            .O(N__6789),
            .I(N__6786));
    Span12Mux_v I__1327 (
            .O(N__6786),
            .I(N__6783));
    Odrv12 I__1326 (
            .O(N__6783),
            .I(A_c_3));
    CascadeMux I__1325 (
            .O(N__6780),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ));
    InMux I__1324 (
            .O(N__6777),
            .I(N__6774));
    LocalMux I__1323 (
            .O(N__6774),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    CascadeMux I__1322 (
            .O(N__6771),
            .I(N__6768));
    InMux I__1321 (
            .O(N__6768),
            .I(N__6762));
    InMux I__1320 (
            .O(N__6767),
            .I(N__6762));
    LocalMux I__1319 (
            .O(N__6762),
            .I(N__6759));
    Span4Mux_v I__1318 (
            .O(N__6759),
            .I(N__6756));
    Span4Mux_v I__1317 (
            .O(N__6756),
            .I(N__6753));
    Sp12to4 I__1316 (
            .O(N__6753),
            .I(N__6750));
    Span12Mux_h I__1315 (
            .O(N__6750),
            .I(N__6747));
    Odrv12 I__1314 (
            .O(N__6747),
            .I(A_c_14));
    InMux I__1313 (
            .O(N__6744),
            .I(N__6741));
    LocalMux I__1312 (
            .O(N__6741),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__1311 (
            .O(N__6738),
            .I(N__6733));
    InMux I__1310 (
            .O(N__6737),
            .I(N__6728));
    InMux I__1309 (
            .O(N__6736),
            .I(N__6728));
    LocalMux I__1308 (
            .O(N__6733),
            .I(N__6725));
    LocalMux I__1307 (
            .O(N__6728),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    Odrv4 I__1306 (
            .O(N__6725),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__1305 (
            .O(N__6720),
            .I(N__6716));
    InMux I__1304 (
            .O(N__6719),
            .I(N__6713));
    LocalMux I__1303 (
            .O(N__6716),
            .I(N__6710));
    LocalMux I__1302 (
            .O(N__6713),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    Odrv12 I__1301 (
            .O(N__6710),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__1300 (
            .O(N__6705),
            .I(N__6702));
    LocalMux I__1299 (
            .O(N__6702),
            .I(N__6699));
    Odrv12 I__1298 (
            .O(N__6699),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ));
    InMux I__1297 (
            .O(N__6696),
            .I(N__6687));
    InMux I__1296 (
            .O(N__6695),
            .I(N__6680));
    InMux I__1295 (
            .O(N__6694),
            .I(N__6680));
    InMux I__1294 (
            .O(N__6693),
            .I(N__6680));
    InMux I__1293 (
            .O(N__6692),
            .I(N__6677));
    InMux I__1292 (
            .O(N__6691),
            .I(N__6672));
    InMux I__1291 (
            .O(N__6690),
            .I(N__6672));
    LocalMux I__1290 (
            .O(N__6687),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__1289 (
            .O(N__6680),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__1288 (
            .O(N__6677),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    LocalMux I__1287 (
            .O(N__6672),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    CascadeMux I__1286 (
            .O(N__6663),
            .I(N__6659));
    CascadeMux I__1285 (
            .O(N__6662),
            .I(N__6654));
    InMux I__1284 (
            .O(N__6659),
            .I(N__6648));
    InMux I__1283 (
            .O(N__6658),
            .I(N__6648));
    InMux I__1282 (
            .O(N__6657),
            .I(N__6645));
    InMux I__1281 (
            .O(N__6654),
            .I(N__6642));
    InMux I__1280 (
            .O(N__6653),
            .I(N__6639));
    LocalMux I__1279 (
            .O(N__6648),
            .I(N__6636));
    LocalMux I__1278 (
            .O(N__6645),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1277 (
            .O(N__6642),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1276 (
            .O(N__6639),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    Odrv4 I__1275 (
            .O(N__6636),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    CascadeMux I__1274 (
            .O(N__6627),
            .I(N__6619));
    CascadeMux I__1273 (
            .O(N__6626),
            .I(N__6616));
    InMux I__1272 (
            .O(N__6625),
            .I(N__6613));
    InMux I__1271 (
            .O(N__6624),
            .I(N__6608));
    InMux I__1270 (
            .O(N__6623),
            .I(N__6608));
    InMux I__1269 (
            .O(N__6622),
            .I(N__6605));
    InMux I__1268 (
            .O(N__6619),
            .I(N__6600));
    InMux I__1267 (
            .O(N__6616),
            .I(N__6600));
    LocalMux I__1266 (
            .O(N__6613),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1265 (
            .O(N__6608),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1264 (
            .O(N__6605),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1263 (
            .O(N__6600),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__1262 (
            .O(N__6591),
            .I(N__6581));
    InMux I__1261 (
            .O(N__6590),
            .I(N__6576));
    InMux I__1260 (
            .O(N__6589),
            .I(N__6576));
    InMux I__1259 (
            .O(N__6588),
            .I(N__6573));
    InMux I__1258 (
            .O(N__6587),
            .I(N__6564));
    InMux I__1257 (
            .O(N__6586),
            .I(N__6564));
    InMux I__1256 (
            .O(N__6585),
            .I(N__6564));
    InMux I__1255 (
            .O(N__6584),
            .I(N__6564));
    LocalMux I__1254 (
            .O(N__6581),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__1253 (
            .O(N__6576),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__1252 (
            .O(N__6573),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__1251 (
            .O(N__6564),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    CascadeMux I__1250 (
            .O(N__6555),
            .I(N__6551));
    InMux I__1249 (
            .O(N__6554),
            .I(N__6544));
    InMux I__1248 (
            .O(N__6551),
            .I(N__6541));
    InMux I__1247 (
            .O(N__6550),
            .I(N__6536));
    InMux I__1246 (
            .O(N__6549),
            .I(N__6536));
    InMux I__1245 (
            .O(N__6548),
            .I(N__6531));
    InMux I__1244 (
            .O(N__6547),
            .I(N__6531));
    LocalMux I__1243 (
            .O(N__6544),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1242 (
            .O(N__6541),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1241 (
            .O(N__6536),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1240 (
            .O(N__6531),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    InMux I__1239 (
            .O(N__6522),
            .I(N__6519));
    LocalMux I__1238 (
            .O(N__6519),
            .I(\U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0 ));
    CascadeMux I__1237 (
            .O(N__6516),
            .I(N__6513));
    InMux I__1236 (
            .O(N__6513),
            .I(N__6510));
    LocalMux I__1235 (
            .O(N__6510),
            .I(N__6507));
    Odrv4 I__1234 (
            .O(N__6507),
            .I(\U712_REG_SM.DS_EN_RNOZ0Z_0 ));
    InMux I__1233 (
            .O(N__6504),
            .I(N__6501));
    LocalMux I__1232 (
            .O(N__6501),
            .I(\U712_REG_SM.N_300 ));
    InMux I__1231 (
            .O(N__6498),
            .I(N__6494));
    InMux I__1230 (
            .O(N__6497),
            .I(N__6491));
    LocalMux I__1229 (
            .O(N__6494),
            .I(\U712_REG_SM.N_228 ));
    LocalMux I__1228 (
            .O(N__6491),
            .I(\U712_REG_SM.N_228 ));
    InMux I__1227 (
            .O(N__6486),
            .I(N__6483));
    LocalMux I__1226 (
            .O(N__6483),
            .I(N__6480));
    Span4Mux_h I__1225 (
            .O(N__6480),
            .I(N__6476));
    InMux I__1224 (
            .O(N__6479),
            .I(N__6473));
    Odrv4 I__1223 (
            .O(N__6476),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__1222 (
            .O(N__6473),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    IoInMux I__1221 (
            .O(N__6468),
            .I(N__6465));
    LocalMux I__1220 (
            .O(N__6465),
            .I(N__6461));
    InMux I__1219 (
            .O(N__6464),
            .I(N__6457));
    Span12Mux_s2_v I__1218 (
            .O(N__6461),
            .I(N__6454));
    CascadeMux I__1217 (
            .O(N__6460),
            .I(N__6451));
    LocalMux I__1216 (
            .O(N__6457),
            .I(N__6448));
    Span12Mux_v I__1215 (
            .O(N__6454),
            .I(N__6445));
    InMux I__1214 (
            .O(N__6451),
            .I(N__6442));
    Span4Mux_v I__1213 (
            .O(N__6448),
            .I(N__6439));
    Odrv12 I__1212 (
            .O(N__6445),
            .I(REGENn_c));
    LocalMux I__1211 (
            .O(N__6442),
            .I(REGENn_c));
    Odrv4 I__1210 (
            .O(N__6439),
            .I(REGENn_c));
    InMux I__1209 (
            .O(N__6432),
            .I(N__6429));
    LocalMux I__1208 (
            .O(N__6429),
            .I(N__6426));
    Odrv4 I__1207 (
            .O(N__6426),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__1206 (
            .O(N__6423),
            .I(N__6420));
    LocalMux I__1205 (
            .O(N__6420),
            .I(N__6417));
    Span12Mux_s9_v I__1204 (
            .O(N__6417),
            .I(N__6414));
    Odrv12 I__1203 (
            .O(N__6414),
            .I(CMA_c_2));
    InMux I__1202 (
            .O(N__6411),
            .I(N__6408));
    LocalMux I__1201 (
            .O(N__6408),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i ));
    InMux I__1200 (
            .O(N__6405),
            .I(N__6402));
    LocalMux I__1199 (
            .O(N__6402),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    InMux I__1198 (
            .O(N__6399),
            .I(N__6396));
    LocalMux I__1197 (
            .O(N__6396),
            .I(N__6393));
    Span4Mux_h I__1196 (
            .O(N__6393),
            .I(N__6390));
    Odrv4 I__1195 (
            .O(N__6390),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    IoInMux I__1194 (
            .O(N__6387),
            .I(N__6384));
    LocalMux I__1193 (
            .O(N__6384),
            .I(N__6381));
    Span4Mux_s3_v I__1192 (
            .O(N__6381),
            .I(N__6378));
    Span4Mux_v I__1191 (
            .O(N__6378),
            .I(N__6375));
    Odrv4 I__1190 (
            .O(N__6375),
            .I(CMA_c_1));
    InMux I__1189 (
            .O(N__6372),
            .I(N__6359));
    InMux I__1188 (
            .O(N__6371),
            .I(N__6359));
    InMux I__1187 (
            .O(N__6370),
            .I(N__6359));
    InMux I__1186 (
            .O(N__6369),
            .I(N__6356));
    InMux I__1185 (
            .O(N__6368),
            .I(N__6349));
    InMux I__1184 (
            .O(N__6367),
            .I(N__6349));
    InMux I__1183 (
            .O(N__6366),
            .I(N__6349));
    LocalMux I__1182 (
            .O(N__6359),
            .I(\U712_CHIP_RAM.N_36 ));
    LocalMux I__1181 (
            .O(N__6356),
            .I(\U712_CHIP_RAM.N_36 ));
    LocalMux I__1180 (
            .O(N__6349),
            .I(\U712_CHIP_RAM.N_36 ));
    InMux I__1179 (
            .O(N__6342),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    InMux I__1178 (
            .O(N__6339),
            .I(N__6335));
    InMux I__1177 (
            .O(N__6338),
            .I(N__6332));
    LocalMux I__1176 (
            .O(N__6335),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1175 (
            .O(N__6332),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    CEMux I__1174 (
            .O(N__6327),
            .I(N__6324));
    LocalMux I__1173 (
            .O(N__6324),
            .I(N__6320));
    CEMux I__1172 (
            .O(N__6323),
            .I(N__6317));
    Span4Mux_v I__1171 (
            .O(N__6320),
            .I(N__6314));
    LocalMux I__1170 (
            .O(N__6317),
            .I(N__6311));
    Span4Mux_h I__1169 (
            .O(N__6314),
            .I(N__6306));
    Span4Mux_v I__1168 (
            .O(N__6311),
            .I(N__6306));
    Span4Mux_h I__1167 (
            .O(N__6306),
            .I(N__6303));
    Odrv4 I__1166 (
            .O(N__6303),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__1165 (
            .O(N__6300),
            .I(N__6297));
    LocalMux I__1164 (
            .O(N__6297),
            .I(N__6294));
    Odrv4 I__1163 (
            .O(N__6294),
            .I(\U712_CHIP_RAM.N_285 ));
    InMux I__1162 (
            .O(N__6291),
            .I(N__6285));
    InMux I__1161 (
            .O(N__6290),
            .I(N__6282));
    InMux I__1160 (
            .O(N__6289),
            .I(N__6277));
    InMux I__1159 (
            .O(N__6288),
            .I(N__6277));
    LocalMux I__1158 (
            .O(N__6285),
            .I(N__6271));
    LocalMux I__1157 (
            .O(N__6282),
            .I(N__6271));
    LocalMux I__1156 (
            .O(N__6277),
            .I(N__6268));
    InMux I__1155 (
            .O(N__6276),
            .I(N__6265));
    Odrv4 I__1154 (
            .O(N__6271),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__1153 (
            .O(N__6268),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1152 (
            .O(N__6265),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    CascadeMux I__1151 (
            .O(N__6258),
            .I(N__6253));
    InMux I__1150 (
            .O(N__6257),
            .I(N__6243));
    InMux I__1149 (
            .O(N__6256),
            .I(N__6243));
    InMux I__1148 (
            .O(N__6253),
            .I(N__6243));
    CascadeMux I__1147 (
            .O(N__6252),
            .I(N__6238));
    InMux I__1146 (
            .O(N__6251),
            .I(N__6233));
    InMux I__1145 (
            .O(N__6250),
            .I(N__6233));
    LocalMux I__1144 (
            .O(N__6243),
            .I(N__6230));
    CascadeMux I__1143 (
            .O(N__6242),
            .I(N__6227));
    InMux I__1142 (
            .O(N__6241),
            .I(N__6221));
    InMux I__1141 (
            .O(N__6238),
            .I(N__6221));
    LocalMux I__1140 (
            .O(N__6233),
            .I(N__6218));
    Span4Mux_v I__1139 (
            .O(N__6230),
            .I(N__6215));
    InMux I__1138 (
            .O(N__6227),
            .I(N__6210));
    InMux I__1137 (
            .O(N__6226),
            .I(N__6210));
    LocalMux I__1136 (
            .O(N__6221),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1135 (
            .O(N__6218),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1134 (
            .O(N__6215),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1133 (
            .O(N__6210),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1132 (
            .O(N__6201),
            .I(N__6198));
    LocalMux I__1131 (
            .O(N__6198),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_a3_0_a3_0 ));
    InMux I__1130 (
            .O(N__6195),
            .I(N__6192));
    LocalMux I__1129 (
            .O(N__6192),
            .I(N__6189));
    Span4Mux_v I__1128 (
            .O(N__6189),
            .I(N__6185));
    InMux I__1127 (
            .O(N__6188),
            .I(N__6182));
    Odrv4 I__1126 (
            .O(N__6185),
            .I(\U712_CHIP_RAM.N_342 ));
    LocalMux I__1125 (
            .O(N__6182),
            .I(\U712_CHIP_RAM.N_342 ));
    InMux I__1124 (
            .O(N__6177),
            .I(N__6174));
    LocalMux I__1123 (
            .O(N__6174),
            .I(N__6171));
    Span4Mux_v I__1122 (
            .O(N__6171),
            .I(N__6165));
    InMux I__1121 (
            .O(N__6170),
            .I(N__6162));
    InMux I__1120 (
            .O(N__6169),
            .I(N__6157));
    InMux I__1119 (
            .O(N__6168),
            .I(N__6157));
    Odrv4 I__1118 (
            .O(N__6165),
            .I(\U712_CHIP_RAM.N_328 ));
    LocalMux I__1117 (
            .O(N__6162),
            .I(\U712_CHIP_RAM.N_328 ));
    LocalMux I__1116 (
            .O(N__6157),
            .I(\U712_CHIP_RAM.N_328 ));
    CascadeMux I__1115 (
            .O(N__6150),
            .I(N__6146));
    CascadeMux I__1114 (
            .O(N__6149),
            .I(N__6143));
    InMux I__1113 (
            .O(N__6146),
            .I(N__6137));
    InMux I__1112 (
            .O(N__6143),
            .I(N__6137));
    InMux I__1111 (
            .O(N__6142),
            .I(N__6129));
    LocalMux I__1110 (
            .O(N__6137),
            .I(N__6126));
    InMux I__1109 (
            .O(N__6136),
            .I(N__6123));
    InMux I__1108 (
            .O(N__6135),
            .I(N__6119));
    CascadeMux I__1107 (
            .O(N__6134),
            .I(N__6114));
    InMux I__1106 (
            .O(N__6133),
            .I(N__6111));
    InMux I__1105 (
            .O(N__6132),
            .I(N__6103));
    LocalMux I__1104 (
            .O(N__6129),
            .I(N__6096));
    Span4Mux_h I__1103 (
            .O(N__6126),
            .I(N__6096));
    LocalMux I__1102 (
            .O(N__6123),
            .I(N__6096));
    CascadeMux I__1101 (
            .O(N__6122),
            .I(N__6092));
    LocalMux I__1100 (
            .O(N__6119),
            .I(N__6087));
    InMux I__1099 (
            .O(N__6118),
            .I(N__6084));
    InMux I__1098 (
            .O(N__6117),
            .I(N__6078));
    InMux I__1097 (
            .O(N__6114),
            .I(N__6078));
    LocalMux I__1096 (
            .O(N__6111),
            .I(N__6075));
    InMux I__1095 (
            .O(N__6110),
            .I(N__6070));
    InMux I__1094 (
            .O(N__6109),
            .I(N__6070));
    InMux I__1093 (
            .O(N__6108),
            .I(N__6063));
    InMux I__1092 (
            .O(N__6107),
            .I(N__6063));
    InMux I__1091 (
            .O(N__6106),
            .I(N__6063));
    LocalMux I__1090 (
            .O(N__6103),
            .I(N__6060));
    Span4Mux_v I__1089 (
            .O(N__6096),
            .I(N__6057));
    InMux I__1088 (
            .O(N__6095),
            .I(N__6048));
    InMux I__1087 (
            .O(N__6092),
            .I(N__6048));
    InMux I__1086 (
            .O(N__6091),
            .I(N__6048));
    InMux I__1085 (
            .O(N__6090),
            .I(N__6048));
    Span4Mux_v I__1084 (
            .O(N__6087),
            .I(N__6043));
    LocalMux I__1083 (
            .O(N__6084),
            .I(N__6043));
    InMux I__1082 (
            .O(N__6083),
            .I(N__6040));
    LocalMux I__1081 (
            .O(N__6078),
            .I(N__6037));
    Span4Mux_h I__1080 (
            .O(N__6075),
            .I(N__6030));
    LocalMux I__1079 (
            .O(N__6070),
            .I(N__6030));
    LocalMux I__1078 (
            .O(N__6063),
            .I(N__6030));
    Odrv12 I__1077 (
            .O(N__6060),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1076 (
            .O(N__6057),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1075 (
            .O(N__6048),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1074 (
            .O(N__6043),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1073 (
            .O(N__6040),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1072 (
            .O(N__6037),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1071 (
            .O(N__6030),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__1070 (
            .O(N__6015),
            .I(N__6008));
    CascadeMux I__1069 (
            .O(N__6014),
            .I(N__6004));
    CascadeMux I__1068 (
            .O(N__6013),
            .I(N__6001));
    InMux I__1067 (
            .O(N__6012),
            .I(N__5994));
    InMux I__1066 (
            .O(N__6011),
            .I(N__5994));
    InMux I__1065 (
            .O(N__6008),
            .I(N__5991));
    InMux I__1064 (
            .O(N__6007),
            .I(N__5988));
    InMux I__1063 (
            .O(N__6004),
            .I(N__5985));
    InMux I__1062 (
            .O(N__6001),
            .I(N__5982));
    CascadeMux I__1061 (
            .O(N__6000),
            .I(N__5975));
    CascadeMux I__1060 (
            .O(N__5999),
            .I(N__5972));
    LocalMux I__1059 (
            .O(N__5994),
            .I(N__5963));
    LocalMux I__1058 (
            .O(N__5991),
            .I(N__5963));
    LocalMux I__1057 (
            .O(N__5988),
            .I(N__5963));
    LocalMux I__1056 (
            .O(N__5985),
            .I(N__5960));
    LocalMux I__1055 (
            .O(N__5982),
            .I(N__5957));
    InMux I__1054 (
            .O(N__5981),
            .I(N__5954));
    InMux I__1053 (
            .O(N__5980),
            .I(N__5951));
    InMux I__1052 (
            .O(N__5979),
            .I(N__5948));
    InMux I__1051 (
            .O(N__5978),
            .I(N__5941));
    InMux I__1050 (
            .O(N__5975),
            .I(N__5941));
    InMux I__1049 (
            .O(N__5972),
            .I(N__5941));
    InMux I__1048 (
            .O(N__5971),
            .I(N__5936));
    InMux I__1047 (
            .O(N__5970),
            .I(N__5936));
    Span4Mux_v I__1046 (
            .O(N__5963),
            .I(N__5933));
    Odrv4 I__1045 (
            .O(N__5960),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1044 (
            .O(N__5957),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1043 (
            .O(N__5954),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1042 (
            .O(N__5951),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1041 (
            .O(N__5948),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1040 (
            .O(N__5941),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1039 (
            .O(N__5936),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1038 (
            .O(N__5933),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1037 (
            .O(N__5916),
            .I(N__5908));
    InMux I__1036 (
            .O(N__5915),
            .I(N__5908));
    CascadeMux I__1035 (
            .O(N__5914),
            .I(N__5900));
    InMux I__1034 (
            .O(N__5913),
            .I(N__5895));
    LocalMux I__1033 (
            .O(N__5908),
            .I(N__5891));
    CascadeMux I__1032 (
            .O(N__5907),
            .I(N__5887));
    InMux I__1031 (
            .O(N__5906),
            .I(N__5883));
    InMux I__1030 (
            .O(N__5905),
            .I(N__5878));
    InMux I__1029 (
            .O(N__5904),
            .I(N__5878));
    InMux I__1028 (
            .O(N__5903),
            .I(N__5873));
    InMux I__1027 (
            .O(N__5900),
            .I(N__5873));
    CascadeMux I__1026 (
            .O(N__5899),
            .I(N__5870));
    InMux I__1025 (
            .O(N__5898),
            .I(N__5865));
    LocalMux I__1024 (
            .O(N__5895),
            .I(N__5862));
    InMux I__1023 (
            .O(N__5894),
            .I(N__5859));
    Span4Mux_v I__1022 (
            .O(N__5891),
            .I(N__5856));
    InMux I__1021 (
            .O(N__5890),
            .I(N__5849));
    InMux I__1020 (
            .O(N__5887),
            .I(N__5849));
    InMux I__1019 (
            .O(N__5886),
            .I(N__5849));
    LocalMux I__1018 (
            .O(N__5883),
            .I(N__5842));
    LocalMux I__1017 (
            .O(N__5878),
            .I(N__5842));
    LocalMux I__1016 (
            .O(N__5873),
            .I(N__5842));
    InMux I__1015 (
            .O(N__5870),
            .I(N__5835));
    InMux I__1014 (
            .O(N__5869),
            .I(N__5835));
    InMux I__1013 (
            .O(N__5868),
            .I(N__5835));
    LocalMux I__1012 (
            .O(N__5865),
            .I(N__5830));
    Span4Mux_h I__1011 (
            .O(N__5862),
            .I(N__5830));
    LocalMux I__1010 (
            .O(N__5859),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1009 (
            .O(N__5856),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1008 (
            .O(N__5849),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1007 (
            .O(N__5842),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1006 (
            .O(N__5835),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1005 (
            .O(N__5830),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__1004 (
            .O(N__5817),
            .I(N__5806));
    InMux I__1003 (
            .O(N__5816),
            .I(N__5806));
    InMux I__1002 (
            .O(N__5815),
            .I(N__5801));
    InMux I__1001 (
            .O(N__5814),
            .I(N__5801));
    InMux I__1000 (
            .O(N__5813),
            .I(N__5798));
    InMux I__999 (
            .O(N__5812),
            .I(N__5795));
    InMux I__998 (
            .O(N__5811),
            .I(N__5784));
    LocalMux I__997 (
            .O(N__5806),
            .I(N__5778));
    LocalMux I__996 (
            .O(N__5801),
            .I(N__5775));
    LocalMux I__995 (
            .O(N__5798),
            .I(N__5771));
    LocalMux I__994 (
            .O(N__5795),
            .I(N__5768));
    InMux I__993 (
            .O(N__5794),
            .I(N__5765));
    InMux I__992 (
            .O(N__5793),
            .I(N__5758));
    InMux I__991 (
            .O(N__5792),
            .I(N__5758));
    InMux I__990 (
            .O(N__5791),
            .I(N__5758));
    InMux I__989 (
            .O(N__5790),
            .I(N__5753));
    InMux I__988 (
            .O(N__5789),
            .I(N__5753));
    InMux I__987 (
            .O(N__5788),
            .I(N__5748));
    InMux I__986 (
            .O(N__5787),
            .I(N__5748));
    LocalMux I__985 (
            .O(N__5784),
            .I(N__5745));
    InMux I__984 (
            .O(N__5783),
            .I(N__5738));
    InMux I__983 (
            .O(N__5782),
            .I(N__5738));
    InMux I__982 (
            .O(N__5781),
            .I(N__5738));
    Span4Mux_v I__981 (
            .O(N__5778),
            .I(N__5733));
    Span4Mux_h I__980 (
            .O(N__5775),
            .I(N__5733));
    InMux I__979 (
            .O(N__5774),
            .I(N__5730));
    Odrv4 I__978 (
            .O(N__5771),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__977 (
            .O(N__5768),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__976 (
            .O(N__5765),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__975 (
            .O(N__5758),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__974 (
            .O(N__5753),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__973 (
            .O(N__5748),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__972 (
            .O(N__5745),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__971 (
            .O(N__5738),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__970 (
            .O(N__5733),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__969 (
            .O(N__5730),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__968 (
            .O(N__5709),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_2_i_1_cascade_ ));
    InMux I__967 (
            .O(N__5706),
            .I(N__5702));
    InMux I__966 (
            .O(N__5705),
            .I(N__5691));
    LocalMux I__965 (
            .O(N__5702),
            .I(N__5688));
    InMux I__964 (
            .O(N__5701),
            .I(N__5685));
    InMux I__963 (
            .O(N__5700),
            .I(N__5682));
    InMux I__962 (
            .O(N__5699),
            .I(N__5677));
    InMux I__961 (
            .O(N__5698),
            .I(N__5677));
    InMux I__960 (
            .O(N__5697),
            .I(N__5672));
    InMux I__959 (
            .O(N__5696),
            .I(N__5672));
    InMux I__958 (
            .O(N__5695),
            .I(N__5663));
    InMux I__957 (
            .O(N__5694),
            .I(N__5660));
    LocalMux I__956 (
            .O(N__5691),
            .I(N__5655));
    Span4Mux_h I__955 (
            .O(N__5688),
            .I(N__5655));
    LocalMux I__954 (
            .O(N__5685),
            .I(N__5652));
    LocalMux I__953 (
            .O(N__5682),
            .I(N__5645));
    LocalMux I__952 (
            .O(N__5677),
            .I(N__5645));
    LocalMux I__951 (
            .O(N__5672),
            .I(N__5645));
    InMux I__950 (
            .O(N__5671),
            .I(N__5638));
    InMux I__949 (
            .O(N__5670),
            .I(N__5638));
    InMux I__948 (
            .O(N__5669),
            .I(N__5638));
    InMux I__947 (
            .O(N__5668),
            .I(N__5633));
    InMux I__946 (
            .O(N__5667),
            .I(N__5633));
    InMux I__945 (
            .O(N__5666),
            .I(N__5630));
    LocalMux I__944 (
            .O(N__5663),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__943 (
            .O(N__5660),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__942 (
            .O(N__5655),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__941 (
            .O(N__5652),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__940 (
            .O(N__5645),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__939 (
            .O(N__5638),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__938 (
            .O(N__5633),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__937 (
            .O(N__5630),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    CascadeMux I__936 (
            .O(N__5613),
            .I(N__5610));
    InMux I__935 (
            .O(N__5610),
            .I(N__5607));
    LocalMux I__934 (
            .O(N__5607),
            .I(N__5604));
    Span4Mux_h I__933 (
            .O(N__5604),
            .I(N__5601));
    Odrv4 I__932 (
            .O(N__5601),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_2_i_2 ));
    InMux I__931 (
            .O(N__5598),
            .I(N__5593));
    InMux I__930 (
            .O(N__5597),
            .I(N__5588));
    InMux I__929 (
            .O(N__5596),
            .I(N__5588));
    LocalMux I__928 (
            .O(N__5593),
            .I(\U712_REG_SM.N_210 ));
    LocalMux I__927 (
            .O(N__5588),
            .I(\U712_REG_SM.N_210 ));
    InMux I__926 (
            .O(N__5583),
            .I(N__5577));
    InMux I__925 (
            .O(N__5582),
            .I(N__5570));
    InMux I__924 (
            .O(N__5581),
            .I(N__5570));
    InMux I__923 (
            .O(N__5580),
            .I(N__5570));
    LocalMux I__922 (
            .O(N__5577),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__921 (
            .O(N__5570),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    CascadeMux I__920 (
            .O(N__5565),
            .I(\U712_REG_SM.N_248_cascade_ ));
    InMux I__919 (
            .O(N__5562),
            .I(N__5555));
    InMux I__918 (
            .O(N__5561),
            .I(N__5552));
    InMux I__917 (
            .O(N__5560),
            .I(N__5549));
    InMux I__916 (
            .O(N__5559),
            .I(N__5544));
    InMux I__915 (
            .O(N__5558),
            .I(N__5544));
    LocalMux I__914 (
            .O(N__5555),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__913 (
            .O(N__5552),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__912 (
            .O(N__5549),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__911 (
            .O(N__5544),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__910 (
            .O(N__5535),
            .I(N__5532));
    LocalMux I__909 (
            .O(N__5532),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_1_0 ));
    InMux I__908 (
            .O(N__5529),
            .I(N__5526));
    LocalMux I__907 (
            .O(N__5526),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    InMux I__906 (
            .O(N__5523),
            .I(bfn_10_8_0_));
    InMux I__905 (
            .O(N__5520),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__904 (
            .O(N__5517),
            .I(N__5514));
    LocalMux I__903 (
            .O(N__5514),
            .I(N__5511));
    Odrv4 I__902 (
            .O(N__5511),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__901 (
            .O(N__5508),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__900 (
            .O(N__5505),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    CascadeMux I__899 (
            .O(N__5502),
            .I(N__5498));
    InMux I__898 (
            .O(N__5501),
            .I(N__5495));
    InMux I__897 (
            .O(N__5498),
            .I(N__5492));
    LocalMux I__896 (
            .O(N__5495),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__895 (
            .O(N__5492),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__894 (
            .O(N__5487),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__893 (
            .O(N__5484),
            .I(N__5480));
    InMux I__892 (
            .O(N__5483),
            .I(N__5477));
    LocalMux I__891 (
            .O(N__5480),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__890 (
            .O(N__5477),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__889 (
            .O(N__5472),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__888 (
            .O(N__5469),
            .I(N__5465));
    InMux I__887 (
            .O(N__5468),
            .I(N__5462));
    LocalMux I__886 (
            .O(N__5465),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__885 (
            .O(N__5462),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__884 (
            .O(N__5457),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__883 (
            .O(N__5454),
            .I(N__5450));
    InMux I__882 (
            .O(N__5453),
            .I(N__5447));
    LocalMux I__881 (
            .O(N__5450),
            .I(\U712_CHIP_RAM.N_211 ));
    LocalMux I__880 (
            .O(N__5447),
            .I(\U712_CHIP_RAM.N_211 ));
    InMux I__879 (
            .O(N__5442),
            .I(N__5439));
    LocalMux I__878 (
            .O(N__5439),
            .I(N__5436));
    Odrv4 I__877 (
            .O(N__5436),
            .I(\U712_CHIP_RAM.N_64_1 ));
    InMux I__876 (
            .O(N__5433),
            .I(N__5426));
    InMux I__875 (
            .O(N__5432),
            .I(N__5426));
    InMux I__874 (
            .O(N__5431),
            .I(N__5423));
    LocalMux I__873 (
            .O(N__5426),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ));
    LocalMux I__872 (
            .O(N__5423),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ));
    CascadeMux I__871 (
            .O(N__5418),
            .I(\U712_CHIP_RAM.N_64_1_cascade_ ));
    CascadeMux I__870 (
            .O(N__5415),
            .I(N__5411));
    InMux I__869 (
            .O(N__5414),
            .I(N__5407));
    InMux I__868 (
            .O(N__5411),
            .I(N__5404));
    InMux I__867 (
            .O(N__5410),
            .I(N__5401));
    LocalMux I__866 (
            .O(N__5407),
            .I(N__5396));
    LocalMux I__865 (
            .O(N__5404),
            .I(N__5396));
    LocalMux I__864 (
            .O(N__5401),
            .I(\U712_CHIP_RAM.N_340 ));
    Odrv4 I__863 (
            .O(N__5396),
            .I(\U712_CHIP_RAM.N_340 ));
    CascadeMux I__862 (
            .O(N__5391),
            .I(\U712_CHIP_RAM.N_340_cascade_ ));
    InMux I__861 (
            .O(N__5388),
            .I(N__5383));
    CascadeMux I__860 (
            .O(N__5387),
            .I(N__5379));
    InMux I__859 (
            .O(N__5386),
            .I(N__5372));
    LocalMux I__858 (
            .O(N__5383),
            .I(N__5369));
    InMux I__857 (
            .O(N__5382),
            .I(N__5366));
    InMux I__856 (
            .O(N__5379),
            .I(N__5363));
    InMux I__855 (
            .O(N__5378),
            .I(N__5358));
    InMux I__854 (
            .O(N__5377),
            .I(N__5358));
    InMux I__853 (
            .O(N__5376),
            .I(N__5355));
    InMux I__852 (
            .O(N__5375),
            .I(N__5352));
    LocalMux I__851 (
            .O(N__5372),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7 ));
    Odrv4 I__850 (
            .O(N__5369),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7 ));
    LocalMux I__849 (
            .O(N__5366),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7 ));
    LocalMux I__848 (
            .O(N__5363),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7 ));
    LocalMux I__847 (
            .O(N__5358),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7 ));
    LocalMux I__846 (
            .O(N__5355),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7 ));
    LocalMux I__845 (
            .O(N__5352),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7 ));
    InMux I__844 (
            .O(N__5337),
            .I(N__5334));
    LocalMux I__843 (
            .O(N__5334),
            .I(\U712_CHIP_RAM.N_267 ));
    CascadeMux I__842 (
            .O(N__5331),
            .I(\U712_CHIP_RAM.N_281_cascade_ ));
    InMux I__841 (
            .O(N__5328),
            .I(N__5325));
    LocalMux I__840 (
            .O(N__5325),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_0_i_0 ));
    InMux I__839 (
            .O(N__5322),
            .I(N__5316));
    InMux I__838 (
            .O(N__5321),
            .I(N__5316));
    LocalMux I__837 (
            .O(N__5316),
            .I(\U712_CHIP_RAM.N_207_i ));
    InMux I__836 (
            .O(N__5313),
            .I(N__5310));
    LocalMux I__835 (
            .O(N__5310),
            .I(N__5307));
    Span4Mux_v I__834 (
            .O(N__5307),
            .I(N__5304));
    Sp12to4 I__833 (
            .O(N__5304),
            .I(N__5301));
    Span12Mux_h I__832 (
            .O(N__5301),
            .I(N__5298));
    Odrv12 I__831 (
            .O(N__5298),
            .I(A_c_11));
    InMux I__830 (
            .O(N__5295),
            .I(N__5292));
    LocalMux I__829 (
            .O(N__5292),
            .I(N__5289));
    Span12Mux_v I__828 (
            .O(N__5289),
            .I(N__5286));
    Span12Mux_h I__827 (
            .O(N__5286),
            .I(N__5283));
    Odrv12 I__826 (
            .O(N__5283),
            .I(A_c_4));
    InMux I__825 (
            .O(N__5280),
            .I(N__5277));
    LocalMux I__824 (
            .O(N__5277),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    SRMux I__823 (
            .O(N__5274),
            .I(N__5271));
    LocalMux I__822 (
            .O(N__5271),
            .I(N__5268));
    Span4Mux_h I__821 (
            .O(N__5268),
            .I(N__5265));
    Odrv4 I__820 (
            .O(N__5265),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__819 (
            .O(N__5262),
            .I(N__5259));
    LocalMux I__818 (
            .O(N__5259),
            .I(N__5256));
    Span4Mux_v I__817 (
            .O(N__5256),
            .I(N__5253));
    Sp12to4 I__816 (
            .O(N__5253),
            .I(N__5250));
    Span12Mux_h I__815 (
            .O(N__5250),
            .I(N__5247));
    Span12Mux_v I__814 (
            .O(N__5247),
            .I(N__5244));
    Odrv12 I__813 (
            .O(N__5244),
            .I(A_c_5));
    InMux I__812 (
            .O(N__5241),
            .I(N__5238));
    LocalMux I__811 (
            .O(N__5238),
            .I(N__5235));
    Span12Mux_h I__810 (
            .O(N__5235),
            .I(N__5232));
    Odrv12 I__809 (
            .O(N__5232),
            .I(A_c_12));
    InMux I__808 (
            .O(N__5229),
            .I(N__5226));
    LocalMux I__807 (
            .O(N__5226),
            .I(N__5223));
    Span4Mux_v I__806 (
            .O(N__5223),
            .I(N__5220));
    Span4Mux_v I__805 (
            .O(N__5220),
            .I(N__5217));
    Sp12to4 I__804 (
            .O(N__5217),
            .I(N__5214));
    Span12Mux_h I__803 (
            .O(N__5214),
            .I(N__5211));
    Odrv12 I__802 (
            .O(N__5211),
            .I(A_c_7));
    CascadeMux I__801 (
            .O(N__5208),
            .I(\U712_CHIP_RAM.N_347_cascade_ ));
    CascadeMux I__800 (
            .O(N__5205),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_1_cascade_ ));
    CascadeMux I__799 (
            .O(N__5202),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_cascade_ ));
    InMux I__798 (
            .O(N__5199),
            .I(N__5196));
    LocalMux I__797 (
            .O(N__5196),
            .I(\U712_CHIP_RAM.N_284 ));
    InMux I__796 (
            .O(N__5193),
            .I(N__5186));
    InMux I__795 (
            .O(N__5192),
            .I(N__5186));
    InMux I__794 (
            .O(N__5191),
            .I(N__5183));
    LocalMux I__793 (
            .O(N__5186),
            .I(\U712_REG_SM.N_215 ));
    LocalMux I__792 (
            .O(N__5183),
            .I(\U712_REG_SM.N_215 ));
    InMux I__791 (
            .O(N__5178),
            .I(N__5174));
    InMux I__790 (
            .O(N__5177),
            .I(N__5171));
    LocalMux I__789 (
            .O(N__5174),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__788 (
            .O(N__5171),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    CascadeMux I__787 (
            .O(N__5166),
            .I(\U712_REG_SM.N_215_cascade_ ));
    CascadeMux I__786 (
            .O(N__5163),
            .I(\U712_REG_SM.N_228_cascade_ ));
    CascadeMux I__785 (
            .O(N__5160),
            .I(\U712_REG_SM.STATE_COUNT_srsts_i_i_0_1_cascade_ ));
    InMux I__784 (
            .O(N__5157),
            .I(N__5154));
    LocalMux I__783 (
            .O(N__5154),
            .I(N__5150));
    IoInMux I__782 (
            .O(N__5153),
            .I(N__5147));
    Span4Mux_v I__781 (
            .O(N__5150),
            .I(N__5144));
    LocalMux I__780 (
            .O(N__5147),
            .I(N__5141));
    Sp12to4 I__779 (
            .O(N__5144),
            .I(N__5138));
    Span4Mux_s3_h I__778 (
            .O(N__5141),
            .I(N__5135));
    Span12Mux_h I__777 (
            .O(N__5138),
            .I(N__5130));
    Sp12to4 I__776 (
            .O(N__5135),
            .I(N__5130));
    Span12Mux_v I__775 (
            .O(N__5130),
            .I(N__5127));
    Odrv12 I__774 (
            .O(N__5127),
            .I(C1_c));
    InMux I__773 (
            .O(N__5124),
            .I(N__5120));
    IoInMux I__772 (
            .O(N__5123),
            .I(N__5117));
    LocalMux I__771 (
            .O(N__5120),
            .I(N__5114));
    LocalMux I__770 (
            .O(N__5117),
            .I(N__5111));
    Span4Mux_v I__769 (
            .O(N__5114),
            .I(N__5108));
    IoSpan4Mux I__768 (
            .O(N__5111),
            .I(N__5105));
    Sp12to4 I__767 (
            .O(N__5108),
            .I(N__5102));
    IoSpan4Mux I__766 (
            .O(N__5105),
            .I(N__5099));
    Span12Mux_h I__765 (
            .O(N__5102),
            .I(N__5096));
    IoSpan4Mux I__764 (
            .O(N__5099),
            .I(N__5093));
    Odrv12 I__763 (
            .O(N__5096),
            .I(C3_c));
    Odrv4 I__762 (
            .O(N__5093),
            .I(C3_c));
    InMux I__761 (
            .O(N__5088),
            .I(N__5085));
    LocalMux I__760 (
            .O(N__5085),
            .I(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_1 ));
    InMux I__759 (
            .O(N__5082),
            .I(N__5079));
    LocalMux I__758 (
            .O(N__5079),
            .I(N__5076));
    Span12Mux_h I__757 (
            .O(N__5076),
            .I(N__5073));
    Odrv12 I__756 (
            .O(N__5073),
            .I(RAS1n_c));
    InMux I__755 (
            .O(N__5070),
            .I(N__5064));
    InMux I__754 (
            .O(N__5069),
            .I(N__5064));
    LocalMux I__753 (
            .O(N__5064),
            .I(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_0 ));
    InMux I__752 (
            .O(N__5061),
            .I(N__5058));
    LocalMux I__751 (
            .O(N__5058),
            .I(N__5055));
    Span4Mux_v I__750 (
            .O(N__5055),
            .I(N__5051));
    InMux I__749 (
            .O(N__5054),
            .I(N__5048));
    Sp12to4 I__748 (
            .O(N__5051),
            .I(N__5045));
    LocalMux I__747 (
            .O(N__5048),
            .I(N__5042));
    Span12Mux_h I__746 (
            .O(N__5045),
            .I(N__5039));
    Span12Mux_h I__745 (
            .O(N__5042),
            .I(N__5036));
    Span12Mux_v I__744 (
            .O(N__5039),
            .I(N__5033));
    Span12Mux_v I__743 (
            .O(N__5036),
            .I(N__5030));
    Odrv12 I__742 (
            .O(N__5033),
            .I(TSn_c));
    Odrv12 I__741 (
            .O(N__5030),
            .I(TSn_c));
    CascadeMux I__740 (
            .O(N__5025),
            .I(N__5022));
    InMux I__739 (
            .O(N__5022),
            .I(N__5019));
    LocalMux I__738 (
            .O(N__5019),
            .I(N__5016));
    Span4Mux_v I__737 (
            .O(N__5016),
            .I(N__5013));
    Span4Mux_v I__736 (
            .O(N__5013),
            .I(N__5010));
    Sp12to4 I__735 (
            .O(N__5010),
            .I(N__5007));
    Span12Mux_h I__734 (
            .O(N__5007),
            .I(N__5004));
    Odrv12 I__733 (
            .O(N__5004),
            .I(REGSPACEn_c));
    InMux I__732 (
            .O(N__5001),
            .I(N__4998));
    LocalMux I__731 (
            .O(N__4998),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_2 ));
    CascadeMux I__730 (
            .O(N__4995),
            .I(N__4991));
    CascadeMux I__729 (
            .O(N__4994),
            .I(N__4988));
    InMux I__728 (
            .O(N__4991),
            .I(N__4985));
    InMux I__727 (
            .O(N__4988),
            .I(N__4982));
    LocalMux I__726 (
            .O(N__4985),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__725 (
            .O(N__4982),
            .I(DBR_SYNCZ0Z_1));
    InMux I__724 (
            .O(N__4977),
            .I(N__4973));
    InMux I__723 (
            .O(N__4976),
            .I(N__4970));
    LocalMux I__722 (
            .O(N__4973),
            .I(DBR_SYNCZ0Z_0));
    LocalMux I__721 (
            .O(N__4970),
            .I(DBR_SYNCZ0Z_0));
    CascadeMux I__720 (
            .O(N__4965),
            .I(\U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_1_2_cascade_ ));
    CascadeMux I__719 (
            .O(N__4962),
            .I(N__4958));
    InMux I__718 (
            .O(N__4961),
            .I(N__4955));
    InMux I__717 (
            .O(N__4958),
            .I(N__4952));
    LocalMux I__716 (
            .O(N__4955),
            .I(\U712_REG_SM.N_245 ));
    LocalMux I__715 (
            .O(N__4952),
            .I(\U712_REG_SM.N_245 ));
    InMux I__714 (
            .O(N__4947),
            .I(N__4944));
    LocalMux I__713 (
            .O(N__4944),
            .I(\U712_CHIP_RAM.N_209 ));
    CascadeMux I__712 (
            .O(N__4941),
            .I(\U712_CHIP_RAM.N_209_cascade_ ));
    InMux I__711 (
            .O(N__4938),
            .I(N__4935));
    LocalMux I__710 (
            .O(N__4935),
            .I(\U712_CHIP_RAM.N_263 ));
    InMux I__709 (
            .O(N__4932),
            .I(N__4929));
    LocalMux I__708 (
            .O(N__4929),
            .I(\U712_CHIP_RAM.N_246 ));
    CascadeMux I__707 (
            .O(N__4926),
            .I(N__4923));
    InMux I__706 (
            .O(N__4923),
            .I(N__4920));
    LocalMux I__705 (
            .O(N__4920),
            .I(N__4911));
    InMux I__704 (
            .O(N__4919),
            .I(N__4908));
    InMux I__703 (
            .O(N__4918),
            .I(N__4904));
    InMux I__702 (
            .O(N__4917),
            .I(N__4901));
    InMux I__701 (
            .O(N__4916),
            .I(N__4898));
    InMux I__700 (
            .O(N__4915),
            .I(N__4893));
    InMux I__699 (
            .O(N__4914),
            .I(N__4893));
    Span4Mux_h I__698 (
            .O(N__4911),
            .I(N__4888));
    LocalMux I__697 (
            .O(N__4908),
            .I(N__4888));
    InMux I__696 (
            .O(N__4907),
            .I(N__4885));
    LocalMux I__695 (
            .O(N__4904),
            .I(N__4882));
    LocalMux I__694 (
            .O(N__4901),
            .I(\U712_CHIP_RAM.N_332 ));
    LocalMux I__693 (
            .O(N__4898),
            .I(\U712_CHIP_RAM.N_332 ));
    LocalMux I__692 (
            .O(N__4893),
            .I(\U712_CHIP_RAM.N_332 ));
    Odrv4 I__691 (
            .O(N__4888),
            .I(\U712_CHIP_RAM.N_332 ));
    LocalMux I__690 (
            .O(N__4885),
            .I(\U712_CHIP_RAM.N_332 ));
    Odrv4 I__689 (
            .O(N__4882),
            .I(\U712_CHIP_RAM.N_332 ));
    InMux I__688 (
            .O(N__4869),
            .I(N__4865));
    InMux I__687 (
            .O(N__4868),
            .I(N__4862));
    LocalMux I__686 (
            .O(N__4865),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__685 (
            .O(N__4862),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__684 (
            .O(N__4857),
            .I(N__4850));
    InMux I__683 (
            .O(N__4856),
            .I(N__4850));
    InMux I__682 (
            .O(N__4855),
            .I(N__4847));
    LocalMux I__681 (
            .O(N__4850),
            .I(N__4844));
    LocalMux I__680 (
            .O(N__4847),
            .I(\U712_CHIP_RAM.N_203 ));
    Odrv4 I__679 (
            .O(N__4844),
            .I(\U712_CHIP_RAM.N_203 ));
    CascadeMux I__678 (
            .O(N__4839),
            .I(\U712_CHIP_RAM.N_203_cascade_ ));
    CascadeMux I__677 (
            .O(N__4836),
            .I(N__4833));
    InMux I__676 (
            .O(N__4833),
            .I(N__4830));
    LocalMux I__675 (
            .O(N__4830),
            .I(N__4827));
    Odrv4 I__674 (
            .O(N__4827),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_3_0 ));
    InMux I__673 (
            .O(N__4824),
            .I(N__4818));
    InMux I__672 (
            .O(N__4823),
            .I(N__4818));
    LocalMux I__671 (
            .O(N__4818),
            .I(\U712_CHIP_RAM.N_341 ));
    CEMux I__670 (
            .O(N__4815),
            .I(N__4812));
    LocalMux I__669 (
            .O(N__4812),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0 ));
    CascadeMux I__668 (
            .O(N__4809),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7_cascade_ ));
    InMux I__667 (
            .O(N__4806),
            .I(N__4803));
    LocalMux I__666 (
            .O(N__4803),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_0_0_i_1 ));
    CascadeMux I__665 (
            .O(N__4800),
            .I(\U712_CHIP_RAM.N_211_cascade_ ));
    InMux I__664 (
            .O(N__4797),
            .I(N__4794));
    LocalMux I__663 (
            .O(N__4794),
            .I(\U712_CHIP_RAM.N_87 ));
    InMux I__662 (
            .O(N__4791),
            .I(N__4788));
    LocalMux I__661 (
            .O(N__4788),
            .I(\U712_CHIP_RAM.N_266 ));
    CascadeMux I__660 (
            .O(N__4785),
            .I(N__4778));
    InMux I__659 (
            .O(N__4784),
            .I(N__4775));
    InMux I__658 (
            .O(N__4783),
            .I(N__4772));
    InMux I__657 (
            .O(N__4782),
            .I(N__4767));
    InMux I__656 (
            .O(N__4781),
            .I(N__4767));
    InMux I__655 (
            .O(N__4778),
            .I(N__4763));
    LocalMux I__654 (
            .O(N__4775),
            .I(N__4756));
    LocalMux I__653 (
            .O(N__4772),
            .I(N__4756));
    LocalMux I__652 (
            .O(N__4767),
            .I(N__4756));
    InMux I__651 (
            .O(N__4766),
            .I(N__4753));
    LocalMux I__650 (
            .O(N__4763),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__649 (
            .O(N__4756),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__648 (
            .O(N__4753),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    CascadeMux I__647 (
            .O(N__4746),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a3_0_0_cascade_ ));
    InMux I__646 (
            .O(N__4743),
            .I(N__4739));
    InMux I__645 (
            .O(N__4742),
            .I(N__4736));
    LocalMux I__644 (
            .O(N__4739),
            .I(N__4733));
    LocalMux I__643 (
            .O(N__4736),
            .I(\U712_CHIP_RAM.N_264 ));
    Odrv4 I__642 (
            .O(N__4733),
            .I(\U712_CHIP_RAM.N_264 ));
    CascadeMux I__641 (
            .O(N__4728),
            .I(\U712_CHIP_RAM.N_264_cascade_ ));
    CascadeMux I__640 (
            .O(N__4725),
            .I(\U712_CHIP_RAM.N_36_cascade_ ));
    InMux I__639 (
            .O(N__4722),
            .I(N__4718));
    InMux I__638 (
            .O(N__4721),
            .I(N__4715));
    LocalMux I__637 (
            .O(N__4718),
            .I(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1 ));
    LocalMux I__636 (
            .O(N__4715),
            .I(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1 ));
    CascadeMux I__635 (
            .O(N__4710),
            .I(\U712_CHIP_RAM.N_342_cascade_ ));
    InMux I__634 (
            .O(N__4707),
            .I(N__4703));
    InMux I__633 (
            .O(N__4706),
            .I(N__4700));
    LocalMux I__632 (
            .O(N__4703),
            .I(\U712_CHIP_RAM.N_381 ));
    LocalMux I__631 (
            .O(N__4700),
            .I(\U712_CHIP_RAM.N_381 ));
    CascadeMux I__630 (
            .O(N__4695),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_ ));
    InMux I__629 (
            .O(N__4692),
            .I(N__4689));
    LocalMux I__628 (
            .O(N__4689),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_0 ));
    CascadeMux I__627 (
            .O(N__4686),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_1_cascade_ ));
    InMux I__626 (
            .O(N__4683),
            .I(N__4680));
    LocalMux I__625 (
            .O(N__4680),
            .I(N__4677));
    Sp12to4 I__624 (
            .O(N__4677),
            .I(N__4674));
    Span12Mux_v I__623 (
            .O(N__4674),
            .I(N__4671));
    Span12Mux_h I__622 (
            .O(N__4671),
            .I(N__4668));
    Odrv12 I__621 (
            .O(N__4668),
            .I(A_c_8));
    InMux I__620 (
            .O(N__4665),
            .I(N__4662));
    LocalMux I__619 (
            .O(N__4662),
            .I(N__4659));
    Span4Mux_v I__618 (
            .O(N__4659),
            .I(N__4656));
    Span4Mux_v I__617 (
            .O(N__4656),
            .I(N__4653));
    Sp12to4 I__616 (
            .O(N__4653),
            .I(N__4650));
    Odrv12 I__615 (
            .O(N__4650),
            .I(A_c_15));
    CascadeMux I__614 (
            .O(N__4647),
            .I(N__4644));
    InMux I__613 (
            .O(N__4644),
            .I(N__4640));
    InMux I__612 (
            .O(N__4643),
            .I(N__4637));
    LocalMux I__611 (
            .O(N__4640),
            .I(\U712_CHIP_RAM.N_270_4 ));
    LocalMux I__610 (
            .O(N__4637),
            .I(\U712_CHIP_RAM.N_270_4 ));
    CascadeMux I__609 (
            .O(N__4632),
            .I(\U712_REG_SM.STATE_COUNT_srsts_i_i_0_3_cascade_ ));
    InMux I__608 (
            .O(N__4629),
            .I(N__4626));
    LocalMux I__607 (
            .O(N__4626),
            .I(\U712_REG_SM.N_289 ));
    CascadeMux I__606 (
            .O(N__4623),
            .I(\U712_REG_SM.N_289_cascade_ ));
    InMux I__605 (
            .O(N__4620),
            .I(N__4608));
    InMux I__604 (
            .O(N__4619),
            .I(N__4608));
    InMux I__603 (
            .O(N__4618),
            .I(N__4608));
    InMux I__602 (
            .O(N__4617),
            .I(N__4608));
    LocalMux I__601 (
            .O(N__4608),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__600 (
            .O(N__4605),
            .I(N__4602));
    LocalMux I__599 (
            .O(N__4602),
            .I(N__4597));
    InMux I__598 (
            .O(N__4601),
            .I(N__4594));
    InMux I__597 (
            .O(N__4600),
            .I(N__4591));
    Span4Mux_h I__596 (
            .O(N__4597),
            .I(N__4583));
    LocalMux I__595 (
            .O(N__4594),
            .I(N__4583));
    LocalMux I__594 (
            .O(N__4591),
            .I(N__4583));
    InMux I__593 (
            .O(N__4590),
            .I(N__4580));
    Span4Mux_v I__592 (
            .O(N__4583),
            .I(N__4577));
    LocalMux I__591 (
            .O(N__4580),
            .I(N__4574));
    Sp12to4 I__590 (
            .O(N__4577),
            .I(N__4571));
    Span4Mux_v I__589 (
            .O(N__4574),
            .I(N__4568));
    Span12Mux_h I__588 (
            .O(N__4571),
            .I(N__4565));
    Span4Mux_h I__587 (
            .O(N__4568),
            .I(N__4562));
    Span12Mux_v I__586 (
            .O(N__4565),
            .I(N__4559));
    Span4Mux_h I__585 (
            .O(N__4562),
            .I(N__4556));
    Odrv12 I__584 (
            .O(N__4559),
            .I(RnW_c));
    Odrv4 I__583 (
            .O(N__4556),
            .I(RnW_c));
    CascadeMux I__582 (
            .O(N__4551),
            .I(\U712_CHIP_RAM.N_261_cascade_ ));
    IoInMux I__581 (
            .O(N__4548),
            .I(N__4545));
    LocalMux I__580 (
            .O(N__4545),
            .I(N__4542));
    IoSpan4Mux I__579 (
            .O(N__4542),
            .I(N__4539));
    Sp12to4 I__578 (
            .O(N__4539),
            .I(N__4536));
    Span12Mux_s7_h I__577 (
            .O(N__4536),
            .I(N__4533));
    Span12Mux_h I__576 (
            .O(N__4533),
            .I(N__4529));
    InMux I__575 (
            .O(N__4532),
            .I(N__4526));
    Odrv12 I__574 (
            .O(N__4529),
            .I(CLK_EN_c));
    LocalMux I__573 (
            .O(N__4526),
            .I(CLK_EN_c));
    InMux I__572 (
            .O(N__4521),
            .I(N__4518));
    LocalMux I__571 (
            .O(N__4518),
            .I(\U712_CHIP_RAM.N_260 ));
    CascadeMux I__570 (
            .O(N__4515),
            .I(N__4512));
    InMux I__569 (
            .O(N__4512),
            .I(N__4508));
    InMux I__568 (
            .O(N__4511),
            .I(N__4505));
    LocalMux I__567 (
            .O(N__4508),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__566 (
            .O(N__4505),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__565 (
            .O(N__4500),
            .I(N__4488));
    InMux I__564 (
            .O(N__4499),
            .I(N__4488));
    InMux I__563 (
            .O(N__4498),
            .I(N__4488));
    InMux I__562 (
            .O(N__4497),
            .I(N__4488));
    LocalMux I__561 (
            .O(N__4488),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__560 (
            .O(N__4485),
            .I(N__4482));
    LocalMux I__559 (
            .O(N__4482),
            .I(N__4478));
    InMux I__558 (
            .O(N__4481),
            .I(N__4475));
    Span4Mux_v I__557 (
            .O(N__4478),
            .I(N__4472));
    LocalMux I__556 (
            .O(N__4475),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv4 I__555 (
            .O(N__4472),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__554 (
            .O(N__4467),
            .I(N__4464));
    LocalMux I__553 (
            .O(N__4464),
            .I(N__4461));
    Odrv4 I__552 (
            .O(N__4461),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    CascadeMux I__551 (
            .O(N__4458),
            .I(N__4455));
    InMux I__550 (
            .O(N__4455),
            .I(N__4452));
    LocalMux I__549 (
            .O(N__4452),
            .I(N__4448));
    InMux I__548 (
            .O(N__4451),
            .I(N__4445));
    Span4Mux_v I__547 (
            .O(N__4448),
            .I(N__4442));
    LocalMux I__546 (
            .O(N__4445),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv4 I__545 (
            .O(N__4442),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__544 (
            .O(N__4437),
            .I(N__4434));
    LocalMux I__543 (
            .O(N__4434),
            .I(N__4431));
    Odrv12 I__542 (
            .O(N__4431),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    CascadeMux I__541 (
            .O(N__4428),
            .I(N__4425));
    InMux I__540 (
            .O(N__4425),
            .I(N__4422));
    LocalMux I__539 (
            .O(N__4422),
            .I(N__4419));
    Span4Mux_h I__538 (
            .O(N__4419),
            .I(N__4415));
    IoInMux I__537 (
            .O(N__4418),
            .I(N__4412));
    Sp12to4 I__536 (
            .O(N__4415),
            .I(N__4409));
    LocalMux I__535 (
            .O(N__4412),
            .I(N__4406));
    Span12Mux_v I__534 (
            .O(N__4409),
            .I(N__4403));
    IoSpan4Mux I__533 (
            .O(N__4406),
            .I(N__4400));
    Odrv12 I__532 (
            .O(N__4403),
            .I(RAMENn_c));
    Odrv4 I__531 (
            .O(N__4400),
            .I(RAMENn_c));
    CascadeMux I__530 (
            .O(N__4395),
            .I(N__4392));
    InMux I__529 (
            .O(N__4392),
            .I(N__4388));
    InMux I__528 (
            .O(N__4391),
            .I(N__4385));
    LocalMux I__527 (
            .O(N__4388),
            .I(REG_TACK));
    LocalMux I__526 (
            .O(N__4385),
            .I(REG_TACK));
    InMux I__525 (
            .O(N__4380),
            .I(N__4377));
    LocalMux I__524 (
            .O(N__4377),
            .I(\U712_REG_SM.N_225 ));
    CascadeMux I__523 (
            .O(N__4374),
            .I(\U712_REG_SM.N_225_cascade_ ));
    InMux I__522 (
            .O(N__4371),
            .I(N__4368));
    LocalMux I__521 (
            .O(N__4368),
            .I(\U712_REG_SM.N_292 ));
    InMux I__520 (
            .O(N__4365),
            .I(N__4362));
    LocalMux I__519 (
            .O(N__4362),
            .I(\U712_REG_SM.REG_TACK_RNOZ0Z_0 ));
    CascadeMux I__518 (
            .O(N__4359),
            .I(\U712_CHIP_RAM.N_332_cascade_ ));
    CascadeMux I__517 (
            .O(N__4356),
            .I(N__4353));
    InMux I__516 (
            .O(N__4353),
            .I(N__4350));
    LocalMux I__515 (
            .O(N__4350),
            .I(\U712_CHIP_RAM.A_m_2_20 ));
    InMux I__514 (
            .O(N__4347),
            .I(N__4344));
    LocalMux I__513 (
            .O(N__4344),
            .I(N__4341));
    Span4Mux_v I__512 (
            .O(N__4341),
            .I(N__4338));
    Sp12to4 I__511 (
            .O(N__4338),
            .I(N__4335));
    Span12Mux_h I__510 (
            .O(N__4335),
            .I(N__4332));
    Span12Mux_v I__509 (
            .O(N__4332),
            .I(N__4329));
    Odrv12 I__508 (
            .O(N__4329),
            .I(A_c_20));
    CascadeMux I__507 (
            .O(N__4326),
            .I(\U712_CHIP_RAM.A_m_2_20_cascade_ ));
    CascadeMux I__506 (
            .O(N__4323),
            .I(\U712_CHIP_RAM.BANK0_esr_RNOZ0Z_1_cascade_ ));
    IoInMux I__505 (
            .O(N__4320),
            .I(N__4317));
    LocalMux I__504 (
            .O(N__4317),
            .I(N__4314));
    Span4Mux_s3_v I__503 (
            .O(N__4314),
            .I(N__4311));
    Span4Mux_v I__502 (
            .O(N__4311),
            .I(N__4308));
    Span4Mux_v I__501 (
            .O(N__4308),
            .I(N__4305));
    Span4Mux_h I__500 (
            .O(N__4305),
            .I(N__4302));
    Odrv4 I__499 (
            .O(N__4302),
            .I(BANK0_c));
    CEMux I__498 (
            .O(N__4299),
            .I(N__4296));
    LocalMux I__497 (
            .O(N__4296),
            .I(N__4293));
    Odrv4 I__496 (
            .O(N__4293),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_10_0_0 ));
    InMux I__495 (
            .O(N__4290),
            .I(N__4287));
    LocalMux I__494 (
            .O(N__4287),
            .I(N__4284));
    Odrv4 I__493 (
            .O(N__4284),
            .I(\U712_CHIP_RAM.CPU_TACK_e_1 ));
    InMux I__492 (
            .O(N__4281),
            .I(N__4277));
    InMux I__491 (
            .O(N__4280),
            .I(N__4274));
    LocalMux I__490 (
            .O(N__4277),
            .I(CPU_TACKm));
    LocalMux I__489 (
            .O(N__4274),
            .I(CPU_TACKm));
    IoInMux I__488 (
            .O(N__4269),
            .I(N__4266));
    LocalMux I__487 (
            .O(N__4266),
            .I(N__4263));
    IoSpan4Mux I__486 (
            .O(N__4263),
            .I(N__4260));
    Span4Mux_s0_h I__485 (
            .O(N__4260),
            .I(N__4257));
    Sp12to4 I__484 (
            .O(N__4257),
            .I(N__4254));
    Span12Mux_s11_h I__483 (
            .O(N__4254),
            .I(N__4250));
    InMux I__482 (
            .O(N__4253),
            .I(N__4247));
    Odrv12 I__481 (
            .O(N__4250),
            .I(TACK_OUTn));
    LocalMux I__480 (
            .O(N__4247),
            .I(TACK_OUTn));
    InMux I__479 (
            .O(N__4242),
            .I(N__4237));
    InMux I__478 (
            .O(N__4241),
            .I(N__4234));
    InMux I__477 (
            .O(N__4240),
            .I(N__4231));
    LocalMux I__476 (
            .O(N__4237),
            .I(N__4228));
    LocalMux I__475 (
            .O(N__4234),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__474 (
            .O(N__4231),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    Odrv4 I__473 (
            .O(N__4228),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__472 (
            .O(N__4221),
            .I(N__4217));
    InMux I__471 (
            .O(N__4220),
            .I(N__4214));
    InMux I__470 (
            .O(N__4217),
            .I(N__4210));
    LocalMux I__469 (
            .O(N__4214),
            .I(N__4207));
    InMux I__468 (
            .O(N__4213),
            .I(N__4204));
    LocalMux I__467 (
            .O(N__4210),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv4 I__466 (
            .O(N__4207),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__465 (
            .O(N__4204),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__464 (
            .O(N__4197),
            .I(N__4194));
    LocalMux I__463 (
            .O(N__4194),
            .I(\U712_CHIP_RAM.N_243 ));
    InMux I__462 (
            .O(N__4191),
            .I(N__4188));
    LocalMux I__461 (
            .O(N__4188),
            .I(N__4185));
    Span12Mux_v I__460 (
            .O(N__4185),
            .I(N__4182));
    Odrv12 I__459 (
            .O(N__4182),
            .I(A_c_13));
    InMux I__458 (
            .O(N__4179),
            .I(N__4176));
    LocalMux I__457 (
            .O(N__4176),
            .I(N__4173));
    Span4Mux_h I__456 (
            .O(N__4173),
            .I(N__4170));
    Sp12to4 I__455 (
            .O(N__4170),
            .I(N__4167));
    Span12Mux_v I__454 (
            .O(N__4167),
            .I(N__4164));
    Odrv12 I__453 (
            .O(N__4164),
            .I(A_c_6));
    InMux I__452 (
            .O(N__4161),
            .I(N__4158));
    LocalMux I__451 (
            .O(N__4158),
            .I(N__4155));
    Span4Mux_h I__450 (
            .O(N__4155),
            .I(N__4152));
    Sp12to4 I__449 (
            .O(N__4152),
            .I(N__4149));
    Span12Mux_v I__448 (
            .O(N__4149),
            .I(N__4146));
    Odrv12 I__447 (
            .O(N__4146),
            .I(A_c_18));
    InMux I__446 (
            .O(N__4143),
            .I(N__4140));
    LocalMux I__445 (
            .O(N__4140),
            .I(N__4137));
    Span4Mux_v I__444 (
            .O(N__4137),
            .I(N__4134));
    Span4Mux_v I__443 (
            .O(N__4134),
            .I(N__4131));
    Sp12to4 I__442 (
            .O(N__4131),
            .I(N__4128));
    Span12Mux_h I__441 (
            .O(N__4128),
            .I(N__4125));
    Odrv12 I__440 (
            .O(N__4125),
            .I(A_c_16));
    IoInMux I__439 (
            .O(N__4122),
            .I(N__4119));
    LocalMux I__438 (
            .O(N__4119),
            .I(N__4116));
    Span12Mux_s4_v I__437 (
            .O(N__4116),
            .I(N__4113));
    Odrv12 I__436 (
            .O(N__4113),
            .I(N_187_i));
    CascadeMux I__435 (
            .O(N__4110),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_0_a3_0_cascade_ ));
    CascadeMux I__434 (
            .O(N__4107),
            .I(N__4104));
    InMux I__433 (
            .O(N__4104),
            .I(N__4101));
    LocalMux I__432 (
            .O(N__4101),
            .I(N__4097));
    InMux I__431 (
            .O(N__4100),
            .I(N__4094));
    Span4Mux_h I__430 (
            .O(N__4097),
            .I(N__4091));
    LocalMux I__429 (
            .O(N__4094),
            .I(\U712_CHIP_RAM.N_273 ));
    Odrv4 I__428 (
            .O(N__4091),
            .I(\U712_CHIP_RAM.N_273 ));
    CascadeMux I__427 (
            .O(N__4086),
            .I(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1_cascade_ ));
    CascadeMux I__426 (
            .O(N__4083),
            .I(\U712_CHIP_RAM.N_328_cascade_ ));
    CascadeMux I__425 (
            .O(N__4080),
            .I(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ));
    CascadeMux I__424 (
            .O(N__4077),
            .I(\U712_CYCLE_TERM.N_223_i_0_en_cascade_ ));
    InMux I__423 (
            .O(N__4074),
            .I(N__4071));
    LocalMux I__422 (
            .O(N__4071),
            .I(N__4068));
    Odrv4 I__421 (
            .O(N__4068),
            .I(TACK_EN_i_ess));
    CEMux I__420 (
            .O(N__4065),
            .I(N__4062));
    LocalMux I__419 (
            .O(N__4062),
            .I(N__4059));
    Span4Mux_v I__418 (
            .O(N__4059),
            .I(N__4056));
    Span4Mux_h I__417 (
            .O(N__4056),
            .I(N__4053));
    Odrv4 I__416 (
            .O(N__4053),
            .I(\U712_CYCLE_TERM.N_223_i_0_en_0 ));
    InMux I__415 (
            .O(N__4050),
            .I(N__4047));
    LocalMux I__414 (
            .O(N__4047),
            .I(N__4043));
    InMux I__413 (
            .O(N__4046),
            .I(N__4040));
    Span4Mux_v I__412 (
            .O(N__4043),
            .I(N__4034));
    LocalMux I__411 (
            .O(N__4040),
            .I(N__4034));
    InMux I__410 (
            .O(N__4039),
            .I(N__4031));
    Span4Mux_h I__409 (
            .O(N__4034),
            .I(N__4028));
    LocalMux I__408 (
            .O(N__4031),
            .I(N__4025));
    Sp12to4 I__407 (
            .O(N__4028),
            .I(N__4022));
    Span4Mux_v I__406 (
            .O(N__4025),
            .I(N__4019));
    Span12Mux_v I__405 (
            .O(N__4022),
            .I(N__4016));
    IoSpan4Mux I__404 (
            .O(N__4019),
            .I(N__4013));
    Odrv12 I__403 (
            .O(N__4016),
            .I(AWEn_c));
    Odrv4 I__402 (
            .O(N__4013),
            .I(AWEn_c));
    IoInMux I__401 (
            .O(N__4008),
            .I(N__4005));
    LocalMux I__400 (
            .O(N__4005),
            .I(N__4002));
    IoSpan4Mux I__399 (
            .O(N__4002),
            .I(N__3999));
    Span4Mux_s3_h I__398 (
            .O(N__3999),
            .I(N__3996));
    Sp12to4 I__397 (
            .O(N__3996),
            .I(N__3993));
    Span12Mux_s6_v I__396 (
            .O(N__3993),
            .I(N__3990));
    Span12Mux_h I__395 (
            .O(N__3990),
            .I(N__3987));
    Odrv12 I__394 (
            .O(N__3987),
            .I(N_242));
    InMux I__393 (
            .O(N__3984),
            .I(N__3980));
    InMux I__392 (
            .O(N__3983),
            .I(N__3977));
    LocalMux I__391 (
            .O(N__3980),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__390 (
            .O(N__3977),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    InMux I__389 (
            .O(N__3972),
            .I(N__3968));
    InMux I__388 (
            .O(N__3971),
            .I(N__3965));
    LocalMux I__387 (
            .O(N__3968),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    LocalMux I__386 (
            .O(N__3965),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    CascadeMux I__385 (
            .O(N__3960),
            .I(N__3956));
    InMux I__384 (
            .O(N__3959),
            .I(N__3953));
    InMux I__383 (
            .O(N__3956),
            .I(N__3950));
    LocalMux I__382 (
            .O(N__3953),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__381 (
            .O(N__3950),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__380 (
            .O(N__3945),
            .I(N__3941));
    InMux I__379 (
            .O(N__3944),
            .I(N__3938));
    LocalMux I__378 (
            .O(N__3941),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    LocalMux I__377 (
            .O(N__3938),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    CascadeMux I__376 (
            .O(N__3933),
            .I(\U712_CHIP_RAM.N_381_cascade_ ));
    IoInMux I__375 (
            .O(N__3930),
            .I(N__3927));
    LocalMux I__374 (
            .O(N__3927),
            .I(N__3924));
    Span12Mux_s9_v I__373 (
            .O(N__3924),
            .I(N__3921));
    Odrv12 I__372 (
            .O(N__3921),
            .I(VBENn_c));
    InMux I__371 (
            .O(N__3918),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    InMux I__370 (
            .O(N__3915),
            .I(N__3911));
    InMux I__369 (
            .O(N__3914),
            .I(N__3908));
    LocalMux I__368 (
            .O(N__3911),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__367 (
            .O(N__3908),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__366 (
            .O(N__3903),
            .I(N__3899));
    InMux I__365 (
            .O(N__3902),
            .I(N__3896));
    LocalMux I__364 (
            .O(N__3899),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__363 (
            .O(N__3896),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    IoInMux I__362 (
            .O(N__3891),
            .I(N__3888));
    LocalMux I__361 (
            .O(N__3888),
            .I(N__3884));
    CascadeMux I__360 (
            .O(N__3887),
            .I(N__3881));
    Span12Mux_s7_v I__359 (
            .O(N__3884),
            .I(N__3878));
    InMux I__358 (
            .O(N__3881),
            .I(N__3875));
    Odrv12 I__357 (
            .O(N__3878),
            .I(DBDIR_c));
    LocalMux I__356 (
            .O(N__3875),
            .I(DBDIR_c));
    CascadeMux I__355 (
            .O(N__3870),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0_cascade_ ));
    InMux I__354 (
            .O(N__3867),
            .I(N__3862));
    InMux I__353 (
            .O(N__3866),
            .I(N__3857));
    InMux I__352 (
            .O(N__3865),
            .I(N__3857));
    LocalMux I__351 (
            .O(N__3862),
            .I(N__3854));
    LocalMux I__350 (
            .O(N__3857),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_a3_0_0 ));
    Odrv4 I__349 (
            .O(N__3854),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_a3_0_0 ));
    IoInMux I__348 (
            .O(N__3849),
            .I(N__3846));
    LocalMux I__347 (
            .O(N__3846),
            .I(N__3843));
    Span4Mux_s2_v I__346 (
            .O(N__3843),
            .I(N__3840));
    Span4Mux_v I__345 (
            .O(N__3840),
            .I(N__3837));
    Span4Mux_h I__344 (
            .O(N__3837),
            .I(N__3834));
    Odrv4 I__343 (
            .O(N__3834),
            .I(CLK80_PLL_i_i));
    IoInMux I__342 (
            .O(N__3831),
            .I(N__3828));
    LocalMux I__341 (
            .O(N__3828),
            .I(N__3825));
    Span4Mux_s2_h I__340 (
            .O(N__3825),
            .I(N__3822));
    Sp12to4 I__339 (
            .O(N__3822),
            .I(N__3819));
    Span12Mux_v I__338 (
            .O(N__3819),
            .I(N__3816));
    Odrv12 I__337 (
            .O(N__3816),
            .I(N_1012_i));
    InMux I__336 (
            .O(N__3813),
            .I(bfn_7_5_0_));
    InMux I__335 (
            .O(N__3810),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__334 (
            .O(N__3807),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__333 (
            .O(N__3804),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__332 (
            .O(N__3801),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__331 (
            .O(N__3798),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__330 (
            .O(N__3795),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    IoInMux I__329 (
            .O(N__3792),
            .I(N__3789));
    LocalMux I__328 (
            .O(N__3789),
            .I(N__3786));
    IoSpan4Mux I__327 (
            .O(N__3786),
            .I(N__3783));
    Span4Mux_s2_v I__326 (
            .O(N__3783),
            .I(N__3780));
    Sp12to4 I__325 (
            .O(N__3780),
            .I(N__3777));
    Span12Mux_v I__324 (
            .O(N__3777),
            .I(N__3774));
    Odrv12 I__323 (
            .O(N__3774),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__7733));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__7734));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__7731));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__7732));
    defparam IN_MUX_bfv_10_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_8_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_5_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7560),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__5153),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__5123),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_5_1_3.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_5_1_3.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_5_1_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_5_1_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8736),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_obuft_RNO_LC_6_12_3.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_6_12_3.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_6_12_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 TACKn_obuft_RNO_LC_6_12_3 (
            .in0(N__4074),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_1012_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_5_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_5_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(N__3945),
            .in2(_gnd_net_),
            .in3(N__3813),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_7_5_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__7730),
            .ce(),
            .sr(N__5274));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_5_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_5_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_5_1  (
            .in0(_gnd_net_),
            .in1(N__3972),
            .in2(_gnd_net_),
            .in3(N__3810),
            .lcout(\U712_CHIP_RAM.REFRESH5lto1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__7730),
            .ce(),
            .sr(N__5274));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_5_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_5_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_5_2  (
            .in0(_gnd_net_),
            .in1(N__3984),
            .in2(_gnd_net_),
            .in3(N__3807),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__7730),
            .ce(),
            .sr(N__5274));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_5_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_5_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_5_3  (
            .in0(_gnd_net_),
            .in1(N__4481),
            .in2(_gnd_net_),
            .in3(N__3804),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__7730),
            .ce(),
            .sr(N__5274));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_5_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_5_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_5_4  (
            .in0(_gnd_net_),
            .in1(N__3959),
            .in2(_gnd_net_),
            .in3(N__3801),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__7730),
            .ce(),
            .sr(N__5274));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_5_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_5_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_5_5  (
            .in0(_gnd_net_),
            .in1(N__3903),
            .in2(_gnd_net_),
            .in3(N__3798),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__7730),
            .ce(),
            .sr(N__5274));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_5_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_5_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_5_6  (
            .in0(_gnd_net_),
            .in1(N__3915),
            .in2(_gnd_net_),
            .in3(N__3795),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__7730),
            .ce(),
            .sr(N__5274));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_5_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_5_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_5_7  (
            .in0(_gnd_net_),
            .in1(N__4451),
            .in2(_gnd_net_),
            .in3(N__3918),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7730),
            .ce(),
            .sr(N__5274));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_7_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_7_6_3 .LUT_INIT=16'b0011111100101111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_7_6_3  (
            .in0(N__9615),
            .in1(N__7349),
            .in2(N__8456),
            .in3(N__7275),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_7_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_7_6_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(N__3914),
            .in2(_gnd_net_),
            .in3(N__3902),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_7_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_7_7_4 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_7_7_4  (
            .in0(N__4100),
            .in1(N__9619),
            .in2(N__4356),
            .in3(N__6135),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8719),
            .ce(),
            .sr(N__10115));
    defparam \U712_CHIP_RAM.DBDIR_LC_7_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_7_7_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_7_7_7 .LUT_INIT=16'b0111010011110000;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_7_7_7  (
            .in0(N__4050),
            .in1(N__3867),
            .in2(N__3887),
            .in3(N__4917),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8719),
            .ce(),
            .sr(N__10115));
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_7_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_7_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_7_8_2 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_LC_7_8_2  (
            .in0(N__4915),
            .in1(N__9476),
            .in2(N__4107),
            .in3(N__3866),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8723),
            .ce(),
            .sr(N__10109));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_7_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_7_8_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_7_8_5  (
            .in0(N__3865),
            .in1(N__4743),
            .in2(_gnd_net_),
            .in3(N__4914),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_7_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_7_8_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_7_8_6 .LUT_INIT=16'b1100101011111010;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_7_8_6  (
            .in0(N__9358),
            .in1(N__5813),
            .in2(N__3870),
            .in3(N__8040),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8723),
            .ce(),
            .sr(N__10109));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_7_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_7_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__6250),
            .in2(_gnd_net_),
            .in3(N__6118),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_9_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_9_1  (
            .in0(N__6251),
            .in1(N__4046),
            .in2(_gnd_net_),
            .in3(N__4605),
            .lcout(\U712_CHIP_RAM.N_243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_7_9_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_7_9_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(N__4280),
            .in2(_gnd_net_),
            .in3(N__4391),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_7_9_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_7_9_3 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_7_9_3  (
            .in0(N__7698),
            .in1(N__4213),
            .in2(N__4080),
            .in3(N__4511),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_223_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_7_9_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_7_9_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_7_9_4  (
            .in0(N__10139),
            .in1(_gnd_net_),
            .in2(N__4077),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.N_223_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_10_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_10_4 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_10_4 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_10_4  (
            .in0(N__4220),
            .in1(N__7697),
            .in2(_gnd_net_),
            .in3(N__4241),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8730),
            .ce(N__4065),
            .sr(N__10096));
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_7_20_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_7_20_2 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_m2_LC_7_20_2  (
            .in0(N__4590),
            .in1(N__4039),
            .in2(_gnd_net_),
            .in3(N__9523),
            .lcout(N_242),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_5_0 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_5_0  (
            .in0(N__3983),
            .in1(N__3971),
            .in2(N__3960),
            .in3(N__3944),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_2_LC_8_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_2_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_2_LC_8_6_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_2_LC_8_6_0  (
            .in0(N__5814),
            .in1(N__5696),
            .in2(_gnd_net_),
            .in3(N__6168),
            .lcout(\U712_CHIP_RAM.N_381 ),
            .ltout(\U712_CHIP_RAM.N_381_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_6_1 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_6_1  (
            .in0(N__6169),
            .in1(N__4643),
            .in2(N__3933),
            .in3(N__5916),
            .lcout(\U712_CHIP_RAM.CPU_TACK_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a3_LC_8_6_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a3_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a3_LC_8_6_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a3_LC_8_6_2  (
            .in0(N__8523),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9620),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_8_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_8_6_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_8_6_3  (
            .in0(N__4191),
            .in1(_gnd_net_),
            .in2(N__8403),
            .in3(N__4179),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_8_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_8_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_8_6_4  (
            .in0(N__4161),
            .in1(N__4143),
            .in2(_gnd_net_),
            .in3(N__8364),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_187_i_LC_8_6_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_187_i_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_187_i_LC_8_6_5 .LUT_INIT=16'b0001001100110001;
    LogicCell40 \U712_BYTE_ENABLE.N_187_i_LC_8_6_5  (
            .in0(N__9621),
            .in1(N__8766),
            .in2(N__9860),
            .in3(N__10207),
            .lcout(N_187_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_0_LC_8_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_0_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_0_LC_8_6_6 .LUT_INIT=16'b0100000101000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_0_LC_8_6_6  (
            .in0(N__5815),
            .in1(N__5697),
            .in2(N__6015),
            .in3(N__4783),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_0_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_8_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_8_6_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_8_6_7  (
            .in0(N__6133),
            .in1(N__5915),
            .in2(N__4110),
            .in3(N__5382),
            .lcout(\U712_CHIP_RAM.N_273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNI4ICS5_LC_8_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNI4ICS5_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNI4ICS5_LC_8_7_0 .LUT_INIT=16'b1010000010100010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNI4ICS5_LC_8_7_0  (
            .in0(N__4907),
            .in1(N__6289),
            .in2(N__6258),
            .in3(N__4857),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_8_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_8_7_1 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_8_7_1  (
            .in0(N__4742),
            .in1(N__10140),
            .in2(N__4086),
            .in3(N__6136),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_10_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI85LA2_1_LC_8_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI85LA2_1_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI85LA2_1_LC_8_7_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI85LA2_1_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__6007),
            .in2(_gnd_net_),
            .in3(N__5375),
            .lcout(\U712_CHIP_RAM.N_328 ),
            .ltout(\U712_CHIP_RAM.N_328_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_8_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_8_7_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_8_7_3  (
            .in0(N__5774),
            .in1(N__5913),
            .in2(N__4083),
            .in3(N__5666),
            .lcout(\U712_CHIP_RAM.N_332 ),
            .ltout(\U712_CHIP_RAM.N_332_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNI4ICS5_0_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNI4ICS5_0_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNI4ICS5_0_LC_8_7_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNI4ICS5_0_LC_8_7_4  (
            .in0(N__6256),
            .in1(N__6288),
            .in2(N__4359),
            .in3(N__4856),
            .lcout(\U712_CHIP_RAM.A_m_2_20 ),
            .ltout(\U712_CHIP_RAM.A_m_2_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_7_5 .LUT_INIT=16'b0011111111111111;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__4347),
            .in2(N__4326),
            .in3(N__9129),
            .lcout(),
            .ltout(\U712_CHIP_RAM.BANK0_esr_RNOZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_LC_8_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_esr_LC_8_7_6 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_LC_8_7_6  (
            .in0(N__6257),
            .in1(N__4916),
            .in2(N__4323),
            .in3(N__7137),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8715),
            .ce(N__4299),
            .sr(N__10110));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_8_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_8_0 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_8_8_0  (
            .in0(N__6705),
            .in1(N__4240),
            .in2(N__4515),
            .in3(N__4497),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8720),
            .ce(),
            .sr(N__10100));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_8_1 .LUT_INIT=16'b1000100010111000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_8_8_1  (
            .in0(N__4281),
            .in1(N__4797),
            .in2(N__9660),
            .in3(N__4290),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8720),
            .ce(),
            .sr(N__10100));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_8_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_8_2 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_8_2 .LUT_INIT=16'b1111111110100010;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_8_8_2  (
            .in0(N__4253),
            .in1(N__4499),
            .in2(N__7914),
            .in3(N__6736),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8720),
            .ce(),
            .sr(N__10100));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_8_8_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_8_8_3 .LUT_INIT=16'b1011101010110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_8_8_3  (
            .in0(N__4500),
            .in1(N__4242),
            .in2(N__4221),
            .in3(N__7912),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8720),
            .ce(),
            .sr(N__10100));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_8_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_8_8_4 .LUT_INIT=16'b0111001011110000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_8_8_4  (
            .in0(N__6142),
            .in1(N__4197),
            .in2(N__4785),
            .in3(N__4721),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8720),
            .ce(),
            .sr(N__10100));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_8_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6719),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8720),
            .ce(),
            .sr(N__10100));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_8_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6737),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8720),
            .ce(),
            .sr(N__10100));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_8_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_8_8_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_8_8_7  (
            .in0(N__4498),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7908),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8720),
            .ce(),
            .sr(N__10100));
    defparam \U712_CHIP_RAM.REFRESH_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_8_9_0 .LUT_INIT=16'b1111001111111011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_8_9_0  (
            .in0(N__4485),
            .in1(N__4467),
            .in2(N__4458),
            .in3(N__4437),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8724),
            .ce(),
            .sr(N__10097));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_9_7 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_9_7  (
            .in0(N__5054),
            .in1(N__9639),
            .in2(N__4428),
            .in3(N__4869),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8724),
            .ce(),
            .sr(N__10097));
    defparam \U712_REG_SM.REG_TACK_LC_8_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_8_10_2 .LUT_INIT=16'b1011100010101010;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_8_10_2  (
            .in0(N__4365),
            .in1(N__4371),
            .in2(N__4395),
            .in3(N__4380),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8727),
            .ce(),
            .sr(N__10091));
    defparam \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_8_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_8_11_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_8_11_0  (
            .in0(N__4618),
            .in1(N__6550),
            .in2(_gnd_net_),
            .in3(N__6693),
            .lcout(\U712_REG_SM.N_225 ),
            .ltout(\U712_REG_SM.N_225_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_11_1 .LUT_INIT=16'b0001001100010001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_8_11_1  (
            .in0(N__7614),
            .in1(N__4629),
            .in2(N__4374),
            .in3(N__6498),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8731),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_8_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_8_11_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_8_11_2  (
            .in0(N__6692),
            .in1(N__6549),
            .in2(_gnd_net_),
            .in3(N__5191),
            .lcout(\U712_REG_SM.N_292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_8_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_8_11_3 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_8_11_3  (
            .in0(N__5597),
            .in1(N__4601),
            .in2(N__6662),
            .in3(N__4617),
            .lcout(\U712_REG_SM.REG_TACK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_8_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_8_11_4 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_8_11_4  (
            .in0(N__4619),
            .in1(N__7617),
            .in2(_gnd_net_),
            .in3(N__6694),
            .lcout(),
            .ltout(\U712_REG_SM.STATE_COUNT_srsts_i_i_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_8_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_8_11_5 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_8_11_5  (
            .in0(N__6695),
            .in1(N__5192),
            .in2(N__4632),
            .in3(N__4961),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8731),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIEMV42_4_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIEMV42_4_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIEMV42_4_LC_8_11_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIEMV42_4_LC_8_11_6  (
            .in0(N__6657),
            .in1(N__7616),
            .in2(_gnd_net_),
            .in3(N__5596),
            .lcout(\U712_REG_SM.N_289 ),
            .ltout(\U712_REG_SM.N_289_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_8_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_8_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_8_11_7 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_8_11_7  (
            .in0(N__7615),
            .in1(N__5193),
            .in2(N__4623),
            .in3(N__4620),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8731),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_8_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_8_12_7 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_8_12_7  (
            .in0(N__4600),
            .in1(N__6653),
            .in2(_gnd_net_),
            .in3(N__6588),
            .lcout(\U712_REG_SM.DS_EN_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_5_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_5_0  (
            .in0(N__5905),
            .in1(N__4784),
            .in2(N__6150),
            .in3(N__4707),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_261_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_5_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_5_1 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__4532),
            .in2(N__4551),
            .in3(N__4521),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8710),
            .ce(),
            .sr(N__10116));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_5_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_5_2  (
            .in0(N__6012),
            .in1(N__6188),
            .in2(N__6149),
            .in3(N__5388),
            .lcout(\U712_CHIP_RAM.N_260 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS6PC1_2_LC_9_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS6PC1_2_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS6PC1_2_LC_9_5_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIS6PC1_2_LC_9_5_6  (
            .in0(N__5904),
            .in1(N__5816),
            .in2(_gnd_net_),
            .in3(N__5701),
            .lcout(\U712_CHIP_RAM.N_342 ),
            .ltout(\U712_CHIP_RAM.N_342_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_5_7 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_5_7  (
            .in0(N__5817),
            .in1(N__5706),
            .in2(N__4710),
            .in3(N__6011),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_6_0 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_6_0  (
            .in0(N__5414),
            .in1(_gnd_net_),
            .in2(N__4647),
            .in3(N__6170),
            .lcout(\U712_CHIP_RAM.N_284 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2B8VE_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2B8VE_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2B8VE_LC_9_6_1 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2B8VE_LC_9_6_1  (
            .in0(N__5337),
            .in1(N__4706),
            .in2(N__4836),
            .in3(N__4791),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_9_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_9_6_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4695),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_6_3 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_6_3  (
            .in0(N__4692),
            .in1(N__5699),
            .in2(N__6013),
            .in3(N__6117),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_6_4 .LUT_INIT=16'b1011101110111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_6_4  (
            .in0(N__8821),
            .in1(N__5431),
            .in2(N__4686),
            .in3(N__5442),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8712),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_6_5  (
            .in0(N__4683),
            .in1(N__4665),
            .in2(_gnd_net_),
            .in3(N__8369),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_6_6 .LUT_INIT=16'b1010111100111111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_6_6  (
            .in0(N__4782),
            .in1(N__5700),
            .in2(N__6134),
            .in3(N__5903),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_0_0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILL8G1_LC_9_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILL8G1_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNILL8G1_LC_9_6_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNILL8G1_LC_9_6_7  (
            .in0(N__5811),
            .in1(N__5698),
            .in2(N__5914),
            .in3(N__4781),
            .lcout(\U712_CHIP_RAM.N_270_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_9_7_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_9_7_2  (
            .in0(N__7692),
            .in1(N__6300),
            .in2(N__5613),
            .in3(N__5454),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8713),
            .ce(N__4815),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_7_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_7_3  (
            .in0(N__5468),
            .in1(N__5483),
            .in2(N__5502),
            .in3(N__6338),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_9_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_9_7_4 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__5788),
            .in2(N__4809),
            .in3(N__5979),
            .lcout(\U712_CHIP_RAM.N_211 ),
            .ltout(\U712_CHIP_RAM.N_211_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_7_5 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__4806),
            .in2(N__4800),
            .in3(N__4932),
            .lcout(\U712_CHIP_RAM.N_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_9_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_9_7_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_9_7_7  (
            .in0(N__5787),
            .in1(N__7693),
            .in2(N__5387),
            .in3(N__4947),
            .lcout(\U712_CHIP_RAM.N_266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_9_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_9_8_0 .LUT_INIT=16'b1000001010000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_9_8_0  (
            .in0(N__5781),
            .in1(N__5670),
            .in2(N__6000),
            .in3(N__4766),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_9_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_9_8_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_9_8_1  (
            .in0(N__5869),
            .in1(N__6110),
            .in2(N__4746),
            .in3(N__5377),
            .lcout(\U712_CHIP_RAM.N_264 ),
            .ltout(\U712_CHIP_RAM.N_264_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_9_8_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_9_8_2  (
            .in0(N__7662),
            .in1(N__4938),
            .in2(N__4728),
            .in3(N__4919),
            .lcout(\U712_CHIP_RAM.N_36 ),
            .ltout(\U712_CHIP_RAM.N_36_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_3 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_3  (
            .in0(N__5410),
            .in1(N__5517),
            .in2(N__4725),
            .in3(N__4722),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8716),
            .ce(N__6327),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_1_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_1_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_1_LC_9_8_4 .LUT_INIT=16'b0000010000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_1_LC_9_8_4  (
            .in0(N__6109),
            .in1(N__5669),
            .in2(N__5999),
            .in3(N__5868),
            .lcout(\U712_CHIP_RAM.N_209 ),
            .ltout(\U712_CHIP_RAM.N_209_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_9_8_5 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__5782),
            .in2(N__4941),
            .in3(N__5378),
            .lcout(\U712_CHIP_RAM.N_263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_6 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_6  (
            .in0(N__6201),
            .in1(N__6369),
            .in2(N__4926),
            .in3(N__5529),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8716),
            .ce(N__6327),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_8_7 .LUT_INIT=16'b1111000010100011;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_8_7  (
            .in0(N__5671),
            .in1(N__5783),
            .in2(N__5899),
            .in3(N__5978),
            .lcout(\U712_CHIP_RAM.N_246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNILCLN6_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNILCLN6_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNILCLN6_LC_9_9_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNILCLN6_LC_9_9_0  (
            .in0(N__4855),
            .in1(N__4824),
            .in2(N__5415),
            .in3(N__4918),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861_1_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861_1_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861_1_LC_9_9_1 .LUT_INIT=16'b0011011100111111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861_1_LC_9_9_1  (
            .in0(N__5069),
            .in1(N__4868),
            .in2(N__4994),
            .in3(N__5088),
            .lcout(\U712_CHIP_RAM.N_203 ),
            .ltout(\U712_CHIP_RAM.N_203_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH0703_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH0703_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH0703_LC_9_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH0703_LC_9_9_2  (
            .in0(N__7661),
            .in1(N__4823),
            .in2(N__4839),
            .in3(N__6083),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_3  (
            .in0(N__9513),
            .in1(N__5001),
            .in2(N__6242),
            .in3(N__7119),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8721),
            .ce(),
            .sr(N__10092));
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIRILU_LC_9_9_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIRILU_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__6276),
            .in2(_gnd_net_),
            .in3(N__6226),
            .lcout(\U712_CHIP_RAM.N_341 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_SYNC_1_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_1_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_1_LC_9_9_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_SYNC_1_LC_9_9_5  (
            .in0(N__5070),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8721),
            .ce(),
            .sr(N__10092));
    defparam \U712_CHIP_RAM.REFRESH_SYNC_0_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_0_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_SYNC_0_LC_9_9_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.REFRESH_SYNC_0_LC_9_9_6  (
            .in0(N__5082),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9162),
            .lcout(\U712_CHIP_RAM.REFRESH_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8721),
            .ce(),
            .sr(N__10092));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_10_1 .LUT_INIT=16'b0000010111001101;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_9_10_1  (
            .in0(N__5061),
            .in1(N__5178),
            .in2(N__5025),
            .in3(N__8512),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8725),
            .ce(),
            .sr(N__10086));
    defparam DBR_SYNC_0_LC_9_10_3.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_9_10_3.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_9_10_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 DBR_SYNC_0_LC_9_10_3 (
            .in0(N__7811),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8725),
            .ce(),
            .sr(N__10086));
    defparam DBR_SYNC_1_LC_9_10_5.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_9_10_5.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_9_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_9_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4977),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8725),
            .ce(),
            .sr(N__10086));
    defparam \U712_CHIP_RAM.CAS_SYNC_2_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_2_LC_9_10_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_2_LC_9_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_2_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8538),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8725),
            .ce(),
            .sr(N__10086));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_9_11_0 .LUT_INIT=16'b1000000011000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_9_11_0  (
            .in0(N__6696),
            .in1(N__7612),
            .in2(N__4962),
            .in3(N__7085),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8728),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI07K21_1_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI07K21_1_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI07K21_1_LC_9_11_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI07K21_1_LC_9_11_1  (
            .in0(N__6586),
            .in1(N__6623),
            .in2(N__4995),
            .in3(N__4976),
            .lcout(),
            .ltout(\U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI35EO1_1_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI35EO1_1_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI35EO1_1_LC_9_11_2 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI35EO1_1_LC_9_11_2  (
            .in0(N__5582),
            .in1(_gnd_net_),
            .in2(N__4965),
            .in3(N__5560),
            .lcout(\U712_REG_SM.N_245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_9_11_3 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_9_11_3  (
            .in0(N__6585),
            .in1(N__5559),
            .in2(N__6627),
            .in3(N__5580),
            .lcout(\U712_REG_SM.N_215 ),
            .ltout(\U712_REG_SM.N_215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_9_11_4 .LUT_INIT=16'b1111001111110011;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__5177),
            .in2(N__5166),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.N_228 ),
            .ltout(\U712_REG_SM.N_228_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_11_5 .LUT_INIT=16'b1101010111110111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_11_5  (
            .in0(N__7613),
            .in1(N__6479),
            .in2(N__5163),
            .in3(N__6554),
            .lcout(),
            .ltout(\U712_REG_SM.STATE_COUNT_srsts_i_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_11_6 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_9_11_6  (
            .in0(N__6624),
            .in1(N__6587),
            .in2(N__5160),
            .in3(N__7749),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8728),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_9_11_7 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_9_11_7  (
            .in0(N__6584),
            .in1(N__5558),
            .in2(N__6626),
            .in3(N__5581),
            .lcout(\U712_REG_SM.N_210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_12_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5157),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8732),
            .ce(),
            .sr(N__10081));
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_12_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5562),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8732),
            .ce(),
            .sr(N__10081));
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_12_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6591),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8732),
            .ce(),
            .sr(N__10081));
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_12_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5124),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8732),
            .ce(),
            .sr(N__10081));
    defparam \U712_REG_SM.REG_CYCLE_LC_9_19_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_19_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_19_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_9_19_2  (
            .in0(N__6464),
            .in1(N__7696),
            .in2(_gnd_net_),
            .in3(N__7789),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8893),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_10_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_10_5_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_10_5_0  (
            .in0(N__8813),
            .in1(N__7530),
            .in2(N__8269),
            .in3(N__8396),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_5_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_5_2  (
            .in0(N__5262),
            .in1(N__5241),
            .in2(_gnd_net_),
            .in3(N__8397),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_5_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_5_5  (
            .in0(N__5229),
            .in1(N__9688),
            .in2(_gnd_net_),
            .in3(N__8577),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_347_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_6 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_6  (
            .in0(N__7336),
            .in1(_gnd_net_),
            .in2(N__5208),
            .in3(N__8398),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_10_6_0 .LUT_INIT=16'b0000000000111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_10_6_0  (
            .in0(N__8270),
            .in1(N__7532),
            .in2(N__8399),
            .in3(N__8814),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_0_LC_10_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_0_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_0_LC_10_6_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_0_LC_10_6_1  (
            .in0(N__7533),
            .in1(N__8360),
            .in2(_gnd_net_),
            .in3(N__8271),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_6_2 .LUT_INIT=16'b0111111101101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_6_2  (
            .in0(N__5705),
            .in1(N__6132),
            .in2(N__6014),
            .in3(N__5906),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_3  (
            .in0(N__5386),
            .in1(N__7694),
            .in2(N__5205),
            .in3(N__5812),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_6_4 .LUT_INIT=16'b1000100010001011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_6_4  (
            .in0(N__8272),
            .in1(N__5432),
            .in2(N__5202),
            .in3(N__5199),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8711),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_6_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_6_5  (
            .in0(N__9683),
            .in1(N__5280),
            .in2(N__8430),
            .in3(N__7941),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIISK15_2_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIISK15_2_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIISK15_2_LC_10_6_6 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIISK15_2_LC_10_6_6  (
            .in0(N__7695),
            .in1(N__5535),
            .in2(_gnd_net_),
            .in3(N__5453),
            .lcout(\U712_CHIP_RAM.N_64_1 ),
            .ltout(\U712_CHIP_RAM.N_64_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_6_7 .LUT_INIT=16'b1101110111011000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_6_7  (
            .in0(N__5433),
            .in1(N__7540),
            .in2(N__5418),
            .in3(N__5328),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8711),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(N__7685),
            .in2(_gnd_net_),
            .in3(N__6106),
            .lcout(\U712_CHIP_RAM.N_340 ),
            .ltout(\U712_CHIP_RAM.N_340_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_10_7_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_10_7_1  (
            .in0(N__5886),
            .in1(N__5321),
            .in2(N__5391),
            .in3(N__5376),
            .lcout(\U712_CHIP_RAM.N_267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_10_7_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_10_7_3  (
            .in0(N__5890),
            .in1(N__5790),
            .in2(_gnd_net_),
            .in3(N__5971),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_281_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_7_4 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_7_4  (
            .in0(N__5322),
            .in1(_gnd_net_),
            .in2(N__5331),
            .in3(N__6108),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_10_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_10_7_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_10_7_5  (
            .in0(_gnd_net_),
            .in1(N__5667),
            .in2(_gnd_net_),
            .in3(N__5970),
            .lcout(\U712_CHIP_RAM.N_207_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_6  (
            .in0(N__5313),
            .in1(N__5295),
            .in2(_gnd_net_),
            .in3(N__8368),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNINN5O1_2_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNINN5O1_2_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNINN5O1_2_LC_10_7_7 .LUT_INIT=16'b0001000100011100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNINN5O1_2_LC_10_7_7  (
            .in0(N__6107),
            .in1(N__5789),
            .in2(N__5907),
            .in3(N__5668),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_8_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__5794),
            .in2(_gnd_net_),
            .in3(N__5523),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(bfn_10_8_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_8_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_8_1  (
            .in0(N__6370),
            .in1(N__5981),
            .in2(_gnd_net_),
            .in3(N__5520),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__8714),
            .ce(N__6323),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_8_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(N__5695),
            .in2(_gnd_net_),
            .in3(N__5508),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_8_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_8_3  (
            .in0(N__6371),
            .in1(N__5894),
            .in2(_gnd_net_),
            .in3(N__5505),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__8714),
            .ce(N__6323),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_8_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_8_4  (
            .in0(N__6366),
            .in1(N__5501),
            .in2(_gnd_net_),
            .in3(N__5487),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__8714),
            .ce(N__6323),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_8_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_8_5  (
            .in0(N__6372),
            .in1(N__5484),
            .in2(_gnd_net_),
            .in3(N__5472),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__8714),
            .ce(N__6323),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_8_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_8_6  (
            .in0(N__6367),
            .in1(N__5469),
            .in2(_gnd_net_),
            .in3(N__5457),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__8714),
            .ce(N__6323),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_8_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_8_7  (
            .in0(N__6339),
            .in1(N__6368),
            .in2(_gnd_net_),
            .in3(N__6342),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8714),
            .ce(N__6323),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_10_9_1 .LUT_INIT=16'b0101000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_10_9_1  (
            .in0(N__5793),
            .in1(N__6290),
            .in2(N__6252),
            .in3(N__6091),
            .lcout(\U712_CHIP_RAM.N_285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_9_2 .LUT_INIT=16'b0000101010001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_9_2  (
            .in0(N__7663),
            .in1(N__6291),
            .in2(N__6122),
            .in3(N__6241),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_a3_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_9_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_9_3  (
            .in0(N__6195),
            .in1(N__6095),
            .in2(_gnd_net_),
            .in3(N__6177),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8717),
            .ce(),
            .sr(N__10087));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_2_1_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_2_1_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_2_1_LC_10_9_5 .LUT_INIT=16'b1100110000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_2_1_LC_10_9_5  (
            .in0(N__5791),
            .in1(N__6090),
            .in2(_gnd_net_),
            .in3(N__5980),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_2_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_1_1_LC_10_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_1_1_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_1_1_LC_10_9_6 .LUT_INIT=16'b1111101111110110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_1_1_LC_10_9_6  (
            .in0(N__5898),
            .in1(N__5792),
            .in2(N__5709),
            .in3(N__5694),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_2_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_10_11_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_10_11_0  (
            .in0(N__6658),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5598),
            .lcout(\U712_REG_SM.ASn_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_3_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_3_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_3_LC_10_11_2 .LUT_INIT=16'b0111011111101110;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_3_LC_10_11_2  (
            .in0(N__6690),
            .in1(N__6622),
            .in2(_gnd_net_),
            .in3(N__6589),
            .lcout(),
            .ltout(\U712_REG_SM.N_248_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_10_11_3 .LUT_INIT=16'b1111000111110101;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_2_LC_10_11_3  (
            .in0(N__6547),
            .in1(N__5583),
            .in2(N__5565),
            .in3(N__5561),
            .lcout(\U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_10_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_10_11_4 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_10_11_4  (
            .in0(N__6691),
            .in1(N__6548),
            .in2(N__6663),
            .in3(N__7747),
            .lcout(\U712_REG_SM.N_300 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_10_11_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_10_11_6  (
            .in0(N__6625),
            .in1(N__6590),
            .in2(N__6555),
            .in3(N__7746),
            .lcout(\U712_REG_SM.N_226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_LC_10_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_10_12_0 .LUT_INIT=16'b1010101010001011;
    LogicCell40 \U712_REG_SM.DS_EN_LC_10_12_0  (
            .in0(N__10307),
            .in1(N__6522),
            .in2(N__6516),
            .in3(N__6504),
            .lcout(DS_ENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8729),
            .ce(),
            .sr(N__10078));
    defparam \U712_REG_SM.REGENn_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_10_12_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_10_12_5 .LUT_INIT=16'b1110101011111010;
    LogicCell40 \U712_REG_SM.REGENn_LC_10_12_5  (
            .in0(N__7098),
            .in1(N__6497),
            .in2(N__6460),
            .in3(N__6486),
            .lcout(REGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8729),
            .ce(),
            .sr(N__10078));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_4_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_11_4_4  (
            .in0(N__7203),
            .in1(N__8121),
            .in2(N__7359),
            .in3(N__6432),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8701),
            .ce(N__7385),
            .sr(N__10111));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_11_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_11_5_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__10138),
            .in2(_gnd_net_),
            .in3(N__6411),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_5_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_5_6  (
            .in0(N__9705),
            .in1(N__6405),
            .in2(N__8457),
            .in3(N__7929),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_11_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_11_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_11_6_2  (
            .in0(N__7293),
            .in1(N__6399),
            .in2(_gnd_net_),
            .in3(N__6777),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8706),
            .ce(N__7386),
            .sr(N__10098));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_6_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_6_5  (
            .in0(N__7531),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8255),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_11_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_11_6_7  (
            .in0(N__6819),
            .in1(N__6744),
            .in2(_gnd_net_),
            .in3(N__6885),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8706),
            .ce(N__7386),
            .sr(N__10098));
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5_1_LC_11_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5_1_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5_1_LC_11_7_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5_1_LC_11_7_0  (
            .in0(N__8405),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9640),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_7_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_7_1  (
            .in0(N__6858),
            .in1(N__6840),
            .in2(_gnd_net_),
            .in3(N__8404),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_4 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_4  (
            .in0(N__7467),
            .in1(N__8132),
            .in2(N__9684),
            .in3(N__6767),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_7_5  (
            .in0(N__6813),
            .in1(N__6795),
            .in2(_gnd_net_),
            .in3(N__8406),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_6 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_6  (
            .in0(N__8407),
            .in1(N__9641),
            .in2(N__6780),
            .in3(N__7953),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_7 .LUT_INIT=16'b1110001011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_7  (
            .in0(N__8133),
            .in1(N__9642),
            .in2(N__6771),
            .in3(N__7468),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_8_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_8_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__6738),
            .in2(_gnd_net_),
            .in3(N__6720),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_LC_11_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_LC_11_11_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_LC_11_11_2 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U712_REG_SM.ASn_LC_11_11_2  (
            .in0(N__7055),
            .in1(N__7097),
            .in2(_gnd_net_),
            .in3(N__7086),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8722),
            .ce(),
            .sr(N__10079));
    defparam CONSTANT_ONE_LUT4_LC_12_1_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_3_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_3_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_12_3_0  (
            .in0(N__7550),
            .in1(N__8459),
            .in2(N__8835),
            .in3(N__8279),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8697),
            .ce(N__7407),
            .sr(N__10108));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_5_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_12_5_0  (
            .in0(N__7204),
            .in1(N__7284),
            .in2(N__7356),
            .in3(N__6900),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8700),
            .ce(N__7387),
            .sr(N__10095));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_5_1 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_12_5_1  (
            .in0(N__6996),
            .in1(N__7481),
            .in2(N__9722),
            .in3(N__9174),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8700),
            .ce(N__7387),
            .sr(N__10095));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_5_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_12_5_2  (
            .in0(N__7205),
            .in1(N__9234),
            .in2(N__7357),
            .in3(N__6960),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8700),
            .ce(N__7387),
            .sr(N__10095));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_5_4 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_12_5_4  (
            .in0(N__8103),
            .in1(N__7348),
            .in2(N__7209),
            .in3(N__7254),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8700),
            .ce(N__7387),
            .sr(N__10095));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_3  (
            .in0(N__9696),
            .in1(N__6906),
            .in2(N__8460),
            .in3(N__7992),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_6_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_6_5  (
            .in0(N__9697),
            .in1(N__6894),
            .in2(N__8461),
            .in3(N__8619),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_6_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_6_7  (
            .in0(N__9698),
            .in1(N__7248),
            .in2(N__8462),
            .in3(N__7146),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_7_1 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_7_1  (
            .in0(N__9646),
            .in1(N__7239),
            .in2(N__8458),
            .in3(N__8625),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_12_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_12_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_12_7_2 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_12_7_2  (
            .in0(N__7191),
            .in1(N__7346),
            .in2(N__7227),
            .in3(N__8109),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8705),
            .ce(N__7403),
            .sr(N__10085));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_7_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_12_7_6  (
            .in0(N__7192),
            .in1(N__7347),
            .in2(N__8094),
            .in3(N__7173),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8705),
            .ce(N__7403),
            .sr(N__10085));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_12_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_12_8_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_12_8_0  (
            .in0(N__8961),
            .in1(N__9125),
            .in2(_gnd_net_),
            .in3(N__9222),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__8561),
            .sr(N__10083));
    defparam \U712_CHIP_RAM.DMA_A20_LC_12_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_12_9_6 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_12_9_6  (
            .in0(N__9099),
            .in1(N__7104),
            .in2(N__8960),
            .in3(N__7133),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__10080));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_12_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_12_10_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__8534),
            .in2(_gnd_net_),
            .in3(N__8750),
            .lcout(\U712_CHIP_RAM.un5_DMA_CYCLE_START_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS10_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS10_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS10_LC_12_10_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS10_LC_12_10_2  (
            .in0(N__7804),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8901),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10 ),
            .ltout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_12_10_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7917),
            .in3(N__10137),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESS10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pll_RNI8MQ3_LC_12_11_5.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_12_11_5.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_12_11_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 pll_RNI8MQ3_LC_12_11_5 (
            .in0(N__7913),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_11_6 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_11_6  (
            .in0(N__10136),
            .in1(N__7812),
            .in2(_gnd_net_),
            .in3(N__7748),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESS9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_20_1.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_20_1.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_20_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7657),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RASn_LC_13_2_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_13_2_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_13_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_13_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7551),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8698),
            .ce(),
            .sr(N__10117));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_5_4 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_13_5_4  (
            .in0(N__7482),
            .in1(N__7449),
            .in2(N__9723),
            .in3(N__8913),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8703),
            .ce(N__7396),
            .sr(N__10101));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_6_7 .LUT_INIT=16'b0000010011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_6_7  (
            .in0(N__9695),
            .in1(N__7265),
            .in2(N__7358),
            .in3(N__8443),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_7_0  (
            .in0(N__9100),
            .in1(N__8027),
            .in2(_gnd_net_),
            .in3(N__8082),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8895),
            .ce(N__8866),
            .sr(N__10093));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_7_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_7_1  (
            .in0(N__8028),
            .in1(N__9101),
            .in2(_gnd_net_),
            .in3(N__7982),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8895),
            .ce(N__8866),
            .sr(N__10093));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_7_2 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_7_2  (
            .in0(N__7983),
            .in1(N__9276),
            .in2(N__9122),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8895),
            .ce(N__8866),
            .sr(N__10093));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_7_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_7_4  (
            .in0(N__8208),
            .in1(_gnd_net_),
            .in2(N__9123),
            .in3(N__9330),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8895),
            .ce(N__8866),
            .sr(N__10093));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_6  (
            .in0(N__8172),
            .in1(_gnd_net_),
            .in2(N__9124),
            .in3(N__8609),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8895),
            .ce(N__8866),
            .sr(N__10093));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_7_7  (
            .in0(N__8610),
            .in1(N__9221),
            .in2(_gnd_net_),
            .in3(N__9111),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8895),
            .ce(N__8866),
            .sr(N__10093));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_8_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_13_8_0  (
            .in0(N__8081),
            .in1(N__9084),
            .in2(_gnd_net_),
            .in3(N__8020),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__8565),
            .sr(N__10088));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_8_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_8_1  (
            .in0(N__8021),
            .in1(_gnd_net_),
            .in2(N__9118),
            .in3(N__7980),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__8565),
            .sr(N__10088));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_2  (
            .in0(N__7981),
            .in1(N__9088),
            .in2(_gnd_net_),
            .in3(N__9271),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__8565),
            .sr(N__10088));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_8_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_8_3  (
            .in0(N__9272),
            .in1(_gnd_net_),
            .in2(N__9119),
            .in3(N__9328),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__8565),
            .sr(N__10088));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_4  (
            .in0(N__9329),
            .in1(N__9092),
            .in2(_gnd_net_),
            .in3(N__8205),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__8565),
            .sr(N__10088));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_5  (
            .in0(N__8168),
            .in1(_gnd_net_),
            .in2(N__9120),
            .in3(N__8206),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__8565),
            .sr(N__10088));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7  (
            .in0(N__9220),
            .in1(_gnd_net_),
            .in2(N__9121),
            .in3(N__8608),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__8565),
            .sr(N__10088));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_0  (
            .in0(N__8167),
            .in1(N__9040),
            .in2(_gnd_net_),
            .in3(N__8607),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__8557),
            .sr(N__10084));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_10_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_13_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8751),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8718),
            .ce(),
            .sr(N__10082));
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_LC_13_20_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a3_LC_13_20_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a3_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__9522),
            .in2(_gnd_net_),
            .in3(N__8519),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_14_2_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_14_2_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_14_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_14_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8466),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8699),
            .ce(),
            .sr(N__10119));
    defparam \U712_CHIP_RAM.WEn_LC_14_3_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_14_3_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_14_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_14_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8280),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8702),
            .ce(),
            .sr(N__10118));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_6  (
            .in0(N__8207),
            .in1(N__9076),
            .in2(_gnd_net_),
            .in3(N__8166),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8897),
            .ce(N__8870),
            .sr(N__10099));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_6  (
            .in0(N__9324),
            .in1(N__9041),
            .in2(_gnd_net_),
            .in3(N__9257),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8896),
            .ce(N__8871),
            .sr(N__10094));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_7  (
            .in0(N__9210),
            .in1(_gnd_net_),
            .in2(N__9083),
            .in3(N__8947),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8896),
            .ce(N__8871),
            .sr(N__10094));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_9_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_9_7  (
            .in0(N__9158),
            .in1(N__9014),
            .in2(_gnd_net_),
            .in3(N__8946),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8894),
            .ce(N__8856),
            .sr(N__10089));
    defparam \U712_CHIP_RAM.CRCSn_LC_15_3_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_15_3_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_15_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_15_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8834),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8704),
            .ce(),
            .sr(N__10120));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_15_8_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_15_8_2 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_15_8_2  (
            .in0(N__10292),
            .in1(_gnd_net_),
            .in2(N__9770),
            .in3(N__9725),
            .lcout(\U712_BYTE_ENABLE.N_313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_15_8_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_15_8_3 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_15_8_3  (
            .in0(N__9724),
            .in1(N__9762),
            .in2(N__9875),
            .in3(N__10291),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_315_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_LC_15_8_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_LC_15_8_4 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_LC_15_8_4  (
            .in0(N__9374),
            .in1(N__9987),
            .in2(N__8769),
            .in3(N__9514),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_15_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_15_10_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_15_10_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_15_10_4  (
            .in0(N__9449),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9982),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8726),
            .ce(),
            .sr(N__10090));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_LC_16_7_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_LC_16_7_2 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_LC_16_7_2  (
            .in0(N__9392),
            .in1(N__9945),
            .in2(N__9986),
            .in3(N__9528),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_16_8_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_16_8_0 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_16_8_0  (
            .in0(N__10286),
            .in1(N__9766),
            .in2(N__9876),
            .in3(N__9718),
            .lcout(\U712_BYTE_ENABLE.N_311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_LC_16_8_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_LC_16_8_2 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_0_LC_16_8_2  (
            .in0(N__9939),
            .in1(N__9450),
            .in2(N__9524),
            .in3(N__9375),
            .lcout(\U712_BYTE_ENABLE.un1_CLMBEn_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_20_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_20_1 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_20_1  (
            .in0(N__10200),
            .in1(N__10274),
            .in2(_gnd_net_),
            .in3(N__10319),
            .lcout(N_170),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_174_i_LC_17_6_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_174_i_LC_17_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_174_i_LC_17_6_1 .LUT_INIT=16'b0001010101000101;
    LogicCell40 \U712_BYTE_ENABLE.N_174_i_LC_17_6_1  (
            .in0(N__9915),
            .in1(N__9879),
            .in2(N__9726),
            .in3(N__10231),
            .lcout(N_174_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_172_i_LC_17_7_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_172_i_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_172_i_LC_17_7_2 .LUT_INIT=16'b0001001000110011;
    LogicCell40 \U712_BYTE_ENABLE.N_172_i_LC_17_7_2  (
            .in0(N__9877),
            .in1(N__9336),
            .in2(N__10232),
            .in3(N__9647),
            .lcout(N_172_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_176_i_LC_17_7_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_176_i_LC_17_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_176_i_LC_17_7_6 .LUT_INIT=16'b0001001000110011;
    LogicCell40 \U712_BYTE_ENABLE.N_176_i_LC_17_7_6  (
            .in0(N__9878),
            .in1(N__9801),
            .in2(N__10233),
            .in3(N__9648),
            .lcout(N_176_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_17_8_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_17_8_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_17_8_0  (
            .in0(N__9774),
            .in1(N__10296),
            .in2(_gnd_net_),
            .in3(N__9709),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_LC_17_8_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_LC_17_8_1 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_LC_17_8_1  (
            .in0(N__9518),
            .in1(N__9442),
            .in2(N__9399),
            .in3(N__9385),
            .lcout(\U712_BYTE_ENABLE.un1_CUUBEn_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_17_20_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_17_20_2 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_17_20_2  (
            .in0(N__10320),
            .in1(N__10287),
            .in2(_gnd_net_),
            .in3(N__10216),
            .lcout(N_168),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 23 2024 21:58:14

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RAMENn : out std_logic;
    RASn : out std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__10315\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_OUT_i_i\ : std_logic;
signal \CLK40_OUT_i_i\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.un6_REG_CYCLE_START_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_GOZ0\ : std_logic;
signal \C1_c\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_r_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH6lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_0\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_168_0_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_2\ : std_logic;
signal \U712_REG_SM.N_175_cascade_\ : std_logic;
signal \U712_REG_SM.N_171_0\ : std_logic;
signal \U712_REG_SM.N_194_cascade_\ : std_logic;
signal \U712_REG_SM.N_169_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_1\ : std_logic;
signal \U712_REG_SM.N_170_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_174_cascade_\ : std_logic;
signal \U712_REG_SM.N_162_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_172_0\ : std_logic;
signal \U712_REG_SM.N_162_0\ : std_logic;
signal \U712_REG_SM.N_195\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_163_0\ : std_logic;
signal \U712_REG_SM.N_194\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_186_0\ : std_logic;
signal \N_510_i\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_43_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_a2_0_4_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\ : std_logic;
signal \U712_REG_SM.DS_EN_7_0\ : std_logic;
signal \U712_REG_SM.N_187\ : std_logic;
signal \U712_REG_SM.N_157_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_159_0\ : std_logic;
signal \U712_REG_SM.N_159_0_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.N_165_0\ : std_logic;
signal \U712_REG_SM.N_165_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_170_0\ : std_logic;
signal \U712_REG_SM.N_173_0\ : std_logic;
signal \U712_REG_SM.LDS_OUT_2_0_0\ : std_logic;
signal \U712_REG_SM.UDS_OUT_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_105_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_105\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER17_1\ : std_logic;
signal \U712_CHIP_RAM.N_50_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_43\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_tz_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_68\ : std_logic;
signal \U712_CHIP_RAM.N_98\ : std_logic;
signal \U712_CHIP_RAM.N_55_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_57_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_92_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_44\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_3\ : std_logic;
signal \U712_CHIP_RAM.N_106_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.N_100\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_6\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.un6_CPU_CYCLE_START_cascade_\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.N_49\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \CLK40_OUT_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \DRDDIR_0_i\ : std_logic;
signal \CLMBEn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1\ : std_logic;
signal \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1_cascade_\ : std_logic;
signal \CLLBEn_c\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_167_0\ : std_logic;
signal \U712_BYTE_ENABLE.LLBE_0\ : std_logic;
signal \U712_BYTE_ENABLE.LMBE_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.N_78_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_76_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_58\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c2\ : std_logic;
signal \U712_CHIP_RAM.N_46\ : std_logic;
signal \U712_CHIP_RAM.N_77\ : std_logic;
signal \U712_CHIP_RAM.N_99\ : std_logic;
signal \U712_CHIP_RAM.N_99_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_79\ : std_logic;
signal \U712_CHIP_RAM.N_93_1\ : std_logic;
signal \U712_CHIP_RAM.N_52\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_54\ : std_logic;
signal \U712_CHIP_RAM.N_50\ : std_logic;
signal \U712_CHIP_RAM.N_54_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_START_2_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_0_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_70_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_106\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER53_3_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_40\ : std_logic;
signal \U712_CHIP_RAM.N_40_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_51\ : std_logic;
signal \U712_CHIP_RAM.N_59\ : std_logic;
signal \U712_CHIP_RAM.N_59_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_45_0_0_en\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_0\ : std_logic;
signal \U712_BYTE_ENABLE.UMBE_0\ : std_logic;
signal \CUMBEn_c\ : std_logic;
signal \U712_BYTE_ENABLE.UUBE_0\ : std_logic;
signal \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_0\ : std_logic;
signal \CUUBEn_c\ : std_logic;
signal \U712_REG_SM.LDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_LDSn_i\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.N_33\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.N_35_cascade_\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.N_34\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.DBENn_7_0_a2_0\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_CYCLE_TERM.N_45_0_0_en_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS4\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.UDS_OUTZ0\ : std_logic;
signal \U712_REG_SM.DS_ENZ0\ : std_logic;
signal \U712_REG_SM_un1_UDSn_i\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_5_cascade_\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.N_32\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.N_36\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.N_31\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_6\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.N_37\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_7_cascade_\ : std_logic;
signal \A_c_18\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_38\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_OUT_i\,
            REFERENCECLK => \N__3711\,
            RESETB => \N__7125\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_OUT\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10315\,
            DIN => \N__10314\,
            DOUT => \N__10313\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10315\,
            PADOUT => \N__10314\,
            PADIN => \N__10313\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5436\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10306\,
            DIN => \N__10305\,
            DOUT => \N__10304\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10306\,
            PADOUT => \N__10305\,
            PADIN => \N__10304\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10297\,
            DIN => \N__10296\,
            DOUT => \N__10295\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10297\,
            PADOUT => \N__10296\,
            PADIN => \N__10295\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8568\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10288\,
            DIN => \N__10287\,
            DOUT => \N__10286\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10288\,
            PADOUT => \N__10287\,
            PADIN => \N__10286\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4983\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10279\,
            DIN => \N__10278\,
            DOUT => \N__10277\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10279\,
            PADOUT => \N__10278\,
            PADIN => \N__10277\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10270\,
            DIN => \N__10269\,
            DOUT => \N__10268\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10270\,
            PADOUT => \N__10269\,
            PADIN => \N__10268\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10261\,
            DIN => \N__10260\,
            DOUT => \N__10259\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10261\,
            PADOUT => \N__10260\,
            PADIN => \N__10259\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10252\,
            DIN => \N__10251\,
            DOUT => \N__10250\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10252\,
            PADOUT => \N__10251\,
            PADIN => \N__10250\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10243\,
            DIN => \N__10242\,
            DOUT => \N__10241\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10243\,
            PADOUT => \N__10242\,
            PADIN => \N__10241\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10234\,
            DIN => \N__10233\,
            DOUT => \N__10232\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10234\,
            PADOUT => \N__10233\,
            PADIN => \N__10232\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10225\,
            DIN => \N__10224\,
            DOUT => \N__10223\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10225\,
            PADOUT => \N__10224\,
            PADIN => \N__10223\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9129\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10216\,
            DIN => \N__10215\,
            DOUT => \N__10214\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10216\,
            PADOUT => \N__10215\,
            PADIN => \N__10214\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6989\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10207\,
            DIN => \N__10206\,
            DOUT => \N__10205\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10207\,
            PADOUT => \N__10206\,
            PADIN => \N__10205\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10198\,
            DIN => \N__10197\,
            DOUT => \N__10196\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10198\,
            PADOUT => \N__10197\,
            PADIN => \N__10196\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10189\,
            DIN => \N__10188\,
            DOUT => \N__10187\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10189\,
            PADOUT => \N__10188\,
            PADIN => \N__10187\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4077\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10180\,
            DIN => \N__10179\,
            DOUT => \N__10178\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10180\,
            PADOUT => \N__10179\,
            PADIN => \N__10178\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10171\,
            DIN => \N__10170\,
            DOUT => \N__10169\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10171\,
            PADOUT => \N__10170\,
            PADIN => \N__10169\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10162\,
            DIN => \N__10161\,
            DOUT => \N__10160\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10162\,
            PADOUT => \N__10161\,
            PADIN => \N__10160\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7803\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10153\,
            DIN => \N__10152\,
            DOUT => \N__10151\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10153\,
            PADOUT => \N__10152\,
            PADIN => \N__10151\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10144\,
            DIN => \N__10143\,
            DOUT => \N__10142\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10144\,
            PADOUT => \N__10143\,
            PADIN => \N__10142\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8517\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10135\,
            DIN => \N__10134\,
            DOUT => \N__10133\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10135\,
            PADOUT => \N__10134\,
            PADIN => \N__10133\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10126\,
            DIN => \N__10125\,
            DOUT => \N__10124\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10126\,
            PADOUT => \N__10125\,
            PADIN => \N__10124\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10117\,
            DIN => \N__10116\,
            DOUT => \N__10115\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10117\,
            PADOUT => \N__10116\,
            PADIN => \N__10115\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10108\,
            DIN => \N__10107\,
            DOUT => \N__10106\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10108\,
            PADOUT => \N__10107\,
            PADIN => \N__10106\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10099\,
            DIN => \N__10098\,
            DOUT => \N__10097\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10099\,
            PADOUT => \N__10098\,
            PADIN => \N__10097\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10090\,
            DIN => \N__10089\,
            DOUT => \N__10088\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10090\,
            PADOUT => \N__10089\,
            PADIN => \N__10088\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10081\,
            DIN => \N__10080\,
            DOUT => \N__10079\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10081\,
            PADOUT => \N__10080\,
            PADIN => \N__10079\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10072\,
            DIN => \N__10071\,
            DOUT => \N__10070\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10072\,
            PADOUT => \N__10071\,
            PADIN => \N__10070\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10063\,
            DIN => \N__10062\,
            DOUT => \N__10061\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10063\,
            PADOUT => \N__10062\,
            PADIN => \N__10061\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10054\,
            DIN => \N__10053\,
            DOUT => \N__10052\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10054\,
            PADOUT => \N__10053\,
            PADIN => \N__10052\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7650\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10045\,
            DIN => \N__10044\,
            DOUT => \N__10043\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10045\,
            PADOUT => \N__10044\,
            PADIN => \N__10043\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10036\,
            DIN => \N__10035\,
            DOUT => \N__10034\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10036\,
            PADOUT => \N__10035\,
            PADIN => \N__10034\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10027\,
            DIN => \N__10026\,
            DOUT => \N__10025\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10027\,
            PADOUT => \N__10026\,
            PADIN => \N__10025\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10018\,
            DIN => \N__10017\,
            DOUT => \N__10016\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10018\,
            PADOUT => \N__10017\,
            PADIN => \N__10016\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10009\,
            DIN => \N__10008\,
            DOUT => \N__10007\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10009\,
            PADOUT => \N__10008\,
            PADIN => \N__10007\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3789\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10000\,
            DIN => \N__9999\,
            DOUT => \N__9998\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10000\,
            PADOUT => \N__9999\,
            PADIN => \N__9998\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6372\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9991\,
            DIN => \N__9990\,
            DOUT => \N__9989\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9991\,
            PADOUT => \N__9990\,
            PADIN => \N__9989\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9982\,
            DIN => \N__9981\,
            DOUT => \N__9980\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9982\,
            PADOUT => \N__9981\,
            PADIN => \N__9980\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8793\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9973\,
            DIN => \N__9972\,
            DOUT => \N__9971\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9973\,
            PADOUT => \N__9972\,
            PADIN => \N__9971\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9964\,
            DIN => \N__9963\,
            DOUT => \N__9962\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9964\,
            PADOUT => \N__9963\,
            PADIN => \N__9962\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9955\,
            DIN => \N__9954\,
            DOUT => \N__9953\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9955\,
            PADOUT => \N__9954\,
            PADIN => \N__9953\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3804\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9946\,
            DIN => \N__9945\,
            DOUT => \N__9944\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9946\,
            PADOUT => \N__9945\,
            PADIN => \N__9944\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9937\,
            DIN => \N__9936\,
            DOUT => \N__9935\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9937\,
            PADOUT => \N__9936\,
            PADIN => \N__9935\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4137\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9928\,
            DIN => \N__9927\,
            DOUT => \N__9926\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9928\,
            PADOUT => \N__9927\,
            PADIN => \N__9926\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6348\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9919\,
            DIN => \N__9918\,
            DOUT => \N__9917\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9919\,
            PADOUT => \N__9918\,
            PADIN => \N__9917\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9910\,
            DIN => \N__9909\,
            DOUT => \N__9908\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9910\,
            PADOUT => \N__9909\,
            PADIN => \N__9908\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9901\,
            DIN => \N__9900\,
            DOUT => \N__9899\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9901\,
            PADOUT => \N__9900\,
            PADIN => \N__9899\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9892\,
            DIN => \N__9891\,
            DOUT => \N__9890\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9892\,
            PADOUT => \N__9891\,
            PADIN => \N__9890\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9108\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9883\,
            DIN => \N__9882\,
            DOUT => \N__9881\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9883\,
            PADOUT => \N__9882\,
            PADIN => \N__9881\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9874\,
            DIN => \N__9873\,
            DOUT => \N__9872\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9874\,
            PADOUT => \N__9873\,
            PADIN => \N__9872\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6702\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9865\,
            DIN => \N__9864\,
            DOUT => \N__9863\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9865\,
            PADOUT => \N__9864\,
            PADIN => \N__9863\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7149\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9856\,
            DIN => \N__9855\,
            DOUT => \N__9854\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9856\,
            PADOUT => \N__9855\,
            PADIN => \N__9854\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5457\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9847\,
            DIN => \N__9846\,
            DOUT => \N__9845\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9847\,
            PADOUT => \N__9846\,
            PADIN => \N__9845\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7590\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9838\,
            DIN => \N__9837\,
            DOUT => \N__9836\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9838\,
            PADOUT => \N__9837\,
            PADIN => \N__9836\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4133\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9829\,
            DIN => \N__9828\,
            DOUT => \N__9827\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9829\,
            PADOUT => \N__9828\,
            PADIN => \N__9827\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9820\,
            DIN => \N__9819\,
            DOUT => \N__9818\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9820\,
            PADOUT => \N__9819\,
            PADIN => \N__9818\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9811\,
            DIN => \N__9810\,
            DOUT => \N__9809\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9811\,
            PADOUT => \N__9810\,
            PADIN => \N__9809\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4959\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9802\,
            DIN => \N__9801\,
            DOUT => \N__9800\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9802\,
            PADOUT => \N__9801\,
            PADIN => \N__9800\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8922\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9793\,
            DIN => \N__9792\,
            DOUT => \N__9791\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9793\,
            PADOUT => \N__9792\,
            PADIN => \N__9791\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5022\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9784\,
            DIN => \N__9783\,
            DOUT => \N__9782\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9784\,
            PADOUT => \N__9783\,
            PADIN => \N__9782\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6456\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9775\,
            DIN => \N__9774\,
            DOUT => \N__9773\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9775\,
            PADOUT => \N__9774\,
            PADIN => \N__9773\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9766\,
            DIN => \N__9765\,
            DOUT => \N__9764\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9766\,
            PADOUT => \N__9765\,
            PADIN => \N__9764\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9757\,
            DIN => \N__9756\,
            DOUT => \N__9755\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9757\,
            PADOUT => \N__9756\,
            PADIN => \N__9755\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9748\,
            DIN => \N__9747\,
            DOUT => \N__9746\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9748\,
            PADOUT => \N__9747\,
            PADIN => \N__9746\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9739\,
            DIN => \N__9738\,
            DOUT => \N__9737\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9739\,
            PADOUT => \N__9738\,
            PADIN => \N__9737\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7437\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9730\,
            DIN => \N__9729\,
            DOUT => \N__9728\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9730\,
            PADOUT => \N__9729\,
            PADIN => \N__9728\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9721\,
            DIN => \N__9720\,
            DOUT => \N__9719\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9721\,
            PADOUT => \N__9720\,
            PADIN => \N__9719\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6411\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9712\,
            DIN => \N__9711\,
            DOUT => \N__9710\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9712\,
            PADOUT => \N__9711\,
            PADIN => \N__9710\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4089\,
            DIN0 => OPEN,
            DOUT0 => \N__4608\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9703\,
            DIN => \N__9702\,
            DOUT => \N__9701\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9703\,
            PADOUT => \N__9702\,
            PADIN => \N__9701\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6759\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9694\,
            DIN => \N__9693\,
            DOUT => \N__9692\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9694\,
            PADOUT => \N__9693\,
            PADIN => \N__9692\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9685\,
            DIN => \N__9684\,
            DOUT => \N__9683\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9685\,
            PADOUT => \N__9684\,
            PADIN => \N__9683\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9676\,
            DIN => \N__9675\,
            DOUT => \N__9674\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9676\,
            PADOUT => \N__9675\,
            PADIN => \N__9674\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7671\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9667\,
            DIN => \N__9666\,
            DOUT => \N__9665\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9667\,
            PADOUT => \N__9666\,
            PADIN => \N__9665\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9658\,
            DIN => \N__9657\,
            DOUT => \N__9656\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9658\,
            PADOUT => \N__9657\,
            PADIN => \N__9656\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9649\,
            DIN => \N__9648\,
            DOUT => \N__9647\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9649\,
            PADOUT => \N__9648\,
            PADIN => \N__9647\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9640\,
            DIN => \N__9639\,
            DOUT => \N__9638\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9640\,
            PADOUT => \N__9639\,
            PADIN => \N__9638\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9631\,
            DIN => \N__9630\,
            DOUT => \N__9629\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9631\,
            PADOUT => \N__9630\,
            PADIN => \N__9629\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7779\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9622\,
            DIN => \N__9621\,
            DOUT => \N__9620\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9622\,
            PADOUT => \N__9621\,
            PADIN => \N__9620\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7254\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9613\,
            DIN => \N__9612\,
            DOUT => \N__9611\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9613\,
            PADOUT => \N__9612\,
            PADIN => \N__9611\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4926\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9604\,
            DIN => \N__9603\,
            DOUT => \N__9602\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9604\,
            PADOUT => \N__9603\,
            PADIN => \N__9602\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2276\ : InMux
    port map (
            O => \N__9585\,
            I => \N__9582\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__9582\,
            I => \N__9578\
        );

    \I__2274\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9575\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__9578\,
            I => \N__9572\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__9575\,
            I => \N__9569\
        );

    \I__2271\ : Span4Mux_h
    port map (
            O => \N__9572\,
            I => \N__9564\
        );

    \I__2270\ : Span4Mux_v
    port map (
            O => \N__9569\,
            I => \N__9564\
        );

    \I__2269\ : Sp12to4
    port map (
            O => \N__9564\,
            I => \N__9561\
        );

    \I__2268\ : Span12Mux_h
    port map (
            O => \N__9561\,
            I => \N__9558\
        );

    \I__2267\ : Odrv12
    port map (
            O => \N__9558\,
            I => \RAS0n_c\
        );

    \I__2266\ : InMux
    port map (
            O => \N__9555\,
            I => \N__9551\
        );

    \I__2265\ : InMux
    port map (
            O => \N__9554\,
            I => \N__9548\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__9551\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__9548\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2262\ : InMux
    port map (
            O => \N__9543\,
            I => \N__9540\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__9540\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__2260\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9534\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__9534\,
            I => \N__9507\
        );

    \I__2258\ : ClkMux
    port map (
            O => \N__9533\,
            I => \N__9372\
        );

    \I__2257\ : ClkMux
    port map (
            O => \N__9532\,
            I => \N__9372\
        );

    \I__2256\ : ClkMux
    port map (
            O => \N__9531\,
            I => \N__9372\
        );

    \I__2255\ : ClkMux
    port map (
            O => \N__9530\,
            I => \N__9372\
        );

    \I__2254\ : ClkMux
    port map (
            O => \N__9529\,
            I => \N__9372\
        );

    \I__2253\ : ClkMux
    port map (
            O => \N__9528\,
            I => \N__9372\
        );

    \I__2252\ : ClkMux
    port map (
            O => \N__9527\,
            I => \N__9372\
        );

    \I__2251\ : ClkMux
    port map (
            O => \N__9526\,
            I => \N__9372\
        );

    \I__2250\ : ClkMux
    port map (
            O => \N__9525\,
            I => \N__9372\
        );

    \I__2249\ : ClkMux
    port map (
            O => \N__9524\,
            I => \N__9372\
        );

    \I__2248\ : ClkMux
    port map (
            O => \N__9523\,
            I => \N__9372\
        );

    \I__2247\ : ClkMux
    port map (
            O => \N__9522\,
            I => \N__9372\
        );

    \I__2246\ : ClkMux
    port map (
            O => \N__9521\,
            I => \N__9372\
        );

    \I__2245\ : ClkMux
    port map (
            O => \N__9520\,
            I => \N__9372\
        );

    \I__2244\ : ClkMux
    port map (
            O => \N__9519\,
            I => \N__9372\
        );

    \I__2243\ : ClkMux
    port map (
            O => \N__9518\,
            I => \N__9372\
        );

    \I__2242\ : ClkMux
    port map (
            O => \N__9517\,
            I => \N__9372\
        );

    \I__2241\ : ClkMux
    port map (
            O => \N__9516\,
            I => \N__9372\
        );

    \I__2240\ : ClkMux
    port map (
            O => \N__9515\,
            I => \N__9372\
        );

    \I__2239\ : ClkMux
    port map (
            O => \N__9514\,
            I => \N__9372\
        );

    \I__2238\ : ClkMux
    port map (
            O => \N__9513\,
            I => \N__9372\
        );

    \I__2237\ : ClkMux
    port map (
            O => \N__9512\,
            I => \N__9372\
        );

    \I__2236\ : ClkMux
    port map (
            O => \N__9511\,
            I => \N__9372\
        );

    \I__2235\ : ClkMux
    port map (
            O => \N__9510\,
            I => \N__9372\
        );

    \I__2234\ : Glb2LocalMux
    port map (
            O => \N__9507\,
            I => \N__9372\
        );

    \I__2233\ : ClkMux
    port map (
            O => \N__9506\,
            I => \N__9372\
        );

    \I__2232\ : ClkMux
    port map (
            O => \N__9505\,
            I => \N__9372\
        );

    \I__2231\ : ClkMux
    port map (
            O => \N__9504\,
            I => \N__9372\
        );

    \I__2230\ : ClkMux
    port map (
            O => \N__9503\,
            I => \N__9372\
        );

    \I__2229\ : ClkMux
    port map (
            O => \N__9502\,
            I => \N__9372\
        );

    \I__2228\ : ClkMux
    port map (
            O => \N__9501\,
            I => \N__9372\
        );

    \I__2227\ : ClkMux
    port map (
            O => \N__9500\,
            I => \N__9372\
        );

    \I__2226\ : ClkMux
    port map (
            O => \N__9499\,
            I => \N__9372\
        );

    \I__2225\ : ClkMux
    port map (
            O => \N__9498\,
            I => \N__9372\
        );

    \I__2224\ : ClkMux
    port map (
            O => \N__9497\,
            I => \N__9372\
        );

    \I__2223\ : ClkMux
    port map (
            O => \N__9496\,
            I => \N__9372\
        );

    \I__2222\ : ClkMux
    port map (
            O => \N__9495\,
            I => \N__9372\
        );

    \I__2221\ : ClkMux
    port map (
            O => \N__9494\,
            I => \N__9372\
        );

    \I__2220\ : ClkMux
    port map (
            O => \N__9493\,
            I => \N__9372\
        );

    \I__2219\ : ClkMux
    port map (
            O => \N__9492\,
            I => \N__9372\
        );

    \I__2218\ : ClkMux
    port map (
            O => \N__9491\,
            I => \N__9372\
        );

    \I__2217\ : ClkMux
    port map (
            O => \N__9490\,
            I => \N__9372\
        );

    \I__2216\ : ClkMux
    port map (
            O => \N__9489\,
            I => \N__9372\
        );

    \I__2215\ : ClkMux
    port map (
            O => \N__9488\,
            I => \N__9372\
        );

    \I__2214\ : ClkMux
    port map (
            O => \N__9487\,
            I => \N__9372\
        );

    \I__2213\ : ClkMux
    port map (
            O => \N__9486\,
            I => \N__9372\
        );

    \I__2212\ : ClkMux
    port map (
            O => \N__9485\,
            I => \N__9372\
        );

    \I__2211\ : ClkMux
    port map (
            O => \N__9484\,
            I => \N__9372\
        );

    \I__2210\ : ClkMux
    port map (
            O => \N__9483\,
            I => \N__9372\
        );

    \I__2209\ : ClkMux
    port map (
            O => \N__9482\,
            I => \N__9372\
        );

    \I__2208\ : ClkMux
    port map (
            O => \N__9481\,
            I => \N__9372\
        );

    \I__2207\ : ClkMux
    port map (
            O => \N__9480\,
            I => \N__9372\
        );

    \I__2206\ : ClkMux
    port map (
            O => \N__9479\,
            I => \N__9372\
        );

    \I__2205\ : GlobalMux
    port map (
            O => \N__9372\,
            I => \CLK80_OUT\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__9369\,
            I => \N__9366\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9366\,
            I => \N__9346\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9365\,
            I => \N__9346\
        );

    \I__2201\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9346\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9346\
        );

    \I__2199\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9343\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9361\,
            I => \N__9340\
        );

    \I__2197\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9337\
        );

    \I__2196\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9334\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9331\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9357\,
            I => \N__9326\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9356\,
            I => \N__9326\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9355\,
            I => \N__9323\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__9346\,
            I => \N__9315\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__9343\,
            I => \N__9307\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__9340\,
            I => \N__9304\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__9337\,
            I => \N__9298\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__9334\,
            I => \N__9289\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9331\,
            I => \N__9286\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__9326\,
            I => \N__9280\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__9323\,
            I => \N__9273\
        );

    \I__2183\ : SRMux
    port map (
            O => \N__9322\,
            I => \N__9177\
        );

    \I__2182\ : SRMux
    port map (
            O => \N__9321\,
            I => \N__9177\
        );

    \I__2181\ : SRMux
    port map (
            O => \N__9320\,
            I => \N__9177\
        );

    \I__2180\ : SRMux
    port map (
            O => \N__9319\,
            I => \N__9177\
        );

    \I__2179\ : SRMux
    port map (
            O => \N__9318\,
            I => \N__9177\
        );

    \I__2178\ : Glb2LocalMux
    port map (
            O => \N__9315\,
            I => \N__9177\
        );

    \I__2177\ : SRMux
    port map (
            O => \N__9314\,
            I => \N__9177\
        );

    \I__2176\ : SRMux
    port map (
            O => \N__9313\,
            I => \N__9177\
        );

    \I__2175\ : SRMux
    port map (
            O => \N__9312\,
            I => \N__9177\
        );

    \I__2174\ : SRMux
    port map (
            O => \N__9311\,
            I => \N__9177\
        );

    \I__2173\ : SRMux
    port map (
            O => \N__9310\,
            I => \N__9177\
        );

    \I__2172\ : Glb2LocalMux
    port map (
            O => \N__9307\,
            I => \N__9177\
        );

    \I__2171\ : Glb2LocalMux
    port map (
            O => \N__9304\,
            I => \N__9177\
        );

    \I__2170\ : SRMux
    port map (
            O => \N__9303\,
            I => \N__9177\
        );

    \I__2169\ : SRMux
    port map (
            O => \N__9302\,
            I => \N__9177\
        );

    \I__2168\ : SRMux
    port map (
            O => \N__9301\,
            I => \N__9177\
        );

    \I__2167\ : Glb2LocalMux
    port map (
            O => \N__9298\,
            I => \N__9177\
        );

    \I__2166\ : SRMux
    port map (
            O => \N__9297\,
            I => \N__9177\
        );

    \I__2165\ : SRMux
    port map (
            O => \N__9296\,
            I => \N__9177\
        );

    \I__2164\ : SRMux
    port map (
            O => \N__9295\,
            I => \N__9177\
        );

    \I__2163\ : SRMux
    port map (
            O => \N__9294\,
            I => \N__9177\
        );

    \I__2162\ : SRMux
    port map (
            O => \N__9293\,
            I => \N__9177\
        );

    \I__2161\ : SRMux
    port map (
            O => \N__9292\,
            I => \N__9177\
        );

    \I__2160\ : Glb2LocalMux
    port map (
            O => \N__9289\,
            I => \N__9177\
        );

    \I__2159\ : Glb2LocalMux
    port map (
            O => \N__9286\,
            I => \N__9177\
        );

    \I__2158\ : SRMux
    port map (
            O => \N__9285\,
            I => \N__9177\
        );

    \I__2157\ : SRMux
    port map (
            O => \N__9284\,
            I => \N__9177\
        );

    \I__2156\ : SRMux
    port map (
            O => \N__9283\,
            I => \N__9177\
        );

    \I__2155\ : Glb2LocalMux
    port map (
            O => \N__9280\,
            I => \N__9177\
        );

    \I__2154\ : SRMux
    port map (
            O => \N__9279\,
            I => \N__9177\
        );

    \I__2153\ : SRMux
    port map (
            O => \N__9278\,
            I => \N__9177\
        );

    \I__2152\ : SRMux
    port map (
            O => \N__9277\,
            I => \N__9177\
        );

    \I__2151\ : SRMux
    port map (
            O => \N__9276\,
            I => \N__9177\
        );

    \I__2150\ : Glb2LocalMux
    port map (
            O => \N__9273\,
            I => \N__9177\
        );

    \I__2149\ : SRMux
    port map (
            O => \N__9272\,
            I => \N__9177\
        );

    \I__2148\ : SRMux
    port map (
            O => \N__9271\,
            I => \N__9177\
        );

    \I__2147\ : SRMux
    port map (
            O => \N__9270\,
            I => \N__9177\
        );

    \I__2146\ : SRMux
    port map (
            O => \N__9269\,
            I => \N__9177\
        );

    \I__2145\ : SRMux
    port map (
            O => \N__9268\,
            I => \N__9177\
        );

    \I__2144\ : SRMux
    port map (
            O => \N__9267\,
            I => \N__9177\
        );

    \I__2143\ : SRMux
    port map (
            O => \N__9266\,
            I => \N__9177\
        );

    \I__2142\ : SRMux
    port map (
            O => \N__9265\,
            I => \N__9177\
        );

    \I__2141\ : SRMux
    port map (
            O => \N__9264\,
            I => \N__9177\
        );

    \I__2140\ : GlobalMux
    port map (
            O => \N__9177\,
            I => \N__9174\
        );

    \I__2139\ : gio2CtrlBuf
    port map (
            O => \N__9174\,
            I => \RESETn_c_i_g\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9168\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9168\,
            I => \N__9164\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9167\,
            I => \N__9161\
        );

    \I__2135\ : Span4Mux_h
    port map (
            O => \N__9164\,
            I => \N__9156\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9161\,
            I => \N__9156\
        );

    \I__2133\ : Span4Mux_h
    port map (
            O => \N__9156\,
            I => \N__9153\
        );

    \I__2132\ : Sp12to4
    port map (
            O => \N__9153\,
            I => \N__9150\
        );

    \I__2131\ : Span12Mux_v
    port map (
            O => \N__9150\,
            I => \N__9147\
        );

    \I__2130\ : Odrv12
    port map (
            O => \N__9147\,
            I => \DRA_c_1\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9141\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__9141\,
            I => \N__9138\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__9138\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9132\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__9132\,
            I => \U712_CHIP_RAM.N_38\
        );

    \I__2124\ : IoInMux
    port map (
            O => \N__9129\,
            I => \N__9126\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__9126\,
            I => \N__9123\
        );

    \I__2122\ : IoSpan4Mux
    port map (
            O => \N__9123\,
            I => \N__9120\
        );

    \I__2121\ : Sp12to4
    port map (
            O => \N__9120\,
            I => \N__9117\
        );

    \I__2120\ : Span12Mux_s1_h
    port map (
            O => \N__9117\,
            I => \N__9114\
        );

    \I__2119\ : Span12Mux_h
    port map (
            O => \N__9114\,
            I => \N__9111\
        );

    \I__2118\ : Odrv12
    port map (
            O => \N__9111\,
            I => \CMA_c_7\
        );

    \I__2117\ : IoInMux
    port map (
            O => \N__9108\,
            I => \N__9105\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__9105\,
            I => \N__9102\
        );

    \I__2115\ : Span12Mux_s9_v
    port map (
            O => \N__9102\,
            I => \N__9099\
        );

    \I__2114\ : Odrv12
    port map (
            O => \N__9099\,
            I => \CMA_c_10\
        );

    \I__2113\ : CEMux
    port map (
            O => \N__9096\,
            I => \N__9092\
        );

    \I__2112\ : CEMux
    port map (
            O => \N__9095\,
            I => \N__9088\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__9092\,
            I => \N__9085\
        );

    \I__2110\ : CEMux
    port map (
            O => \N__9091\,
            I => \N__9082\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__9088\,
            I => \N__9077\
        );

    \I__2108\ : Span4Mux_h
    port map (
            O => \N__9085\,
            I => \N__9072\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__9082\,
            I => \N__9072\
        );

    \I__2106\ : CEMux
    port map (
            O => \N__9081\,
            I => \N__9069\
        );

    \I__2105\ : CEMux
    port map (
            O => \N__9080\,
            I => \N__9066\
        );

    \I__2104\ : Span4Mux_v
    port map (
            O => \N__9077\,
            I => \N__9057\
        );

    \I__2103\ : Span4Mux_v
    port map (
            O => \N__9072\,
            I => \N__9057\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__9069\,
            I => \N__9057\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9066\,
            I => \N__9054\
        );

    \I__2100\ : CEMux
    port map (
            O => \N__9065\,
            I => \N__9051\
        );

    \I__2099\ : CEMux
    port map (
            O => \N__9064\,
            I => \N__9048\
        );

    \I__2098\ : Span4Mux_h
    port map (
            O => \N__9057\,
            I => \N__9045\
        );

    \I__2097\ : Span4Mux_h
    port map (
            O => \N__9054\,
            I => \N__9042\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__9051\,
            I => \N__9037\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__9048\,
            I => \N__9037\
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__9045\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__2093\ : Odrv4
    port map (
            O => \N__9042\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__2092\ : Odrv12
    port map (
            O => \N__9037\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__9030\,
            I => \N__9025\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__9029\,
            I => \N__9022\
        );

    \I__2089\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9014\
        );

    \I__2088\ : InMux
    port map (
            O => \N__9025\,
            I => \N__9009\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9022\,
            I => \N__9009\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__9021\,
            I => \N__9006\
        );

    \I__2085\ : InMux
    port map (
            O => \N__9020\,
            I => \N__9002\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9019\,
            I => \N__8999\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9018\,
            I => \N__8994\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9017\,
            I => \N__8994\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__9014\,
            I => \N__8991\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9009\,
            I => \N__8988\
        );

    \I__2079\ : InMux
    port map (
            O => \N__9006\,
            I => \N__8981\
        );

    \I__2078\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8981\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__9002\,
            I => \N__8976\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__8999\,
            I => \N__8976\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__8994\,
            I => \N__8971\
        );

    \I__2074\ : Span4Mux_h
    port map (
            O => \N__8991\,
            I => \N__8971\
        );

    \I__2073\ : Span4Mux_h
    port map (
            O => \N__8988\,
            I => \N__8968\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__8987\,
            I => \N__8964\
        );

    \I__2071\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8959\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__8981\,
            I => \N__8956\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__8976\,
            I => \N__8951\
        );

    \I__2068\ : Span4Mux_v
    port map (
            O => \N__8971\,
            I => \N__8951\
        );

    \I__2067\ : Span4Mux_h
    port map (
            O => \N__8968\,
            I => \N__8948\
        );

    \I__2066\ : InMux
    port map (
            O => \N__8967\,
            I => \N__8945\
        );

    \I__2065\ : InMux
    port map (
            O => \N__8964\,
            I => \N__8942\
        );

    \I__2064\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8937\
        );

    \I__2063\ : InMux
    port map (
            O => \N__8962\,
            I => \N__8937\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__8959\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__8956\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__8951\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2059\ : Odrv4
    port map (
            O => \N__8948\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__8945\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__8942\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__8937\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\
        );

    \I__2055\ : IoInMux
    port map (
            O => \N__8922\,
            I => \N__8919\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__8919\,
            I => \N__8916\
        );

    \I__2053\ : Span4Mux_s3_h
    port map (
            O => \N__8916\,
            I => \N__8913\
        );

    \I__2052\ : Span4Mux_v
    port map (
            O => \N__8913\,
            I => \N__8910\
        );

    \I__2051\ : Span4Mux_h
    port map (
            O => \N__8910\,
            I => \N__8907\
        );

    \I__2050\ : Span4Mux_h
    port map (
            O => \N__8907\,
            I => \N__8904\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__8904\,
            I => \WEn_c\
        );

    \I__2048\ : InMux
    port map (
            O => \N__8901\,
            I => \N__8892\
        );

    \I__2047\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8887\
        );

    \I__2046\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8882\
        );

    \I__2045\ : InMux
    port map (
            O => \N__8898\,
            I => \N__8882\
        );

    \I__2044\ : InMux
    port map (
            O => \N__8897\,
            I => \N__8878\
        );

    \I__2043\ : InMux
    port map (
            O => \N__8896\,
            I => \N__8875\
        );

    \I__2042\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8872\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__8892\,
            I => \N__8869\
        );

    \I__2040\ : InMux
    port map (
            O => \N__8891\,
            I => \N__8864\
        );

    \I__2039\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8864\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__8887\,
            I => \N__8861\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__8882\,
            I => \N__8858\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__8881\,
            I => \N__8855\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__8878\,
            I => \N__8851\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__8875\,
            I => \N__8840\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__8872\,
            I => \N__8840\
        );

    \I__2032\ : Span4Mux_v
    port map (
            O => \N__8869\,
            I => \N__8840\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__8864\,
            I => \N__8840\
        );

    \I__2030\ : Span4Mux_h
    port map (
            O => \N__8861\,
            I => \N__8840\
        );

    \I__2029\ : Span4Mux_h
    port map (
            O => \N__8858\,
            I => \N__8837\
        );

    \I__2028\ : InMux
    port map (
            O => \N__8855\,
            I => \N__8831\
        );

    \I__2027\ : InMux
    port map (
            O => \N__8854\,
            I => \N__8828\
        );

    \I__2026\ : Span4Mux_v
    port map (
            O => \N__8851\,
            I => \N__8825\
        );

    \I__2025\ : Span4Mux_h
    port map (
            O => \N__8840\,
            I => \N__8822\
        );

    \I__2024\ : Span4Mux_h
    port map (
            O => \N__8837\,
            I => \N__8819\
        );

    \I__2023\ : InMux
    port map (
            O => \N__8836\,
            I => \N__8816\
        );

    \I__2022\ : InMux
    port map (
            O => \N__8835\,
            I => \N__8813\
        );

    \I__2021\ : InMux
    port map (
            O => \N__8834\,
            I => \N__8810\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__8831\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__8828\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__8825\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__8822\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__8819\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__8816\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__8813\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__8810\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__2012\ : IoInMux
    port map (
            O => \N__8793\,
            I => \N__8790\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__8790\,
            I => \N__8787\
        );

    \I__2010\ : Span4Mux_s3_v
    port map (
            O => \N__8787\,
            I => \N__8784\
        );

    \I__2009\ : Span4Mux_v
    port map (
            O => \N__8784\,
            I => \N__8781\
        );

    \I__2008\ : Span4Mux_h
    port map (
            O => \N__8781\,
            I => \N__8778\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__8778\,
            I => \RASn_c\
        );

    \I__2006\ : CEMux
    port map (
            O => \N__8775\,
            I => \N__8771\
        );

    \I__2005\ : CEMux
    port map (
            O => \N__8774\,
            I => \N__8766\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__8771\,
            I => \N__8762\
        );

    \I__2003\ : CEMux
    port map (
            O => \N__8770\,
            I => \N__8759\
        );

    \I__2002\ : CEMux
    port map (
            O => \N__8769\,
            I => \N__8756\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__8766\,
            I => \N__8753\
        );

    \I__2000\ : CEMux
    port map (
            O => \N__8765\,
            I => \N__8750\
        );

    \I__1999\ : Span4Mux_v
    port map (
            O => \N__8762\,
            I => \N__8747\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__8759\,
            I => \N__8744\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__8756\,
            I => \N__8741\
        );

    \I__1996\ : Span4Mux_v
    port map (
            O => \N__8753\,
            I => \N__8736\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__8750\,
            I => \N__8736\
        );

    \I__1994\ : Span4Mux_h
    port map (
            O => \N__8747\,
            I => \N__8731\
        );

    \I__1993\ : Span4Mux_v
    port map (
            O => \N__8744\,
            I => \N__8731\
        );

    \I__1992\ : Span4Mux_h
    port map (
            O => \N__8741\,
            I => \N__8728\
        );

    \I__1991\ : Span4Mux_h
    port map (
            O => \N__8736\,
            I => \N__8725\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__8731\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__8728\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__8725\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__8718\,
            I => \N__8711\
        );

    \I__1986\ : InMux
    port map (
            O => \N__8717\,
            I => \N__8705\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__8716\,
            I => \N__8702\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__8715\,
            I => \N__8699\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__8714\,
            I => \N__8695\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8711\,
            I => \N__8691\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__8710\,
            I => \N__8688\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__8709\,
            I => \N__8685\
        );

    \I__1979\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8682\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__8705\,
            I => \N__8679\
        );

    \I__1977\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8676\
        );

    \I__1976\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8673\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__8698\,
            I => \N__8670\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8695\,
            I => \N__8667\
        );

    \I__1973\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8663\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__8691\,
            I => \N__8660\
        );

    \I__1971\ : InMux
    port map (
            O => \N__8688\,
            I => \N__8657\
        );

    \I__1970\ : InMux
    port map (
            O => \N__8685\,
            I => \N__8654\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__8682\,
            I => \N__8645\
        );

    \I__1968\ : Span4Mux_v
    port map (
            O => \N__8679\,
            I => \N__8645\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__8676\,
            I => \N__8645\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__8673\,
            I => \N__8645\
        );

    \I__1965\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8642\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__8667\,
            I => \N__8637\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8634\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__8663\,
            I => \N__8630\
        );

    \I__1961\ : Span4Mux_v
    port map (
            O => \N__8660\,
            I => \N__8625\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8657\,
            I => \N__8625\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__8654\,
            I => \N__8620\
        );

    \I__1958\ : Span4Mux_h
    port map (
            O => \N__8645\,
            I => \N__8620\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__8642\,
            I => \N__8617\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__8641\,
            I => \N__8612\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8640\,
            I => \N__8609\
        );

    \I__1954\ : Span4Mux_v
    port map (
            O => \N__8637\,
            I => \N__8604\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__8634\,
            I => \N__8604\
        );

    \I__1952\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8601\
        );

    \I__1951\ : Span4Mux_h
    port map (
            O => \N__8630\,
            I => \N__8598\
        );

    \I__1950\ : Span4Mux_h
    port map (
            O => \N__8625\,
            I => \N__8591\
        );

    \I__1949\ : Span4Mux_h
    port map (
            O => \N__8620\,
            I => \N__8591\
        );

    \I__1948\ : Span4Mux_h
    port map (
            O => \N__8617\,
            I => \N__8591\
        );

    \I__1947\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8586\
        );

    \I__1946\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8586\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8612\,
            I => \N__8583\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__8609\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__8604\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__8601\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__8598\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__8591\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__8586\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__8583\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1937\ : IoInMux
    port map (
            O => \N__8568\,
            I => \N__8565\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8565\,
            I => \N__8562\
        );

    \I__1935\ : Span4Mux_s2_v
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__1934\ : Span4Mux_v
    port map (
            O => \N__8559\,
            I => \N__8556\
        );

    \I__1933\ : Span4Mux_h
    port map (
            O => \N__8556\,
            I => \N__8553\
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__8553\,
            I => \CASn_c\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8546\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8543\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__8546\,
            I => \N__8538\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__8543\,
            I => \N__8538\
        );

    \I__1927\ : Span12Mux_h
    port map (
            O => \N__8538\,
            I => \N__8532\
        );

    \I__1926\ : InMux
    port map (
            O => \N__8537\,
            I => \N__8529\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8536\,
            I => \N__8524\
        );

    \I__1924\ : InMux
    port map (
            O => \N__8535\,
            I => \N__8524\
        );

    \I__1923\ : Odrv12
    port map (
            O => \N__8532\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__8529\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__8524\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1920\ : IoInMux
    port map (
            O => \N__8517\,
            I => \N__8514\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__8514\,
            I => \N__8511\
        );

    \I__1918\ : Span4Mux_s1_v
    port map (
            O => \N__8511\,
            I => \N__8508\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__8508\,
            I => \N__8505\
        );

    \I__1916\ : Span4Mux_v
    port map (
            O => \N__8505\,
            I => \N__8502\
        );

    \I__1915\ : Odrv4
    port map (
            O => \N__8502\,
            I => \CRCSn_c\
        );

    \I__1914\ : InMux
    port map (
            O => \N__8499\,
            I => \N__8496\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8496\,
            I => \N__8493\
        );

    \I__1912\ : Span12Mux_h
    port map (
            O => \N__8493\,
            I => \N__8490\
        );

    \I__1911\ : Odrv12
    port map (
            O => \N__8490\,
            I => \RAS1n_c\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8487\,
            I => \N__8484\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__8484\,
            I => \N__8480\
        );

    \I__1908\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8477\
        );

    \I__1907\ : Span4Mux_h
    port map (
            O => \N__8480\,
            I => \N__8472\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__8477\,
            I => \N__8472\
        );

    \I__1905\ : Sp12to4
    port map (
            O => \N__8472\,
            I => \N__8469\
        );

    \I__1904\ : Span12Mux_v
    port map (
            O => \N__8469\,
            I => \N__8466\
        );

    \I__1903\ : Span12Mux_h
    port map (
            O => \N__8466\,
            I => \N__8463\
        );

    \I__1902\ : Odrv12
    port map (
            O => \N__8463\,
            I => \DRA_c_6\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8457\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__8457\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1899\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8451\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__8451\,
            I => \N__8447\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8444\
        );

    \I__1896\ : Span4Mux_v
    port map (
            O => \N__8447\,
            I => \N__8441\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__8444\,
            I => \N__8438\
        );

    \I__1894\ : Sp12to4
    port map (
            O => \N__8441\,
            I => \N__8435\
        );

    \I__1893\ : Sp12to4
    port map (
            O => \N__8438\,
            I => \N__8432\
        );

    \I__1892\ : Span12Mux_h
    port map (
            O => \N__8435\,
            I => \N__8429\
        );

    \I__1891\ : Span12Mux_v
    port map (
            O => \N__8432\,
            I => \N__8426\
        );

    \I__1890\ : Span12Mux_v
    port map (
            O => \N__8429\,
            I => \N__8423\
        );

    \I__1889\ : Span12Mux_h
    port map (
            O => \N__8426\,
            I => \N__8420\
        );

    \I__1888\ : Odrv12
    port map (
            O => \N__8423\,
            I => \DRA_c_3\
        );

    \I__1887\ : Odrv12
    port map (
            O => \N__8420\,
            I => \DRA_c_3\
        );

    \I__1886\ : InMux
    port map (
            O => \N__8415\,
            I => \N__8412\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8412\,
            I => \N__8409\
        );

    \I__1884\ : Span4Mux_h
    port map (
            O => \N__8409\,
            I => \N__8406\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__8406\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8403\,
            I => \N__8400\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__8400\,
            I => \N__8397\
        );

    \I__1880\ : Span4Mux_h
    port map (
            O => \N__8397\,
            I => \N__8394\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__8394\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__8391\,
            I => \N__8387\
        );

    \I__1877\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8384\
        );

    \I__1876\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8381\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8384\,
            I => \N__8364\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8381\,
            I => \N__8364\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8361\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8379\,
            I => \N__8358\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__8378\,
            I => \N__8353\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8350\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8347\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__8375\,
            I => \N__8340\
        );

    \I__1867\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8335\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8373\,
            I => \N__8335\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8372\,
            I => \N__8330\
        );

    \I__1864\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8330\
        );

    \I__1863\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8325\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8369\,
            I => \N__8325\
        );

    \I__1861\ : Span4Mux_h
    port map (
            O => \N__8364\,
            I => \N__8320\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8361\,
            I => \N__8315\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__8358\,
            I => \N__8315\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8311\
        );

    \I__1857\ : InMux
    port map (
            O => \N__8356\,
            I => \N__8308\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8305\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__8350\,
            I => \N__8302\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8347\,
            I => \N__8299\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8346\,
            I => \N__8295\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8345\,
            I => \N__8288\
        );

    \I__1851\ : InMux
    port map (
            O => \N__8344\,
            I => \N__8288\
        );

    \I__1850\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8288\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8340\,
            I => \N__8285\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8335\,
            I => \N__8278\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__8330\,
            I => \N__8278\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__8325\,
            I => \N__8278\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8324\,
            I => \N__8273\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8323\,
            I => \N__8273\
        );

    \I__1843\ : Span4Mux_v
    port map (
            O => \N__8320\,
            I => \N__8267\
        );

    \I__1842\ : Span4Mux_v
    port map (
            O => \N__8315\,
            I => \N__8267\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8314\,
            I => \N__8264\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8311\,
            I => \N__8253\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8308\,
            I => \N__8253\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8305\,
            I => \N__8253\
        );

    \I__1837\ : Span4Mux_v
    port map (
            O => \N__8302\,
            I => \N__8253\
        );

    \I__1836\ : Span4Mux_h
    port map (
            O => \N__8299\,
            I => \N__8253\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8298\,
            I => \N__8250\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8295\,
            I => \N__8241\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8288\,
            I => \N__8241\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8285\,
            I => \N__8241\
        );

    \I__1831\ : Span4Mux_h
    port map (
            O => \N__8278\,
            I => \N__8241\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8273\,
            I => \N__8236\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8272\,
            I => \N__8233\
        );

    \I__1828\ : Sp12to4
    port map (
            O => \N__8267\,
            I => \N__8228\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8264\,
            I => \N__8228\
        );

    \I__1826\ : Span4Mux_h
    port map (
            O => \N__8253\,
            I => \N__8225\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__8250\,
            I => \N__8220\
        );

    \I__1824\ : Span4Mux_h
    port map (
            O => \N__8241\,
            I => \N__8220\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8240\,
            I => \N__8215\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8239\,
            I => \N__8215\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__8236\,
            I => \CPU_CYCLEm\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8233\,
            I => \CPU_CYCLEm\
        );

    \I__1819\ : Odrv12
    port map (
            O => \N__8228\,
            I => \CPU_CYCLEm\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__8225\,
            I => \CPU_CYCLEm\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__8220\,
            I => \CPU_CYCLEm\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8215\,
            I => \CPU_CYCLEm\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8202\,
            I => \N__8199\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8199\,
            I => \N__8196\
        );

    \I__1813\ : Span12Mux_v
    port map (
            O => \N__8196\,
            I => \N__8193\
        );

    \I__1812\ : Span12Mux_h
    port map (
            O => \N__8193\,
            I => \N__8190\
        );

    \I__1811\ : Odrv12
    port map (
            O => \N__8190\,
            I => \A_c_16\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__8187\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_7_cascade_\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8184\,
            I => \N__8181\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8181\,
            I => \N__8178\
        );

    \I__1807\ : Span12Mux_v
    port map (
            O => \N__8178\,
            I => \N__8175\
        );

    \I__1806\ : Span12Mux_h
    port map (
            O => \N__8175\,
            I => \N__8172\
        );

    \I__1805\ : Odrv12
    port map (
            O => \N__8172\,
            I => \A_c_18\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8169\,
            I => \N__8165\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8168\,
            I => \N__8162\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8165\,
            I => \N__8159\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8162\,
            I => \N__8156\
        );

    \I__1800\ : Span4Mux_v
    port map (
            O => \N__8159\,
            I => \N__8153\
        );

    \I__1799\ : Span12Mux_v
    port map (
            O => \N__8156\,
            I => \N__8148\
        );

    \I__1798\ : Sp12to4
    port map (
            O => \N__8153\,
            I => \N__8148\
        );

    \I__1797\ : Span12Mux_h
    port map (
            O => \N__8148\,
            I => \N__8145\
        );

    \I__1796\ : Odrv12
    port map (
            O => \N__8145\,
            I => \DRA_c_8\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__8142\,
            I => \N__8139\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8136\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8136\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8133\,
            I => \N__8130\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__8130\,
            I => \N__8127\
        );

    \I__1790\ : Span4Mux_v
    port map (
            O => \N__8127\,
            I => \N__8123\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8120\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__8123\,
            I => \N__8117\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__8120\,
            I => \N__8114\
        );

    \I__1786\ : Sp12to4
    port map (
            O => \N__8117\,
            I => \N__8109\
        );

    \I__1785\ : Span12Mux_v
    port map (
            O => \N__8114\,
            I => \N__8109\
        );

    \I__1784\ : Span12Mux_h
    port map (
            O => \N__8109\,
            I => \N__8106\
        );

    \I__1783\ : Odrv12
    port map (
            O => \N__8106\,
            I => \DRA_c_7\
        );

    \I__1782\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8100\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__8100\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__1780\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8094\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8094\,
            I => \N__8090\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8087\
        );

    \I__1777\ : Span4Mux_v
    port map (
            O => \N__8090\,
            I => \N__8082\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8087\,
            I => \N__8082\
        );

    \I__1775\ : Span4Mux_h
    port map (
            O => \N__8082\,
            I => \N__8079\
        );

    \I__1774\ : Span4Mux_v
    port map (
            O => \N__8079\,
            I => \N__8076\
        );

    \I__1773\ : Sp12to4
    port map (
            O => \N__8076\,
            I => \N__8073\
        );

    \I__1772\ : Span12Mux_h
    port map (
            O => \N__8073\,
            I => \N__8070\
        );

    \I__1771\ : Span12Mux_v
    port map (
            O => \N__8070\,
            I => \N__8067\
        );

    \I__1770\ : Odrv12
    port map (
            O => \N__8067\,
            I => \DRA_c_0\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8061\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8061\,
            I => \N__8058\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__8058\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8055\,
            I => \N__8052\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8052\,
            I => \N__8049\
        );

    \I__1764\ : Span4Mux_v
    port map (
            O => \N__8049\,
            I => \N__8045\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8048\,
            I => \N__8042\
        );

    \I__1762\ : Sp12to4
    port map (
            O => \N__8045\,
            I => \N__8039\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8042\,
            I => \N__8036\
        );

    \I__1760\ : Span12Mux_h
    port map (
            O => \N__8039\,
            I => \N__8033\
        );

    \I__1759\ : Span12Mux_v
    port map (
            O => \N__8036\,
            I => \N__8030\
        );

    \I__1758\ : Span12Mux_v
    port map (
            O => \N__8033\,
            I => \N__8027\
        );

    \I__1757\ : Span12Mux_h
    port map (
            O => \N__8030\,
            I => \N__8024\
        );

    \I__1756\ : Odrv12
    port map (
            O => \N__8027\,
            I => \DRA_c_2\
        );

    \I__1755\ : Odrv12
    port map (
            O => \N__8024\,
            I => \DRA_c_2\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8019\,
            I => \N__8016\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__8016\,
            I => \N__8013\
        );

    \I__1752\ : Span4Mux_h
    port map (
            O => \N__8013\,
            I => \N__8010\
        );

    \I__1751\ : Odrv4
    port map (
            O => \N__8010\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8007\,
            I => \N__8004\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__8004\,
            I => \N__7988\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8003\,
            I => \N__7983\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8002\,
            I => \N__7983\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8001\,
            I => \N__7978\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8000\,
            I => \N__7973\
        );

    \I__1744\ : InMux
    port map (
            O => \N__7999\,
            I => \N__7973\
        );

    \I__1743\ : InMux
    port map (
            O => \N__7998\,
            I => \N__7968\
        );

    \I__1742\ : InMux
    port map (
            O => \N__7997\,
            I => \N__7968\
        );

    \I__1741\ : InMux
    port map (
            O => \N__7996\,
            I => \N__7959\
        );

    \I__1740\ : InMux
    port map (
            O => \N__7995\,
            I => \N__7956\
        );

    \I__1739\ : InMux
    port map (
            O => \N__7994\,
            I => \N__7949\
        );

    \I__1738\ : InMux
    port map (
            O => \N__7993\,
            I => \N__7949\
        );

    \I__1737\ : InMux
    port map (
            O => \N__7992\,
            I => \N__7949\
        );

    \I__1736\ : InMux
    port map (
            O => \N__7991\,
            I => \N__7946\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__7988\,
            I => \N__7941\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__7983\,
            I => \N__7941\
        );

    \I__1733\ : InMux
    port map (
            O => \N__7982\,
            I => \N__7938\
        );

    \I__1732\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7934\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__7978\,
            I => \N__7929\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__7973\,
            I => \N__7929\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__7968\,
            I => \N__7926\
        );

    \I__1728\ : InMux
    port map (
            O => \N__7967\,
            I => \N__7923\
        );

    \I__1727\ : InMux
    port map (
            O => \N__7966\,
            I => \N__7912\
        );

    \I__1726\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7912\
        );

    \I__1725\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7912\
        );

    \I__1724\ : InMux
    port map (
            O => \N__7963\,
            I => \N__7912\
        );

    \I__1723\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7912\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__7959\,
            I => \N__7909\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__7956\,
            I => \N__7906\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__7949\,
            I => \N__7901\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__7946\,
            I => \N__7901\
        );

    \I__1718\ : Span4Mux_v
    port map (
            O => \N__7941\,
            I => \N__7894\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__7938\,
            I => \N__7891\
        );

    \I__1716\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7888\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__7934\,
            I => \N__7885\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__7929\,
            I => \N__7876\
        );

    \I__1713\ : Span4Mux_h
    port map (
            O => \N__7926\,
            I => \N__7876\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__7923\,
            I => \N__7876\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__7912\,
            I => \N__7876\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__7909\,
            I => \N__7873\
        );

    \I__1709\ : Span4Mux_h
    port map (
            O => \N__7906\,
            I => \N__7868\
        );

    \I__1708\ : Span4Mux_v
    port map (
            O => \N__7901\,
            I => \N__7868\
        );

    \I__1707\ : InMux
    port map (
            O => \N__7900\,
            I => \N__7861\
        );

    \I__1706\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7861\
        );

    \I__1705\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7861\
        );

    \I__1704\ : InMux
    port map (
            O => \N__7897\,
            I => \N__7858\
        );

    \I__1703\ : Span4Mux_h
    port map (
            O => \N__7894\,
            I => \N__7851\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__7891\,
            I => \N__7851\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__7888\,
            I => \N__7851\
        );

    \I__1700\ : Span4Mux_v
    port map (
            O => \N__7885\,
            I => \N__7846\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__7876\,
            I => \N__7846\
        );

    \I__1698\ : Span4Mux_h
    port map (
            O => \N__7873\,
            I => \N__7841\
        );

    \I__1697\ : Span4Mux_v
    port map (
            O => \N__7868\,
            I => \N__7841\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__7861\,
            I => \N__7838\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__7858\,
            I => \N__7833\
        );

    \I__1694\ : Sp12to4
    port map (
            O => \N__7851\,
            I => \N__7833\
        );

    \I__1693\ : Sp12to4
    port map (
            O => \N__7846\,
            I => \N__7830\
        );

    \I__1692\ : Sp12to4
    port map (
            O => \N__7841\,
            I => \N__7823\
        );

    \I__1691\ : Span12Mux_h
    port map (
            O => \N__7838\,
            I => \N__7823\
        );

    \I__1690\ : Span12Mux_v
    port map (
            O => \N__7833\,
            I => \N__7823\
        );

    \I__1689\ : Span12Mux_h
    port map (
            O => \N__7830\,
            I => \N__7820\
        );

    \I__1688\ : Span12Mux_h
    port map (
            O => \N__7823\,
            I => \N__7817\
        );

    \I__1687\ : Odrv12
    port map (
            O => \N__7820\,
            I => \RESETn_c\
        );

    \I__1686\ : Odrv12
    port map (
            O => \N__7817\,
            I => \RESETn_c\
        );

    \I__1685\ : IoInMux
    port map (
            O => \N__7812\,
            I => \N__7809\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__7809\,
            I => \N__7806\
        );

    \I__1683\ : Odrv12
    port map (
            O => \N__7806\,
            I => \RESETn_c_i\
        );

    \I__1682\ : IoInMux
    port map (
            O => \N__7803\,
            I => \N__7800\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__7800\,
            I => \N__7797\
        );

    \I__1680\ : Span4Mux_s2_v
    port map (
            O => \N__7797\,
            I => \N__7794\
        );

    \I__1679\ : Span4Mux_v
    port map (
            O => \N__7794\,
            I => \N__7791\
        );

    \I__1678\ : Span4Mux_h
    port map (
            O => \N__7791\,
            I => \N__7788\
        );

    \I__1677\ : Odrv4
    port map (
            O => \N__7788\,
            I => \CMA_c_0\
        );

    \I__1676\ : InMux
    port map (
            O => \N__7785\,
            I => \N__7782\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__7782\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__1674\ : IoInMux
    port map (
            O => \N__7779\,
            I => \N__7776\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__7776\,
            I => \N__7773\
        );

    \I__1672\ : IoSpan4Mux
    port map (
            O => \N__7773\,
            I => \N__7770\
        );

    \I__1671\ : IoSpan4Mux
    port map (
            O => \N__7770\,
            I => \N__7767\
        );

    \I__1670\ : Span4Mux_s3_h
    port map (
            O => \N__7767\,
            I => \N__7764\
        );

    \I__1669\ : Span4Mux_h
    port map (
            O => \N__7764\,
            I => \N__7761\
        );

    \I__1668\ : Span4Mux_h
    port map (
            O => \N__7761\,
            I => \N__7758\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__7758\,
            I => \CMA_c_5\
        );

    \I__1666\ : InMux
    port map (
            O => \N__7755\,
            I => \N__7752\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__7752\,
            I => \N__7749\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__7749\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1663\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7743\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7743\,
            I => \N__7740\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__7740\,
            I => \N__7737\
        );

    \I__1660\ : Span4Mux_v
    port map (
            O => \N__7737\,
            I => \N__7734\
        );

    \I__1659\ : Sp12to4
    port map (
            O => \N__7734\,
            I => \N__7731\
        );

    \I__1658\ : Span12Mux_h
    port map (
            O => \N__7731\,
            I => \N__7728\
        );

    \I__1657\ : Odrv12
    port map (
            O => \N__7728\,
            I => \A_c_9\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__7725\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_\
        );

    \I__1655\ : InMux
    port map (
            O => \N__7722\,
            I => \N__7719\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__7719\,
            I => \N__7716\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__7716\,
            I => \N__7713\
        );

    \I__1652\ : Span4Mux_v
    port map (
            O => \N__7713\,
            I => \N__7710\
        );

    \I__1651\ : Sp12to4
    port map (
            O => \N__7710\,
            I => \N__7707\
        );

    \I__1650\ : Span12Mux_h
    port map (
            O => \N__7707\,
            I => \N__7704\
        );

    \I__1649\ : Span12Mux_v
    port map (
            O => \N__7704\,
            I => \N__7701\
        );

    \I__1648\ : Odrv12
    port map (
            O => \N__7701\,
            I => \A_c_2\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7698\,
            I => \N__7695\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__7695\,
            I => \U712_CHIP_RAM.N_31\
        );

    \I__1645\ : InMux
    port map (
            O => \N__7692\,
            I => \N__7689\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7689\,
            I => \N__7686\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__7686\,
            I => \N__7683\
        );

    \I__1642\ : Span4Mux_v
    port map (
            O => \N__7683\,
            I => \N__7680\
        );

    \I__1641\ : Sp12to4
    port map (
            O => \N__7680\,
            I => \N__7677\
        );

    \I__1640\ : Span12Mux_h
    port map (
            O => \N__7677\,
            I => \N__7674\
        );

    \I__1639\ : Odrv12
    port map (
            O => \N__7674\,
            I => \A_c_17\
        );

    \I__1638\ : IoInMux
    port map (
            O => \N__7671\,
            I => \N__7668\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__7668\,
            I => \N__7665\
        );

    \I__1636\ : IoSpan4Mux
    port map (
            O => \N__7665\,
            I => \N__7662\
        );

    \I__1635\ : Span4Mux_s1_h
    port map (
            O => \N__7662\,
            I => \N__7659\
        );

    \I__1634\ : Sp12to4
    port map (
            O => \N__7659\,
            I => \N__7656\
        );

    \I__1633\ : Span12Mux_h
    port map (
            O => \N__7656\,
            I => \N__7653\
        );

    \I__1632\ : Odrv12
    port map (
            O => \N__7653\,
            I => \CMA_c_8\
        );

    \I__1631\ : IoInMux
    port map (
            O => \N__7650\,
            I => \N__7647\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__7647\,
            I => \N__7644\
        );

    \I__1629\ : Span12Mux_s3_h
    port map (
            O => \N__7644\,
            I => \N__7641\
        );

    \I__1628\ : Span12Mux_h
    port map (
            O => \N__7641\,
            I => \N__7638\
        );

    \I__1627\ : Odrv12
    port map (
            O => \N__7638\,
            I => \CMA_c_6\
        );

    \I__1626\ : InMux
    port map (
            O => \N__7635\,
            I => \N__7631\
        );

    \I__1625\ : InMux
    port map (
            O => \N__7634\,
            I => \N__7628\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7631\,
            I => \N__7625\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7628\,
            I => \N__7622\
        );

    \I__1622\ : Span4Mux_h
    port map (
            O => \N__7625\,
            I => \N__7619\
        );

    \I__1621\ : Odrv12
    port map (
            O => \N__7622\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1620\ : Odrv4
    port map (
            O => \N__7619\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__7614\,
            I => \N__7611\
        );

    \I__1618\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7608\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__7608\,
            I => \N__7605\
        );

    \I__1616\ : Span4Mux_v
    port map (
            O => \N__7605\,
            I => \N__7602\
        );

    \I__1615\ : Span4Mux_v
    port map (
            O => \N__7602\,
            I => \N__7599\
        );

    \I__1614\ : Sp12to4
    port map (
            O => \N__7599\,
            I => \N__7596\
        );

    \I__1613\ : Span12Mux_h
    port map (
            O => \N__7596\,
            I => \N__7593\
        );

    \I__1612\ : Odrv12
    port map (
            O => \N__7593\,
            I => \A_c_19\
        );

    \I__1611\ : IoInMux
    port map (
            O => \N__7590\,
            I => \N__7587\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7587\,
            I => \N__7584\
        );

    \I__1609\ : Span12Mux_s3_h
    port map (
            O => \N__7584\,
            I => \N__7581\
        );

    \I__1608\ : Span12Mux_h
    port map (
            O => \N__7581\,
            I => \N__7578\
        );

    \I__1607\ : Odrv12
    port map (
            O => \N__7578\,
            I => \CMA_c_9\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7575\,
            I => \N__7572\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__7572\,
            I => \N__7569\
        );

    \I__1604\ : Span4Mux_v
    port map (
            O => \N__7569\,
            I => \N__7566\
        );

    \I__1603\ : Span4Mux_v
    port map (
            O => \N__7566\,
            I => \N__7563\
        );

    \I__1602\ : Sp12to4
    port map (
            O => \N__7563\,
            I => \N__7560\
        );

    \I__1601\ : Span12Mux_h
    port map (
            O => \N__7560\,
            I => \N__7557\
        );

    \I__1600\ : Odrv12
    port map (
            O => \N__7557\,
            I => \A_c_15\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7554\,
            I => \N__7551\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7551\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_6\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__7548\,
            I => \N__7545\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7542\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7542\,
            I => \N__7539\
        );

    \I__1594\ : Span4Mux_h
    port map (
            O => \N__7539\,
            I => \N__7536\
        );

    \I__1593\ : Span4Mux_v
    port map (
            O => \N__7536\,
            I => \N__7533\
        );

    \I__1592\ : Sp12to4
    port map (
            O => \N__7533\,
            I => \N__7530\
        );

    \I__1591\ : Span12Mux_h
    port map (
            O => \N__7530\,
            I => \N__7527\
        );

    \I__1590\ : Odrv12
    port map (
            O => \N__7527\,
            I => \A_c_8\
        );

    \I__1589\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7521\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__7521\,
            I => \U712_CHIP_RAM.N_37\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7518\,
            I => \N__7514\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7517\,
            I => \N__7511\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7514\,
            I => \N__7506\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7511\,
            I => \N__7506\
        );

    \I__1583\ : Sp12to4
    port map (
            O => \N__7506\,
            I => \N__7503\
        );

    \I__1582\ : Span12Mux_v
    port map (
            O => \N__7503\,
            I => \N__7500\
        );

    \I__1581\ : Span12Mux_h
    port map (
            O => \N__7500\,
            I => \N__7497\
        );

    \I__1580\ : Odrv12
    port map (
            O => \N__7497\,
            I => \DRA_c_4\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7494\,
            I => \N__7491\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__7491\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7488\,
            I => \N__7484\
        );

    \I__1576\ : InMux
    port map (
            O => \N__7487\,
            I => \N__7481\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7484\,
            I => \N__7478\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__7481\,
            I => \N__7475\
        );

    \I__1573\ : Span4Mux_v
    port map (
            O => \N__7478\,
            I => \N__7472\
        );

    \I__1572\ : Span4Mux_h
    port map (
            O => \N__7475\,
            I => \N__7469\
        );

    \I__1571\ : Sp12to4
    port map (
            O => \N__7472\,
            I => \N__7466\
        );

    \I__1570\ : Sp12to4
    port map (
            O => \N__7469\,
            I => \N__7463\
        );

    \I__1569\ : Span12Mux_h
    port map (
            O => \N__7466\,
            I => \N__7460\
        );

    \I__1568\ : Span12Mux_v
    port map (
            O => \N__7463\,
            I => \N__7457\
        );

    \I__1567\ : Span12Mux_v
    port map (
            O => \N__7460\,
            I => \N__7452\
        );

    \I__1566\ : Span12Mux_h
    port map (
            O => \N__7457\,
            I => \N__7452\
        );

    \I__1565\ : Odrv12
    port map (
            O => \N__7452\,
            I => \DRA_c_5\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7449\,
            I => \N__7446\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__7446\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7443\,
            I => \N__7440\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7440\,
            I => \U712_CHIP_RAM.N_32\
        );

    \I__1560\ : IoInMux
    port map (
            O => \N__7437\,
            I => \N__7434\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7434\,
            I => \N__7431\
        );

    \I__1558\ : Span12Mux_s8_v
    port map (
            O => \N__7431\,
            I => \N__7428\
        );

    \I__1557\ : Odrv12
    port map (
            O => \N__7428\,
            I => \CMA_c_1\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7425\,
            I => \N__7422\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7422\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7416\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__7416\,
            I => \N__7413\
        );

    \I__1552\ : Odrv12
    port map (
            O => \N__7413\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1551\ : CEMux
    port map (
            O => \N__7410\,
            I => \N__7406\
        );

    \I__1550\ : CEMux
    port map (
            O => \N__7409\,
            I => \N__7403\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7406\,
            I => \N__7400\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7403\,
            I => \N__7397\
        );

    \I__1547\ : Odrv12
    port map (
            O => \N__7400\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1546\ : Odrv12
    port map (
            O => \N__7397\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1545\ : InMux
    port map (
            O => \N__7392\,
            I => \N__7389\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7389\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7382\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7379\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__7382\,
            I => \N__7373\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7379\,
            I => \N__7373\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7378\,
            I => \N__7370\
        );

    \I__1538\ : Span4Mux_v
    port map (
            O => \N__7373\,
            I => \N__7367\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__7370\,
            I => \N__7364\
        );

    \I__1536\ : Sp12to4
    port map (
            O => \N__7367\,
            I => \N__7361\
        );

    \I__1535\ : Span12Mux_h
    port map (
            O => \N__7364\,
            I => \N__7358\
        );

    \I__1534\ : Span12Mux_h
    port map (
            O => \N__7361\,
            I => \N__7355\
        );

    \I__1533\ : Span12Mux_v
    port map (
            O => \N__7358\,
            I => \N__7352\
        );

    \I__1532\ : Span12Mux_v
    port map (
            O => \N__7355\,
            I => \N__7349\
        );

    \I__1531\ : Odrv12
    port map (
            O => \N__7352\,
            I => \CASLn_c\
        );

    \I__1530\ : Odrv12
    port map (
            O => \N__7349\,
            I => \CASLn_c\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7344\,
            I => \N__7341\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7341\,
            I => \N__7338\
        );

    \I__1527\ : Span4Mux_v
    port map (
            O => \N__7338\,
            I => \N__7333\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7337\,
            I => \N__7330\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7327\
        );

    \I__1524\ : Sp12to4
    port map (
            O => \N__7333\,
            I => \N__7320\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7330\,
            I => \N__7320\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7327\,
            I => \N__7320\
        );

    \I__1521\ : Span12Mux_h
    port map (
            O => \N__7320\,
            I => \N__7317\
        );

    \I__1520\ : Span12Mux_v
    port map (
            O => \N__7317\,
            I => \N__7314\
        );

    \I__1519\ : Odrv12
    port map (
            O => \N__7314\,
            I => \CASUn_c\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7311\,
            I => \N__7307\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7310\,
            I => \N__7304\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__7307\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__7304\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7299\,
            I => \N__7296\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7296\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7290\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7290\,
            I => \N__7286\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7289\,
            I => \N__7283\
        );

    \I__1509\ : Odrv4
    port map (
            O => \N__7286\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7283\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7278\,
            I => \N__7274\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7277\,
            I => \N__7271\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7274\,
            I => \N__7266\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7271\,
            I => \N__7266\
        );

    \I__1503\ : Span4Mux_v
    port map (
            O => \N__7266\,
            I => \N__7262\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7265\,
            I => \N__7259\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__7262\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7259\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__1499\ : IoInMux
    port map (
            O => \N__7254\,
            I => \N__7251\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7251\,
            I => \N__7248\
        );

    \I__1497\ : Span12Mux_s4_v
    port map (
            O => \N__7248\,
            I => \N__7245\
        );

    \I__1496\ : Span12Mux_h
    port map (
            O => \N__7245\,
            I => \N__7242\
        );

    \I__1495\ : Odrv12
    port map (
            O => \N__7242\,
            I => \U712_REG_SM_un1_UDSn_i\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7239\,
            I => \N__7235\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__7238\,
            I => \N__7230\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7235\,
            I => \N__7226\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7234\,
            I => \N__7218\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7233\,
            I => \N__7218\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7230\,
            I => \N__7218\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7229\,
            I => \N__7215\
        );

    \I__1487\ : Span4Mux_v
    port map (
            O => \N__7226\,
            I => \N__7211\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7225\,
            I => \N__7208\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7218\,
            I => \N__7205\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7215\,
            I => \N__7202\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7199\
        );

    \I__1482\ : Span4Mux_v
    port map (
            O => \N__7211\,
            I => \N__7194\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7208\,
            I => \N__7194\
        );

    \I__1480\ : Odrv12
    port map (
            O => \N__7205\,
            I => \DMA_CYCLEm\
        );

    \I__1479\ : Odrv4
    port map (
            O => \N__7202\,
            I => \DMA_CYCLEm\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7199\,
            I => \DMA_CYCLEm\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__7194\,
            I => \DMA_CYCLEm\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7185\,
            I => \N__7181\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7184\,
            I => \N__7178\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7181\,
            I => \N__7175\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7178\,
            I => \N__7172\
        );

    \I__1472\ : Span4Mux_v
    port map (
            O => \N__7175\,
            I => \N__7167\
        );

    \I__1471\ : Span4Mux_v
    port map (
            O => \N__7172\,
            I => \N__7164\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7171\,
            I => \N__7161\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7170\,
            I => \N__7158\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__7167\,
            I => \REG_CYCLEm\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__7164\,
            I => \REG_CYCLEm\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7161\,
            I => \REG_CYCLEm\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7158\,
            I => \REG_CYCLEm\
        );

    \I__1464\ : IoInMux
    port map (
            O => \N__7149\,
            I => \N__7146\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7146\,
            I => \N__7143\
        );

    \I__1462\ : Span4Mux_s3_v
    port map (
            O => \N__7143\,
            I => \N__7140\
        );

    \I__1461\ : Span4Mux_h
    port map (
            O => \N__7140\,
            I => \N__7137\
        );

    \I__1460\ : Sp12to4
    port map (
            O => \N__7137\,
            I => \N__7134\
        );

    \I__1459\ : Span12Mux_v
    port map (
            O => \N__7134\,
            I => \N__7131\
        );

    \I__1458\ : Span12Mux_h
    port map (
            O => \N__7131\,
            I => \N__7128\
        );

    \I__1457\ : Odrv12
    port map (
            O => \N__7128\,
            I => \DRDENn_c\
        );

    \I__1456\ : IoInMux
    port map (
            O => \N__7125\,
            I => \N__7122\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7122\,
            I => \N__7119\
        );

    \I__1454\ : Span4Mux_s2_v
    port map (
            O => \N__7119\,
            I => \N__7116\
        );

    \I__1453\ : Span4Mux_v
    port map (
            O => \N__7116\,
            I => \N__7113\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__7113\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7110\,
            I => \N__7107\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__7107\,
            I => \N__7104\
        );

    \I__1449\ : Span4Mux_v
    port map (
            O => \N__7104\,
            I => \N__7101\
        );

    \I__1448\ : Sp12to4
    port map (
            O => \N__7101\,
            I => \N__7098\
        );

    \I__1447\ : Span12Mux_h
    port map (
            O => \N__7098\,
            I => \N__7095\
        );

    \I__1446\ : Odrv12
    port map (
            O => \N__7095\,
            I => \A_c_14\
        );

    \I__1445\ : CascadeMux
    port map (
            O => \N__7092\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_5_cascade_\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7089\,
            I => \N__7086\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7086\,
            I => \N__7083\
        );

    \I__1442\ : Span12Mux_v
    port map (
            O => \N__7083\,
            I => \N__7080\
        );

    \I__1441\ : Span12Mux_h
    port map (
            O => \N__7080\,
            I => \N__7077\
        );

    \I__1440\ : Odrv12
    port map (
            O => \N__7077\,
            I => \A_c_7\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7071\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__7071\,
            I => \N__7068\
        );

    \I__1437\ : Odrv4
    port map (
            O => \N__7068\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7065\,
            I => \N__7062\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__7062\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7059\,
            I => \N__7056\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7056\,
            I => \N__7053\
        );

    \I__1432\ : Span4Mux_v
    port map (
            O => \N__7053\,
            I => \N__7050\
        );

    \I__1431\ : Sp12to4
    port map (
            O => \N__7050\,
            I => \N__7047\
        );

    \I__1430\ : Span12Mux_h
    port map (
            O => \N__7047\,
            I => \N__7044\
        );

    \I__1429\ : Odrv12
    port map (
            O => \N__7044\,
            I => \A_c_10\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__7041\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7038\,
            I => \N__7035\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__7035\,
            I => \N__7032\
        );

    \I__1425\ : Span12Mux_h
    port map (
            O => \N__7032\,
            I => \N__7029\
        );

    \I__1424\ : Span12Mux_v
    port map (
            O => \N__7029\,
            I => \N__7026\
        );

    \I__1423\ : Odrv12
    port map (
            O => \N__7026\,
            I => \A_c_3\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7023\,
            I => \N__7020\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7020\,
            I => \N__7017\
        );

    \I__1420\ : Odrv12
    port map (
            O => \N__7017\,
            I => \U712_CHIP_RAM.DBENn_7_0_a2_0\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7014\,
            I => \N__7011\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__7011\,
            I => \N__7007\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7010\,
            I => \N__7004\
        );

    \I__1416\ : Span4Mux_v
    port map (
            O => \N__7007\,
            I => \N__7001\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__7004\,
            I => \N__6998\
        );

    \I__1414\ : Span4Mux_h
    port map (
            O => \N__7001\,
            I => \N__6993\
        );

    \I__1413\ : Span4Mux_v
    port map (
            O => \N__6998\,
            I => \N__6993\
        );

    \I__1412\ : Span4Mux_h
    port map (
            O => \N__6993\,
            I => \N__6990\
        );

    \I__1411\ : Sp12to4
    port map (
            O => \N__6990\,
            I => \N__6986\
        );

    \I__1410\ : IoInMux
    port map (
            O => \N__6989\,
            I => \N__6983\
        );

    \I__1409\ : Span12Mux_v
    port map (
            O => \N__6986\,
            I => \N__6980\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__6983\,
            I => \N__6977\
        );

    \I__1407\ : Odrv12
    port map (
            O => \N__6980\,
            I => \AWEn_c\
        );

    \I__1406\ : Odrv4
    port map (
            O => \N__6977\,
            I => \AWEn_c\
        );

    \I__1405\ : InMux
    port map (
            O => \N__6972\,
            I => \N__6968\
        );

    \I__1404\ : InMux
    port map (
            O => \N__6971\,
            I => \N__6965\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__6968\,
            I => \N__6959\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__6965\,
            I => \N__6956\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__6964\,
            I => \N__6953\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__6963\,
            I => \N__6950\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6962\,
            I => \N__6947\
        );

    \I__1398\ : Span4Mux_v
    port map (
            O => \N__6959\,
            I => \N__6944\
        );

    \I__1397\ : Span4Mux_v
    port map (
            O => \N__6956\,
            I => \N__6941\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6953\,
            I => \N__6938\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6950\,
            I => \N__6935\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6947\,
            I => \N__6932\
        );

    \I__1393\ : Sp12to4
    port map (
            O => \N__6944\,
            I => \N__6923\
        );

    \I__1392\ : Sp12to4
    port map (
            O => \N__6941\,
            I => \N__6923\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6938\,
            I => \N__6923\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6935\,
            I => \N__6923\
        );

    \I__1389\ : Span12Mux_v
    port map (
            O => \N__6932\,
            I => \N__6920\
        );

    \I__1388\ : Span12Mux_h
    port map (
            O => \N__6923\,
            I => \N__6917\
        );

    \I__1387\ : Span12Mux_h
    port map (
            O => \N__6920\,
            I => \N__6914\
        );

    \I__1386\ : Span12Mux_v
    port map (
            O => \N__6917\,
            I => \N__6911\
        );

    \I__1385\ : Odrv12
    port map (
            O => \N__6914\,
            I => \RnW_c\
        );

    \I__1384\ : Odrv12
    port map (
            O => \N__6911\,
            I => \RnW_c\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6906\,
            I => \N__6900\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6905\,
            I => \N__6897\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6904\,
            I => \N__6891\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6903\,
            I => \N__6888\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6900\,
            I => \N__6883\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6897\,
            I => \N__6883\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6896\,
            I => \N__6878\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6895\,
            I => \N__6878\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6894\,
            I => \N__6875\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__6891\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__6888\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1372\ : Odrv4
    port map (
            O => \N__6883\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6878\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__6875\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6864\,
            I => \N__6861\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__6861\,
            I => \N__6857\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6860\,
            I => \N__6854\
        );

    \I__1366\ : Span4Mux_h
    port map (
            O => \N__6857\,
            I => \N__6851\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__6854\,
            I => \N__6848\
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__6851\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1363\ : Odrv4
    port map (
            O => \N__6848\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1362\ : CEMux
    port map (
            O => \N__6843\,
            I => \N__6840\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6840\,
            I => \N__6837\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__6837\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0\
        );

    \I__1359\ : InMux
    port map (
            O => \N__6834\,
            I => \N__6831\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__6831\,
            I => \N__6827\
        );

    \I__1357\ : InMux
    port map (
            O => \N__6830\,
            I => \N__6824\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__6827\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__6824\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1354\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6813\
        );

    \I__1353\ : InMux
    port map (
            O => \N__6818\,
            I => \N__6806\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6817\,
            I => \N__6806\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6816\,
            I => \N__6806\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6813\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6806\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6801\,
            I => \N__6798\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__6798\,
            I => \N__6795\
        );

    \I__1346\ : Span12Mux_v
    port map (
            O => \N__6795\,
            I => \N__6792\
        );

    \I__1345\ : Odrv12
    port map (
            O => \N__6792\,
            I => \TACK_EN_i_ess\
        );

    \I__1344\ : CEMux
    port map (
            O => \N__6789\,
            I => \N__6786\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__6786\,
            I => \U712_CYCLE_TERM.N_45_0_0_en_0\
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__6783\,
            I => \N__6780\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6780\,
            I => \N__6776\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6779\,
            I => \N__6773\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__6776\,
            I => \N__6768\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6773\,
            I => \N__6768\
        );

    \I__1337\ : Odrv12
    port map (
            O => \N__6768\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6765\,
            I => \N__6762\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__6762\,
            I => \U712_CHIP_RAM.N_33\
        );

    \I__1334\ : IoInMux
    port map (
            O => \N__6759\,
            I => \N__6756\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__6756\,
            I => \N__6753\
        );

    \I__1332\ : Span12Mux_s2_v
    port map (
            O => \N__6753\,
            I => \N__6750\
        );

    \I__1331\ : Odrv12
    port map (
            O => \N__6750\,
            I => \CMA_c_2\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6744\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6744\,
            I => \N__6741\
        );

    \I__1328\ : Span4Mux_v
    port map (
            O => \N__6741\,
            I => \N__6738\
        );

    \I__1327\ : Sp12to4
    port map (
            O => \N__6738\,
            I => \N__6735\
        );

    \I__1326\ : Span12Mux_h
    port map (
            O => \N__6735\,
            I => \N__6732\
        );

    \I__1325\ : Odrv12
    port map (
            O => \N__6732\,
            I => \A_c_13\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__6729\,
            I => \N__6726\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6726\,
            I => \N__6723\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6723\,
            I => \N__6720\
        );

    \I__1321\ : Span4Mux_v
    port map (
            O => \N__6720\,
            I => \N__6717\
        );

    \I__1320\ : Sp12to4
    port map (
            O => \N__6717\,
            I => \N__6714\
        );

    \I__1319\ : Span12Mux_h
    port map (
            O => \N__6714\,
            I => \N__6711\
        );

    \I__1318\ : Span12Mux_v
    port map (
            O => \N__6711\,
            I => \N__6708\
        );

    \I__1317\ : Odrv12
    port map (
            O => \N__6708\,
            I => \A_c_6\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__6705\,
            I => \U712_CHIP_RAM.N_35_cascade_\
        );

    \I__1315\ : IoInMux
    port map (
            O => \N__6702\,
            I => \N__6699\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__6699\,
            I => \N__6696\
        );

    \I__1313\ : IoSpan4Mux
    port map (
            O => \N__6696\,
            I => \N__6693\
        );

    \I__1312\ : IoSpan4Mux
    port map (
            O => \N__6693\,
            I => \N__6690\
        );

    \I__1311\ : Span4Mux_s2_h
    port map (
            O => \N__6690\,
            I => \N__6687\
        );

    \I__1310\ : Span4Mux_h
    port map (
            O => \N__6687\,
            I => \N__6684\
        );

    \I__1309\ : Sp12to4
    port map (
            O => \N__6684\,
            I => \N__6681\
        );

    \I__1308\ : Odrv12
    port map (
            O => \N__6681\,
            I => \CMA_c_4\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6675\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6675\,
            I => \N__6672\
        );

    \I__1305\ : Span4Mux_v
    port map (
            O => \N__6672\,
            I => \N__6669\
        );

    \I__1304\ : Sp12to4
    port map (
            O => \N__6669\,
            I => \N__6666\
        );

    \I__1303\ : Span12Mux_h
    port map (
            O => \N__6666\,
            I => \N__6663\
        );

    \I__1302\ : Odrv12
    port map (
            O => \N__6663\,
            I => \A_c_12\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__6660\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6657\,
            I => \N__6654\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6654\,
            I => \N__6651\
        );

    \I__1298\ : Sp12to4
    port map (
            O => \N__6651\,
            I => \N__6648\
        );

    \I__1297\ : Span12Mux_v
    port map (
            O => \N__6648\,
            I => \N__6645\
        );

    \I__1296\ : Span12Mux_h
    port map (
            O => \N__6645\,
            I => \N__6642\
        );

    \I__1295\ : Odrv12
    port map (
            O => \N__6642\,
            I => \A_c_5\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6639\,
            I => \N__6636\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6636\,
            I => \U712_CHIP_RAM.N_34\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6633\,
            I => \N__6630\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__6630\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_4\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__6627\,
            I => \N__6624\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6624\,
            I => \N__6621\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6621\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6615\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__6615\,
            I => \N__6612\
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__6612\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6609\,
            I => \N__6606\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6606\,
            I => \N__6603\
        );

    \I__1282\ : Odrv4
    port map (
            O => \N__6603\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6600\,
            I => \N__6597\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__6597\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6590\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6587\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6590\,
            I => \N__6583\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__6587\,
            I => \N__6580\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6577\
        );

    \I__1274\ : Span4Mux_v
    port map (
            O => \N__6583\,
            I => \N__6574\
        );

    \I__1273\ : Span4Mux_h
    port map (
            O => \N__6580\,
            I => \N__6569\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6577\,
            I => \N__6569\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__6574\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__6569\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6564\,
            I => \N__6558\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6555\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6550\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6561\,
            I => \N__6550\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6558\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6555\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__6550\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__6543\,
            I => \N__6540\
        );

    \I__1261\ : InMux
    port map (
            O => \N__6540\,
            I => \N__6536\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6539\,
            I => \N__6533\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6536\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__6533\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6528\,
            I => \N__6525\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__6525\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6519\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6519\,
            I => \N__6516\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__6516\,
            I => \N__6513\
        );

    \I__1252\ : Sp12to4
    port map (
            O => \N__6513\,
            I => \N__6510\
        );

    \I__1251\ : Span12Mux_h
    port map (
            O => \N__6510\,
            I => \N__6507\
        );

    \I__1250\ : Span12Mux_v
    port map (
            O => \N__6507\,
            I => \N__6504\
        );

    \I__1249\ : Odrv12
    port map (
            O => \N__6504\,
            I => \DBRn_c\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__6501\,
            I => \N__6497\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6494\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6497\,
            I => \N__6489\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6494\,
            I => \N__6486\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6493\,
            I => \N__6483\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6480\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6489\,
            I => \N__6477\
        );

    \I__1241\ : Span4Mux_v
    port map (
            O => \N__6486\,
            I => \N__6474\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__6483\,
            I => \N__6471\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__6480\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1238\ : Odrv12
    port map (
            O => \N__6477\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__6474\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__6471\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6462\,
            I => \N__6459\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6459\,
            I => \U712_BYTE_ENABLE.UMBE_0\
        );

    \I__1233\ : IoInMux
    port map (
            O => \N__6456\,
            I => \N__6453\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6453\,
            I => \N__6450\
        );

    \I__1231\ : IoSpan4Mux
    port map (
            O => \N__6450\,
            I => \N__6447\
        );

    \I__1230\ : Span4Mux_s3_v
    port map (
            O => \N__6447\,
            I => \N__6444\
        );

    \I__1229\ : Sp12to4
    port map (
            O => \N__6444\,
            I => \N__6441\
        );

    \I__1228\ : Span12Mux_v
    port map (
            O => \N__6441\,
            I => \N__6438\
        );

    \I__1227\ : Span12Mux_h
    port map (
            O => \N__6438\,
            I => \N__6435\
        );

    \I__1226\ : Odrv12
    port map (
            O => \N__6435\,
            I => \CUMBEn_c\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__6432\,
            I => \N__6429\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6429\,
            I => \N__6426\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6426\,
            I => \N__6423\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__6423\,
            I => \U712_BYTE_ENABLE.UUBE_0\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6420\,
            I => \N__6414\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6419\,
            I => \N__6414\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6414\,
            I => \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_0\
        );

    \I__1218\ : IoInMux
    port map (
            O => \N__6411\,
            I => \N__6408\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__6408\,
            I => \N__6405\
        );

    \I__1216\ : IoSpan4Mux
    port map (
            O => \N__6405\,
            I => \N__6402\
        );

    \I__1215\ : Sp12to4
    port map (
            O => \N__6402\,
            I => \N__6399\
        );

    \I__1214\ : Span12Mux_s7_h
    port map (
            O => \N__6399\,
            I => \N__6396\
        );

    \I__1213\ : Span12Mux_v
    port map (
            O => \N__6396\,
            I => \N__6393\
        );

    \I__1212\ : Odrv12
    port map (
            O => \N__6393\,
            I => \CUUBEn_c\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6387\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6387\,
            I => \N__6384\
        );

    \I__1209\ : Span4Mux_v
    port map (
            O => \N__6384\,
            I => \N__6380\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6383\,
            I => \N__6377\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__6380\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__6377\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__1205\ : IoInMux
    port map (
            O => \N__6372\,
            I => \N__6369\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6369\,
            I => \N__6366\
        );

    \I__1203\ : IoSpan4Mux
    port map (
            O => \N__6366\,
            I => \N__6363\
        );

    \I__1202\ : IoSpan4Mux
    port map (
            O => \N__6363\,
            I => \N__6360\
        );

    \I__1201\ : Span4Mux_s0_v
    port map (
            O => \N__6360\,
            I => \N__6357\
        );

    \I__1200\ : Sp12to4
    port map (
            O => \N__6357\,
            I => \N__6354\
        );

    \I__1199\ : Span12Mux_v
    port map (
            O => \N__6354\,
            I => \N__6351\
        );

    \I__1198\ : Odrv12
    port map (
            O => \N__6351\,
            I => \U712_REG_SM_un1_LDSn_i\
        );

    \I__1197\ : IoInMux
    port map (
            O => \N__6348\,
            I => \N__6345\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6345\,
            I => \N__6342\
        );

    \I__1195\ : Span12Mux_s5_h
    port map (
            O => \N__6342\,
            I => \N__6339\
        );

    \I__1194\ : Span12Mux_h
    port map (
            O => \N__6339\,
            I => \N__6336\
        );

    \I__1193\ : Odrv12
    port map (
            O => \N__6336\,
            I => \CMA_c_3\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6333\,
            I => \N__6330\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__6330\,
            I => \N__6327\
        );

    \I__1190\ : Span4Mux_h
    port map (
            O => \N__6327\,
            I => \N__6324\
        );

    \I__1189\ : Odrv4
    port map (
            O => \N__6324\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__6321\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_START_2_2_cascade_\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6318\,
            I => \N__6313\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6308\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6308\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6313\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6308\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__6303\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_0_sqmuxa_cascade_\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6297\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6297\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_0\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6294\,
            I => \N__6288\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6281\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6292\,
            I => \N__6281\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6281\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6288\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6281\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6276\,
            I => \N__6272\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6275\,
            I => \N__6269\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6272\,
            I => \U712_CHIP_RAM.N_70_2\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6269\,
            I => \U712_CHIP_RAM.N_70_2\
        );

    \I__1169\ : CascadeMux
    port map (
            O => \N__6264\,
            I => \N__6260\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__6263\,
            I => \N__6253\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6250\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6259\,
            I => \N__6247\
        );

    \I__1165\ : InMux
    port map (
            O => \N__6258\,
            I => \N__6244\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__6257\,
            I => \N__6234\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6256\,
            I => \N__6230\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6253\,
            I => \N__6227\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__6250\,
            I => \N__6220\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__6247\,
            I => \N__6220\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6244\,
            I => \N__6220\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6217\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6242\,
            I => \N__6214\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6207\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6240\,
            I => \N__6207\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6207\
        );

    \I__1153\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6204\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6237\,
            I => \N__6197\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6234\,
            I => \N__6197\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6233\,
            I => \N__6197\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6230\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6227\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__6220\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6217\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6214\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6207\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6204\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__6197\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1141\ : CascadeMux
    port map (
            O => \N__6180\,
            I => \N__6175\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6179\,
            I => \N__6170\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6178\,
            I => \N__6170\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6175\,
            I => \N__6167\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6170\,
            I => \U712_CHIP_RAM.N_106\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6167\,
            I => \U712_CHIP_RAM.N_106\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__6162\,
            I => \N__6158\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6152\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6149\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6145\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6156\,
            I => \N__6142\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__6155\,
            I => \N__6139\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6152\,
            I => \N__6136\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6149\,
            I => \N__6133\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__6148\,
            I => \N__6130\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6145\,
            I => \N__6120\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6142\,
            I => \N__6120\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6139\,
            I => \N__6117\
        );

    \I__1123\ : Span4Mux_h
    port map (
            O => \N__6136\,
            I => \N__6112\
        );

    \I__1122\ : Span4Mux_v
    port map (
            O => \N__6133\,
            I => \N__6112\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6130\,
            I => \N__6109\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6129\,
            I => \N__6104\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6128\,
            I => \N__6104\
        );

    \I__1118\ : InMux
    port map (
            O => \N__6127\,
            I => \N__6101\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6126\,
            I => \N__6096\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6096\
        );

    \I__1115\ : Odrv4
    port map (
            O => \N__6120\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6117\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1113\ : Odrv4
    port map (
            O => \N__6112\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6109\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__6104\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6101\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6096\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__6081\,
            I => \N__6078\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6075\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6075\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_3_0\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6072\,
            I => \N__6067\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__6071\,
            I => \N__6064\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6070\,
            I => \N__6061\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6067\,
            I => \N__6058\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6064\,
            I => \N__6055\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6061\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1099\ : Odrv4
    port map (
            O => \N__6058\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__6055\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6048\,
            I => \N__6043\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6047\,
            I => \N__6038\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6046\,
            I => \N__6038\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6043\,
            I => \N__6034\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6038\,
            I => \N__6031\
        );

    \I__1092\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6028\
        );

    \I__1091\ : Span4Mux_h
    port map (
            O => \N__6034\,
            I => \N__6025\
        );

    \I__1090\ : Odrv4
    port map (
            O => \N__6031\,
            I => \U712_CHIP_RAM.N_40\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__6028\,
            I => \U712_CHIP_RAM.N_40\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__6025\,
            I => \U712_CHIP_RAM.N_40\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__6018\,
            I => \U712_CHIP_RAM.N_40_cascade_\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__6015\,
            I => \N__6012\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6012\,
            I => \N__6003\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6011\,
            I => \N__6000\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6010\,
            I => \N__5997\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6009\,
            I => \N__5992\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6008\,
            I => \N__5992\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6007\,
            I => \N__5987\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6006\,
            I => \N__5987\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6003\,
            I => \U712_CHIP_RAM.N_51\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6000\,
            I => \U712_CHIP_RAM.N_51\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5997\,
            I => \U712_CHIP_RAM.N_51\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__5992\,
            I => \U712_CHIP_RAM.N_51\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__5987\,
            I => \U712_CHIP_RAM.N_51\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5976\,
            I => \N__5973\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5973\,
            I => \U712_CHIP_RAM.N_59\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__5970\,
            I => \U712_CHIP_RAM.N_59_cascade_\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5967\,
            I => \N__5962\
        );

    \I__1069\ : InMux
    port map (
            O => \N__5966\,
            I => \N__5958\
        );

    \I__1068\ : InMux
    port map (
            O => \N__5965\,
            I => \N__5955\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5962\,
            I => \N__5949\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5961\,
            I => \N__5946\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5958\,
            I => \N__5941\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__5955\,
            I => \N__5941\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5938\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5933\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5933\
        );

    \I__1060\ : Odrv4
    port map (
            O => \N__5949\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5946\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\
        );

    \I__1058\ : Odrv4
    port map (
            O => \N__5941\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__5938\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__5933\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__5922\,
            I => \N__5919\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5919\,
            I => \N__5906\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5918\,
            I => \N__5906\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__5917\,
            I => \N__5903\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5916\,
            I => \N__5898\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5915\,
            I => \N__5894\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5914\,
            I => \N__5889\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5913\,
            I => \N__5889\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5912\,
            I => \N__5881\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5881\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__5906\,
            I => \N__5878\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5903\,
            I => \N__5875\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5870\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5901\,
            I => \N__5870\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5898\,
            I => \N__5867\
        );

    \I__1040\ : InMux
    port map (
            O => \N__5897\,
            I => \N__5864\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5894\,
            I => \N__5861\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__5889\,
            I => \N__5858\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5854\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5851\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5886\,
            I => \N__5848\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5881\,
            I => \N__5841\
        );

    \I__1033\ : Span4Mux_v
    port map (
            O => \N__5878\,
            I => \N__5841\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5875\,
            I => \N__5841\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__5870\,
            I => \N__5834\
        );

    \I__1030\ : Span4Mux_h
    port map (
            O => \N__5867\,
            I => \N__5834\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5864\,
            I => \N__5834\
        );

    \I__1028\ : Span4Mux_h
    port map (
            O => \N__5861\,
            I => \N__5831\
        );

    \I__1027\ : Span4Mux_h
    port map (
            O => \N__5858\,
            I => \N__5828\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5857\,
            I => \N__5825\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5854\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__5851\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5848\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1022\ : Odrv4
    port map (
            O => \N__5841\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__5834\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1020\ : Odrv4
    port map (
            O => \N__5831\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1019\ : Odrv4
    port map (
            O => \N__5828\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5825\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1017\ : InMux
    port map (
            O => \N__5808\,
            I => \N__5805\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5805\,
            I => \U712_CYCLE_TERM.N_45_0_0_en\
        );

    \I__1015\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5797\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5794\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5791\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5797\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5794\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__5791\,
            I => \U712_CHIP_RAM.N_46\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5781\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5781\,
            I => \U712_CHIP_RAM.N_77\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5778\,
            I => \N__5774\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5771\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__5774\,
            I => \U712_CHIP_RAM.N_99\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__5771\,
            I => \U712_CHIP_RAM.N_99\
        );

    \I__1003\ : CascadeMux
    port map (
            O => \N__5766\,
            I => \U712_CHIP_RAM.N_99_cascade_\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5763\,
            I => \N__5760\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5760\,
            I => \U712_CHIP_RAM.N_79\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5757\,
            I => \N__5751\
        );

    \I__999\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5751\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5751\,
            I => \U712_CHIP_RAM.N_93_1\
        );

    \I__997\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5744\
        );

    \I__996\ : InMux
    port map (
            O => \N__5747\,
            I => \N__5741\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5744\,
            I => \U712_CHIP_RAM.N_52\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5741\,
            I => \U712_CHIP_RAM.N_52\
        );

    \I__993\ : InMux
    port map (
            O => \N__5736\,
            I => \N__5727\
        );

    \I__992\ : InMux
    port map (
            O => \N__5735\,
            I => \N__5724\
        );

    \I__991\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5721\
        );

    \I__990\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5718\
        );

    \I__989\ : InMux
    port map (
            O => \N__5732\,
            I => \N__5713\
        );

    \I__988\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5713\
        );

    \I__987\ : InMux
    port map (
            O => \N__5730\,
            I => \N__5710\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5727\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5724\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5721\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5718\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5713\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5710\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__980\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5694\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__5694\,
            I => \N__5690\
        );

    \I__978\ : InMux
    port map (
            O => \N__5693\,
            I => \N__5687\
        );

    \I__977\ : Odrv4
    port map (
            O => \N__5690\,
            I => \U712_CHIP_RAM.N_54\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5687\,
            I => \U712_CHIP_RAM.N_54\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__5682\,
            I => \N__5674\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__5681\,
            I => \N__5671\
        );

    \I__973\ : InMux
    port map (
            O => \N__5680\,
            I => \N__5667\
        );

    \I__972\ : InMux
    port map (
            O => \N__5679\,
            I => \N__5664\
        );

    \I__971\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5661\
        );

    \I__970\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5656\
        );

    \I__969\ : InMux
    port map (
            O => \N__5674\,
            I => \N__5656\
        );

    \I__968\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5651\
        );

    \I__967\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5651\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5667\,
            I => \N__5648\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__5664\,
            I => \U712_CHIP_RAM.N_50\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5661\,
            I => \U712_CHIP_RAM.N_50\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__5656\,
            I => \U712_CHIP_RAM.N_50\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5651\,
            I => \U712_CHIP_RAM.N_50\
        );

    \I__961\ : Odrv4
    port map (
            O => \N__5648\,
            I => \U712_CHIP_RAM.N_50\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__5637\,
            I => \U712_CHIP_RAM.N_54_cascade_\
        );

    \I__959\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5624\
        );

    \I__958\ : InMux
    port map (
            O => \N__5633\,
            I => \N__5624\
        );

    \I__957\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5621\
        );

    \I__956\ : InMux
    port map (
            O => \N__5631\,
            I => \N__5608\
        );

    \I__955\ : InMux
    port map (
            O => \N__5630\,
            I => \N__5603\
        );

    \I__954\ : InMux
    port map (
            O => \N__5629\,
            I => \N__5603\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5624\,
            I => \N__5598\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__5621\,
            I => \N__5598\
        );

    \I__951\ : InMux
    port map (
            O => \N__5620\,
            I => \N__5595\
        );

    \I__950\ : InMux
    port map (
            O => \N__5619\,
            I => \N__5590\
        );

    \I__949\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5590\
        );

    \I__948\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5583\
        );

    \I__947\ : InMux
    port map (
            O => \N__5616\,
            I => \N__5583\
        );

    \I__946\ : InMux
    port map (
            O => \N__5615\,
            I => \N__5583\
        );

    \I__945\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5574\
        );

    \I__944\ : InMux
    port map (
            O => \N__5613\,
            I => \N__5574\
        );

    \I__943\ : InMux
    port map (
            O => \N__5612\,
            I => \N__5574\
        );

    \I__942\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5574\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5608\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5603\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__939\ : Odrv4
    port map (
            O => \N__5598\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5595\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__5590\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5583\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5574\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__934\ : InMux
    port map (
            O => \N__5559\,
            I => \N__5556\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__5556\,
            I => \N__5553\
        );

    \I__932\ : Span4Mux_v
    port map (
            O => \N__5553\,
            I => \N__5550\
        );

    \I__931\ : Sp12to4
    port map (
            O => \N__5550\,
            I => \N__5547\
        );

    \I__930\ : Span12Mux_h
    port map (
            O => \N__5547\,
            I => \N__5544\
        );

    \I__929\ : Odrv12
    port map (
            O => \N__5544\,
            I => \A_c_11\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__5541\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_\
        );

    \I__927\ : InMux
    port map (
            O => \N__5538\,
            I => \N__5535\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5535\,
            I => \N__5532\
        );

    \I__925\ : Span12Mux_v
    port map (
            O => \N__5532\,
            I => \N__5529\
        );

    \I__924\ : Span12Mux_h
    port map (
            O => \N__5529\,
            I => \N__5526\
        );

    \I__923\ : Odrv12
    port map (
            O => \N__5526\,
            I => \A_c_4\
        );

    \I__922\ : SRMux
    port map (
            O => \N__5523\,
            I => \N__5520\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__5520\,
            I => \N__5517\
        );

    \I__920\ : Span4Mux_h
    port map (
            O => \N__5517\,
            I => \N__5514\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__5514\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__5511\,
            I => \U712_CHIP_RAM.N_78_cascade_\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__5508\,
            I => \U712_CHIP_RAM.N_76_cascade_\
        );

    \I__916\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5499\
        );

    \I__915\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5499\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5499\,
            I => \U712_CHIP_RAM.N_58\
        );

    \I__913\ : InMux
    port map (
            O => \N__5496\,
            I => \N__5490\
        );

    \I__912\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5483\
        );

    \I__911\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5483\
        );

    \I__910\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5483\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5490\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__5483\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\
        );

    \I__907\ : InMux
    port map (
            O => \N__5478\,
            I => \N__5474\
        );

    \I__906\ : InMux
    port map (
            O => \N__5477\,
            I => \N__5471\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5474\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c2\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5471\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c2\
        );

    \I__903\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5463\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5463\,
            I => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__5460\,
            I => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1_cascade_\
        );

    \I__900\ : IoInMux
    port map (
            O => \N__5457\,
            I => \N__5454\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__5454\,
            I => \N__5451\
        );

    \I__898\ : IoSpan4Mux
    port map (
            O => \N__5451\,
            I => \N__5448\
        );

    \I__897\ : Span4Mux_s2_v
    port map (
            O => \N__5448\,
            I => \N__5445\
        );

    \I__896\ : Sp12to4
    port map (
            O => \N__5445\,
            I => \N__5442\
        );

    \I__895\ : Span12Mux_v
    port map (
            O => \N__5442\,
            I => \N__5439\
        );

    \I__894\ : Odrv12
    port map (
            O => \N__5439\,
            I => \CLLBEn_c\
        );

    \I__893\ : IoInMux
    port map (
            O => \N__5436\,
            I => \N__5433\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5433\,
            I => \N__5430\
        );

    \I__891\ : Span4Mux_s1_v
    port map (
            O => \N__5430\,
            I => \N__5427\
        );

    \I__890\ : Sp12to4
    port map (
            O => \N__5427\,
            I => \N__5424\
        );

    \I__889\ : Span12Mux_h
    port map (
            O => \N__5424\,
            I => \N__5419\
        );

    \I__888\ : InMux
    port map (
            O => \N__5423\,
            I => \N__5414\
        );

    \I__887\ : InMux
    port map (
            O => \N__5422\,
            I => \N__5414\
        );

    \I__886\ : Span12Mux_v
    port map (
            O => \N__5419\,
            I => \N__5410\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5414\,
            I => \N__5407\
        );

    \I__884\ : InMux
    port map (
            O => \N__5413\,
            I => \N__5404\
        );

    \I__883\ : Odrv12
    port map (
            O => \N__5410\,
            I => \DBENn_c\
        );

    \I__882\ : Odrv4
    port map (
            O => \N__5407\,
            I => \DBENn_c\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5404\,
            I => \DBENn_c\
        );

    \I__880\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5391\
        );

    \I__879\ : InMux
    port map (
            O => \N__5396\,
            I => \N__5388\
        );

    \I__878\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5385\
        );

    \I__877\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5382\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5391\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5388\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5385\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5382\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__5373\,
            I => \N__5370\
        );

    \I__871\ : InMux
    port map (
            O => \N__5370\,
            I => \N__5367\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5367\,
            I => \N__5362\
        );

    \I__869\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5357\
        );

    \I__868\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5357\
        );

    \I__867\ : Span4Mux_h
    port map (
            O => \N__5362\,
            I => \N__5354\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5357\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__5354\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__864\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5345\
        );

    \I__863\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5342\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5345\,
            I => \U712_REG_SM.N_167_0\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5342\,
            I => \U712_REG_SM.N_167_0\
        );

    \I__860\ : InMux
    port map (
            O => \N__5337\,
            I => \N__5334\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5334\,
            I => \N__5331\
        );

    \I__858\ : Odrv12
    port map (
            O => \N__5331\,
            I => \U712_BYTE_ENABLE.LLBE_0\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__5328\,
            I => \N__5325\
        );

    \I__856\ : InMux
    port map (
            O => \N__5325\,
            I => \N__5322\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__5322\,
            I => \N__5319\
        );

    \I__854\ : Odrv4
    port map (
            O => \N__5319\,
            I => \U712_BYTE_ENABLE.LMBE_0\
        );

    \I__853\ : InMux
    port map (
            O => \N__5316\,
            I => \N__5310\
        );

    \I__852\ : InMux
    port map (
            O => \N__5315\,
            I => \N__5305\
        );

    \I__851\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5305\
        );

    \I__850\ : InMux
    port map (
            O => \N__5313\,
            I => \N__5302\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5310\,
            I => \N__5295\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5305\,
            I => \N__5295\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5302\,
            I => \N__5295\
        );

    \I__846\ : Span4Mux_v
    port map (
            O => \N__5295\,
            I => \N__5292\
        );

    \I__845\ : Span4Mux_v
    port map (
            O => \N__5292\,
            I => \N__5287\
        );

    \I__844\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5282\
        );

    \I__843\ : InMux
    port map (
            O => \N__5290\,
            I => \N__5282\
        );

    \I__842\ : Span4Mux_v
    port map (
            O => \N__5287\,
            I => \N__5279\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5282\,
            I => \N__5276\
        );

    \I__840\ : Sp12to4
    port map (
            O => \N__5279\,
            I => \N__5271\
        );

    \I__839\ : Span12Mux_v
    port map (
            O => \N__5276\,
            I => \N__5271\
        );

    \I__838\ : Odrv12
    port map (
            O => \N__5271\,
            I => \SIZ_c_0\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__5268\,
            I => \N__5265\
        );

    \I__836\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5255\
        );

    \I__835\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5255\
        );

    \I__834\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5255\
        );

    \I__833\ : InMux
    port map (
            O => \N__5262\,
            I => \N__5252\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5255\,
            I => \N__5247\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5252\,
            I => \N__5247\
        );

    \I__830\ : Span4Mux_v
    port map (
            O => \N__5247\,
            I => \N__5244\
        );

    \I__829\ : Span4Mux_v
    port map (
            O => \N__5244\,
            I => \N__5241\
        );

    \I__828\ : Sp12to4
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__827\ : Odrv12
    port map (
            O => \N__5238\,
            I => \A_c_1\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__5235\,
            I => \N__5229\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__5234\,
            I => \N__5226\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__5233\,
            I => \N__5223\
        );

    \I__823\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5214\
        );

    \I__822\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5214\
        );

    \I__821\ : InMux
    port map (
            O => \N__5226\,
            I => \N__5214\
        );

    \I__820\ : InMux
    port map (
            O => \N__5223\,
            I => \N__5211\
        );

    \I__819\ : InMux
    port map (
            O => \N__5222\,
            I => \N__5206\
        );

    \I__818\ : InMux
    port map (
            O => \N__5221\,
            I => \N__5206\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5214\,
            I => \N__5199\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5211\,
            I => \N__5199\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5206\,
            I => \N__5199\
        );

    \I__814\ : Span4Mux_v
    port map (
            O => \N__5199\,
            I => \N__5196\
        );

    \I__813\ : Sp12to4
    port map (
            O => \N__5196\,
            I => \N__5193\
        );

    \I__812\ : Odrv12
    port map (
            O => \N__5193\,
            I => \A_c_0\
        );

    \I__811\ : InMux
    port map (
            O => \N__5190\,
            I => \N__5187\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__5187\,
            I => \N__5184\
        );

    \I__809\ : Span4Mux_v
    port map (
            O => \N__5184\,
            I => \N__5178\
        );

    \I__808\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5173\
        );

    \I__807\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5173\
        );

    \I__806\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5170\
        );

    \I__805\ : Span4Mux_v
    port map (
            O => \N__5178\,
            I => \N__5167\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5173\,
            I => \N__5162\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5170\,
            I => \N__5162\
        );

    \I__802\ : Span4Mux_v
    port map (
            O => \N__5167\,
            I => \N__5159\
        );

    \I__801\ : Sp12to4
    port map (
            O => \N__5162\,
            I => \N__5156\
        );

    \I__800\ : Sp12to4
    port map (
            O => \N__5159\,
            I => \N__5151\
        );

    \I__799\ : Span12Mux_v
    port map (
            O => \N__5156\,
            I => \N__5151\
        );

    \I__798\ : Span12Mux_h
    port map (
            O => \N__5151\,
            I => \N__5148\
        );

    \I__797\ : Odrv12
    port map (
            O => \N__5148\,
            I => \SIZ_c_1\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__5145\,
            I => \N__5141\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__5144\,
            I => \N__5138\
        );

    \I__794\ : InMux
    port map (
            O => \N__5141\,
            I => \N__5134\
        );

    \I__793\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5129\
        );

    \I__792\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5129\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__5134\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5129\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__789\ : InMux
    port map (
            O => \N__5124\,
            I => \N__5121\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5121\,
            I => \U712_CYCLE_TERM.N_49\
        );

    \I__787\ : CascadeMux
    port map (
            O => \N__5118\,
            I => \N__5114\
        );

    \I__786\ : CascadeMux
    port map (
            O => \N__5117\,
            I => \N__5111\
        );

    \I__785\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5107\
        );

    \I__784\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5102\
        );

    \I__783\ : InMux
    port map (
            O => \N__5110\,
            I => \N__5102\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5107\,
            I => \REG_TACK\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5102\,
            I => \REG_TACK\
        );

    \I__780\ : InMux
    port map (
            O => \N__5097\,
            I => \N__5090\
        );

    \I__779\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5090\
        );

    \I__778\ : InMux
    port map (
            O => \N__5095\,
            I => \N__5087\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5090\,
            I => \N__5084\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5087\,
            I => \CPU_TACKm\
        );

    \I__775\ : Odrv4
    port map (
            O => \N__5084\,
            I => \CPU_TACKm\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__5079\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__773\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5073\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5073\,
            I => \N__5068\
        );

    \I__771\ : InMux
    port map (
            O => \N__5072\,
            I => \N__5065\
        );

    \I__770\ : CascadeMux
    port map (
            O => \N__5071\,
            I => \N__5061\
        );

    \I__769\ : Span4Mux_h
    port map (
            O => \N__5068\,
            I => \N__5056\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5065\,
            I => \N__5056\
        );

    \I__767\ : InMux
    port map (
            O => \N__5064\,
            I => \N__5051\
        );

    \I__766\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5051\
        );

    \I__765\ : Span4Mux_h
    port map (
            O => \N__5056\,
            I => \N__5046\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5051\,
            I => \N__5046\
        );

    \I__763\ : Span4Mux_h
    port map (
            O => \N__5046\,
            I => \N__5043\
        );

    \I__762\ : Span4Mux_v
    port map (
            O => \N__5043\,
            I => \N__5040\
        );

    \I__761\ : Span4Mux_v
    port map (
            O => \N__5040\,
            I => \N__5037\
        );

    \I__760\ : Span4Mux_v
    port map (
            O => \N__5037\,
            I => \N__5034\
        );

    \I__759\ : Odrv4
    port map (
            O => \N__5034\,
            I => \CLK40_OUT_i\
        );

    \I__758\ : InMux
    port map (
            O => \N__5031\,
            I => \N__5025\
        );

    \I__757\ : InMux
    port map (
            O => \N__5030\,
            I => \N__5025\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5025\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__755\ : IoInMux
    port map (
            O => \N__5022\,
            I => \N__5019\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5019\,
            I => \N__5016\
        );

    \I__753\ : IoSpan4Mux
    port map (
            O => \N__5016\,
            I => \N__5012\
        );

    \I__752\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5009\
        );

    \I__751\ : Sp12to4
    port map (
            O => \N__5012\,
            I => \N__5005\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__5009\,
            I => \N__5002\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__5008\,
            I => \N__4999\
        );

    \I__748\ : Span12Mux_s9_v
    port map (
            O => \N__5005\,
            I => \N__4996\
        );

    \I__747\ : Span4Mux_v
    port map (
            O => \N__5002\,
            I => \N__4993\
        );

    \I__746\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4990\
        );

    \I__745\ : Odrv12
    port map (
            O => \N__4996\,
            I => \DBDIR_c\
        );

    \I__744\ : Odrv4
    port map (
            O => \N__4993\,
            I => \DBDIR_c\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__4990\,
            I => \DBDIR_c\
        );

    \I__742\ : IoInMux
    port map (
            O => \N__4983\,
            I => \N__4980\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4980\,
            I => \N__4977\
        );

    \I__740\ : Span4Mux_s3_h
    port map (
            O => \N__4977\,
            I => \N__4974\
        );

    \I__739\ : Span4Mux_h
    port map (
            O => \N__4974\,
            I => \N__4971\
        );

    \I__738\ : Sp12to4
    port map (
            O => \N__4971\,
            I => \N__4968\
        );

    \I__737\ : Span12Mux_s6_v
    port map (
            O => \N__4968\,
            I => \N__4965\
        );

    \I__736\ : Span12Mux_h
    port map (
            O => \N__4965\,
            I => \N__4962\
        );

    \I__735\ : Odrv12
    port map (
            O => \N__4962\,
            I => \DRDDIR_0_i\
        );

    \I__734\ : IoInMux
    port map (
            O => \N__4959\,
            I => \N__4956\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4956\,
            I => \N__4953\
        );

    \I__732\ : IoSpan4Mux
    port map (
            O => \N__4953\,
            I => \N__4950\
        );

    \I__731\ : Span4Mux_s0_h
    port map (
            O => \N__4950\,
            I => \N__4947\
        );

    \I__730\ : Sp12to4
    port map (
            O => \N__4947\,
            I => \N__4944\
        );

    \I__729\ : Span12Mux_h
    port map (
            O => \N__4944\,
            I => \N__4941\
        );

    \I__728\ : Span12Mux_v
    port map (
            O => \N__4941\,
            I => \N__4938\
        );

    \I__727\ : Odrv12
    port map (
            O => \N__4938\,
            I => \CLMBEn_c\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__4935\,
            I => \U712_CHIP_RAM.N_106_cascade_\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__4932\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__4929\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_cascade_\
        );

    \I__723\ : IoInMux
    port map (
            O => \N__4926\,
            I => \N__4923\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4923\,
            I => \N__4920\
        );

    \I__721\ : IoSpan4Mux
    port map (
            O => \N__4920\,
            I => \N__4917\
        );

    \I__720\ : Sp12to4
    port map (
            O => \N__4917\,
            I => \N__4914\
        );

    \I__719\ : Span12Mux_s7_h
    port map (
            O => \N__4914\,
            I => \N__4911\
        );

    \I__718\ : Span12Mux_h
    port map (
            O => \N__4911\,
            I => \N__4907\
        );

    \I__717\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4904\
        );

    \I__716\ : Odrv12
    port map (
            O => \N__4907\,
            I => \CLK_EN_c\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4904\,
            I => \CLK_EN_c\
        );

    \I__714\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4895\
        );

    \I__713\ : InMux
    port map (
            O => \N__4898\,
            I => \N__4891\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4895\,
            I => \N__4888\
        );

    \I__711\ : InMux
    port map (
            O => \N__4894\,
            I => \N__4885\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4891\,
            I => \U712_CHIP_RAM.N_100\
        );

    \I__709\ : Odrv4
    port map (
            O => \N__4888\,
            I => \U712_CHIP_RAM.N_100\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4885\,
            I => \U712_CHIP_RAM.N_100\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__4878\,
            I => \N__4875\
        );

    \I__706\ : InMux
    port map (
            O => \N__4875\,
            I => \N__4872\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4872\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0\
        );

    \I__704\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4863\
        );

    \I__703\ : InMux
    port map (
            O => \N__4868\,
            I => \N__4863\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__4863\,
            I => \N__4860\
        );

    \I__701\ : Odrv4
    port map (
            O => \N__4860\,
            I => \U712_CHIP_RAM.CPU_TACK_6\
        );

    \I__700\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4854\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__4854\,
            I => \N__4851\
        );

    \I__698\ : Span12Mux_h
    port map (
            O => \N__4851\,
            I => \N__4848\
        );

    \I__697\ : Span12Mux_v
    port map (
            O => \N__4848\,
            I => \N__4845\
        );

    \I__696\ : Span12Mux_h
    port map (
            O => \N__4845\,
            I => \N__4842\
        );

    \I__695\ : Odrv12
    port map (
            O => \N__4842\,
            I => \RAMSPACEn_c\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__4839\,
            I => \U712_CHIP_RAM.un6_CPU_CYCLE_START_cascade_\
        );

    \I__693\ : InMux
    port map (
            O => \N__4836\,
            I => \N__4833\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4833\,
            I => \N__4829\
        );

    \I__691\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4826\
        );

    \I__690\ : Span4Mux_v
    port map (
            O => \N__4829\,
            I => \N__4823\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4826\,
            I => \N__4820\
        );

    \I__688\ : Span4Mux_h
    port map (
            O => \N__4823\,
            I => \N__4817\
        );

    \I__687\ : Span12Mux_h
    port map (
            O => \N__4820\,
            I => \N__4814\
        );

    \I__686\ : Sp12to4
    port map (
            O => \N__4817\,
            I => \N__4811\
        );

    \I__685\ : Span12Mux_v
    port map (
            O => \N__4814\,
            I => \N__4808\
        );

    \I__684\ : Span12Mux_v
    port map (
            O => \N__4811\,
            I => \N__4805\
        );

    \I__683\ : Odrv12
    port map (
            O => \N__4808\,
            I => \TSn_c\
        );

    \I__682\ : Odrv12
    port map (
            O => \N__4805\,
            I => \TSn_c\
        );

    \I__681\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4796\
        );

    \I__680\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4793\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__4796\,
            I => \N__4790\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__4793\,
            I => \U712_CHIP_RAM.N_68\
        );

    \I__677\ : Odrv4
    port map (
            O => \N__4790\,
            I => \U712_CHIP_RAM.N_68\
        );

    \I__676\ : InMux
    port map (
            O => \N__4785\,
            I => \N__4781\
        );

    \I__675\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4778\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__4781\,
            I => \U712_CHIP_RAM.N_98\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4778\,
            I => \U712_CHIP_RAM.N_98\
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__4773\,
            I => \U712_CHIP_RAM.N_55_cascade_\
        );

    \I__671\ : CascadeMux
    port map (
            O => \N__4770\,
            I => \U712_CHIP_RAM.N_57_cascade_\
        );

    \I__670\ : CascadeMux
    port map (
            O => \N__4767\,
            I => \U712_CHIP_RAM.N_92_cascade_\
        );

    \I__669\ : InMux
    port map (
            O => \N__4764\,
            I => \N__4760\
        );

    \I__668\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4757\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4760\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__4757\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__665\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4745\
        );

    \I__664\ : InMux
    port map (
            O => \N__4751\,
            I => \N__4736\
        );

    \I__663\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4736\
        );

    \I__662\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4736\
        );

    \I__661\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4736\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4745\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4736\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__658\ : InMux
    port map (
            O => \N__4731\,
            I => \N__4725\
        );

    \I__657\ : InMux
    port map (
            O => \N__4730\,
            I => \N__4725\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__4725\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_3\
        );

    \I__655\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4719\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4719\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER17_1\
        );

    \I__653\ : CascadeMux
    port map (
            O => \N__4716\,
            I => \U712_CHIP_RAM.N_50_cascade_\
        );

    \I__652\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4708\
        );

    \I__651\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4705\
        );

    \I__650\ : InMux
    port map (
            O => \N__4711\,
            I => \N__4702\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4708\,
            I => \U712_CHIP_RAM.N_43\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4705\,
            I => \U712_CHIP_RAM.N_43\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4702\,
            I => \U712_CHIP_RAM.N_43\
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__4695\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_tz_1_cascade_\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__4692\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_\
        );

    \I__644\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4686\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4686\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__4683\,
            I => \U712_REG_SM.N_165_0_cascade_\
        );

    \I__641\ : InMux
    port map (
            O => \N__4680\,
            I => \N__4677\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4677\,
            I => \U712_REG_SM.N_170_0\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__4674\,
            I => \N__4667\
        );

    \I__638\ : InMux
    port map (
            O => \N__4673\,
            I => \N__4664\
        );

    \I__637\ : InMux
    port map (
            O => \N__4672\,
            I => \N__4661\
        );

    \I__636\ : InMux
    port map (
            O => \N__4671\,
            I => \N__4656\
        );

    \I__635\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4656\
        );

    \I__634\ : InMux
    port map (
            O => \N__4667\,
            I => \N__4653\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4664\,
            I => \N__4650\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__4661\,
            I => \N__4647\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4656\,
            I => \U712_REG_SM.N_173_0\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4653\,
            I => \U712_REG_SM.N_173_0\
        );

    \I__629\ : Odrv4
    port map (
            O => \N__4650\,
            I => \U712_REG_SM.N_173_0\
        );

    \I__628\ : Odrv4
    port map (
            O => \N__4647\,
            I => \U712_REG_SM.N_173_0\
        );

    \I__627\ : InMux
    port map (
            O => \N__4638\,
            I => \N__4635\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__4635\,
            I => \U712_REG_SM.LDS_OUT_2_0_0\
        );

    \I__625\ : InMux
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__4629\,
            I => \U712_REG_SM.UDS_OUT_2_0_0\
        );

    \I__623\ : CascadeMux
    port map (
            O => \N__4626\,
            I => \U712_CHIP_RAM.N_105_cascade_\
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__4623\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_1_1_cascade_\
        );

    \I__621\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4617\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__4617\,
            I => \U712_CHIP_RAM.N_105\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__4614\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_1_cascade_\
        );

    \I__618\ : CascadeMux
    port map (
            O => \N__4611\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_cascade_\
        );

    \I__617\ : IoInMux
    port map (
            O => \N__4608\,
            I => \N__4605\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4605\,
            I => \N__4602\
        );

    \I__615\ : Span4Mux_s2_h
    port map (
            O => \N__4602\,
            I => \N__4599\
        );

    \I__614\ : Sp12to4
    port map (
            O => \N__4599\,
            I => \N__4596\
        );

    \I__613\ : Span12Mux_v
    port map (
            O => \N__4596\,
            I => \N__4592\
        );

    \I__612\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4589\
        );

    \I__611\ : Odrv12
    port map (
            O => \N__4592\,
            I => \TACK_OUTn\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4589\,
            I => \TACK_OUTn\
        );

    \I__609\ : InMux
    port map (
            O => \N__4584\,
            I => \N__4581\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4581\,
            I => \N__4578\
        );

    \I__607\ : Odrv4
    port map (
            O => \N__4578\,
            I => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__4575\,
            I => \N__4572\
        );

    \I__605\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4569\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4569\,
            I => \U712_REG_SM.DS_EN_7_0\
        );

    \I__603\ : InMux
    port map (
            O => \N__4566\,
            I => \N__4563\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4563\,
            I => \U712_REG_SM.N_187\
        );

    \I__601\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4556\
        );

    \I__600\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4553\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4556\,
            I => \U712_REG_SM.N_157_0\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__4553\,
            I => \U712_REG_SM.N_157_0\
        );

    \I__597\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4541\
        );

    \I__596\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4532\
        );

    \I__595\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4532\
        );

    \I__594\ : InMux
    port map (
            O => \N__4545\,
            I => \N__4532\
        );

    \I__593\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4532\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4541\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4532\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__590\ : InMux
    port map (
            O => \N__4527\,
            I => \N__4524\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4524\,
            I => \N__4519\
        );

    \I__588\ : InMux
    port map (
            O => \N__4523\,
            I => \N__4516\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__4522\,
            I => \N__4513\
        );

    \I__586\ : Span4Mux_v
    port map (
            O => \N__4519\,
            I => \N__4505\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__4516\,
            I => \N__4505\
        );

    \I__584\ : InMux
    port map (
            O => \N__4513\,
            I => \N__4496\
        );

    \I__583\ : InMux
    port map (
            O => \N__4512\,
            I => \N__4496\
        );

    \I__582\ : InMux
    port map (
            O => \N__4511\,
            I => \N__4496\
        );

    \I__581\ : InMux
    port map (
            O => \N__4510\,
            I => \N__4496\
        );

    \I__580\ : Odrv4
    port map (
            O => \N__4505\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__4496\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__578\ : InMux
    port map (
            O => \N__4491\,
            I => \N__4486\
        );

    \I__577\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4483\
        );

    \I__576\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4480\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4486\,
            I => \U712_REG_SM.N_159_0\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4483\,
            I => \U712_REG_SM.N_159_0\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4480\,
            I => \U712_REG_SM.N_159_0\
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__4473\,
            I => \U712_REG_SM.N_159_0_cascade_\
        );

    \I__571\ : InMux
    port map (
            O => \N__4470\,
            I => \N__4465\
        );

    \I__570\ : InMux
    port map (
            O => \N__4469\,
            I => \N__4462\
        );

    \I__569\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4459\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4465\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4462\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4459\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__565\ : InMux
    port map (
            O => \N__4452\,
            I => \N__4449\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4449\,
            I => \U712_REG_SM.N_165_0\
        );

    \I__563\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4437\
        );

    \I__562\ : InMux
    port map (
            O => \N__4445\,
            I => \N__4437\
        );

    \I__561\ : InMux
    port map (
            O => \N__4444\,
            I => \N__4430\
        );

    \I__560\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4430\
        );

    \I__559\ : InMux
    port map (
            O => \N__4442\,
            I => \N__4430\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__4437\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__4430\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__556\ : CascadeMux
    port map (
            O => \N__4425\,
            I => \N__4421\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__4424\,
            I => \N__4417\
        );

    \I__554\ : InMux
    port map (
            O => \N__4421\,
            I => \N__4410\
        );

    \I__553\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4410\
        );

    \I__552\ : InMux
    port map (
            O => \N__4417\,
            I => \N__4403\
        );

    \I__551\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4403\
        );

    \I__550\ : InMux
    port map (
            O => \N__4415\,
            I => \N__4403\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4410\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4403\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__547\ : CascadeMux
    port map (
            O => \N__4398\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_1_cascade_\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__4395\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_2_cascade_\
        );

    \I__545\ : CascadeMux
    port map (
            O => \N__4392\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_0_cascade_\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__4389\,
            I => \N__4383\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__4388\,
            I => \N__4380\
        );

    \I__542\ : InMux
    port map (
            O => \N__4387\,
            I => \N__4377\
        );

    \I__541\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4372\
        );

    \I__540\ : InMux
    port map (
            O => \N__4383\,
            I => \N__4372\
        );

    \I__539\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4369\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4377\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__4372\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4369\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__4362\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_a2_0_4_cascade_\
        );

    \I__534\ : InMux
    port map (
            O => \N__4359\,
            I => \N__4356\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__4356\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_a2_0_1\
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__4353\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__4350\,
            I => \U712_CHIP_RAM.N_43_cascade_\
        );

    \I__530\ : InMux
    port map (
            O => \N__4347\,
            I => \N__4344\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__4344\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6\
        );

    \I__528\ : InMux
    port map (
            O => \N__4341\,
            I => \N__4332\
        );

    \I__527\ : InMux
    port map (
            O => \N__4340\,
            I => \N__4332\
        );

    \I__526\ : InMux
    port map (
            O => \N__4339\,
            I => \N__4332\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__4332\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4\
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__4329\,
            I => \U712_REG_SM.N_162_0_cascade_\
        );

    \I__523\ : InMux
    port map (
            O => \N__4326\,
            I => \N__4320\
        );

    \I__522\ : InMux
    port map (
            O => \N__4325\,
            I => \N__4320\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4320\,
            I => \U712_REG_SM.N_172_0\
        );

    \I__520\ : CascadeMux
    port map (
            O => \N__4317\,
            I => \N__4311\
        );

    \I__519\ : InMux
    port map (
            O => \N__4316\,
            I => \N__4308\
        );

    \I__518\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4303\
        );

    \I__517\ : InMux
    port map (
            O => \N__4314\,
            I => \N__4303\
        );

    \I__516\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4300\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4308\,
            I => \U712_REG_SM.N_162_0\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__4303\,
            I => \U712_REG_SM.N_162_0\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4300\,
            I => \U712_REG_SM.N_162_0\
        );

    \I__512\ : InMux
    port map (
            O => \N__4293\,
            I => \N__4289\
        );

    \I__511\ : InMux
    port map (
            O => \N__4292\,
            I => \N__4286\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__4289\,
            I => \U712_REG_SM.N_195\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4286\,
            I => \U712_REG_SM.N_195\
        );

    \I__508\ : CascadeMux
    port map (
            O => \N__4281\,
            I => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_\
        );

    \I__507\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4274\
        );

    \I__506\ : InMux
    port map (
            O => \N__4277\,
            I => \N__4271\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4274\,
            I => \N__4264\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__4271\,
            I => \N__4264\
        );

    \I__503\ : InMux
    port map (
            O => \N__4270\,
            I => \N__4259\
        );

    \I__502\ : InMux
    port map (
            O => \N__4269\,
            I => \N__4259\
        );

    \I__501\ : Odrv4
    port map (
            O => \N__4264\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4259\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__4254\,
            I => \N__4251\
        );

    \I__498\ : InMux
    port map (
            O => \N__4251\,
            I => \N__4245\
        );

    \I__497\ : InMux
    port map (
            O => \N__4250\,
            I => \N__4245\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4245\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__495\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4235\
        );

    \I__494\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4232\
        );

    \I__493\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4227\
        );

    \I__492\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4227\
        );

    \I__491\ : InMux
    port map (
            O => \N__4238\,
            I => \N__4224\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4235\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4232\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4227\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4224\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__486\ : CascadeMux
    port map (
            O => \N__4215\,
            I => \N__4211\
        );

    \I__485\ : InMux
    port map (
            O => \N__4214\,
            I => \N__4206\
        );

    \I__484\ : InMux
    port map (
            O => \N__4211\,
            I => \N__4203\
        );

    \I__483\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4200\
        );

    \I__482\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4197\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4206\,
            I => \N__4192\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4203\,
            I => \N__4192\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4200\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__4197\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__477\ : Odrv4
    port map (
            O => \N__4192\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__476\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4178\
        );

    \I__475\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4178\
        );

    \I__474\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4175\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__4178\,
            I => \U712_REG_SM.N_163_0\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4175\,
            I => \U712_REG_SM.N_163_0\
        );

    \I__471\ : InMux
    port map (
            O => \N__4170\,
            I => \N__4166\
        );

    \I__470\ : InMux
    port map (
            O => \N__4169\,
            I => \N__4163\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4166\,
            I => \N__4160\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4163\,
            I => \U712_REG_SM.N_194\
        );

    \I__467\ : Odrv4
    port map (
            O => \N__4160\,
            I => \U712_REG_SM.N_194\
        );

    \I__466\ : InMux
    port map (
            O => \N__4155\,
            I => \N__4152\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4152\,
            I => \N__4147\
        );

    \I__464\ : InMux
    port map (
            O => \N__4151\,
            I => \N__4142\
        );

    \I__463\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4142\
        );

    \I__462\ : Odrv4
    port map (
            O => \N__4147\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4142\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__460\ : IoInMux
    port map (
            O => \N__4137\,
            I => \N__4134\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4134\,
            I => \N__4130\
        );

    \I__458\ : IoInMux
    port map (
            O => \N__4133\,
            I => \N__4127\
        );

    \I__457\ : IoSpan4Mux
    port map (
            O => \N__4130\,
            I => \N__4124\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4127\,
            I => \N__4121\
        );

    \I__455\ : Sp12to4
    port map (
            O => \N__4124\,
            I => \N__4118\
        );

    \I__454\ : IoSpan4Mux
    port map (
            O => \N__4121\,
            I => \N__4115\
        );

    \I__453\ : Span12Mux_v
    port map (
            O => \N__4118\,
            I => \N__4112\
        );

    \I__452\ : Sp12to4
    port map (
            O => \N__4115\,
            I => \N__4109\
        );

    \I__451\ : Span12Mux_h
    port map (
            O => \N__4112\,
            I => \N__4104\
        );

    \I__450\ : Span12Mux_v
    port map (
            O => \N__4109\,
            I => \N__4104\
        );

    \I__449\ : Odrv12
    port map (
            O => \N__4104\,
            I => \ASn_c\
        );

    \I__448\ : CEMux
    port map (
            O => \N__4101\,
            I => \N__4098\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__4098\,
            I => \N__4095\
        );

    \I__446\ : Span4Mux_v
    port map (
            O => \N__4095\,
            I => \N__4092\
        );

    \I__445\ : Odrv4
    port map (
            O => \N__4092\,
            I => \U712_REG_SM.N_186_0\
        );

    \I__444\ : IoInMux
    port map (
            O => \N__4089\,
            I => \N__4086\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4086\,
            I => \N__4083\
        );

    \I__442\ : Span12Mux_s10_h
    port map (
            O => \N__4083\,
            I => \N__4080\
        );

    \I__441\ : Odrv12
    port map (
            O => \N__4080\,
            I => \N_510_i\
        );

    \I__440\ : IoInMux
    port map (
            O => \N__4077\,
            I => \N__4074\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4074\,
            I => \N__4071\
        );

    \I__438\ : Span12Mux_s8_v
    port map (
            O => \N__4071\,
            I => \N__4068\
        );

    \I__437\ : Odrv12
    port map (
            O => \N__4068\,
            I => \VBENn_c\
        );

    \I__436\ : CascadeMux
    port map (
            O => \N__4065\,
            I => \U712_REG_SM.N_175_cascade_\
        );

    \I__435\ : InMux
    port map (
            O => \N__4062\,
            I => \N__4059\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__4059\,
            I => \N__4056\
        );

    \I__433\ : Odrv4
    port map (
            O => \N__4056\,
            I => \U712_REG_SM.N_171_0\
        );

    \I__432\ : CascadeMux
    port map (
            O => \N__4053\,
            I => \U712_REG_SM.N_194_cascade_\
        );

    \I__431\ : CascadeMux
    port map (
            O => \N__4050\,
            I => \N__4045\
        );

    \I__430\ : InMux
    port map (
            O => \N__4049\,
            I => \N__4038\
        );

    \I__429\ : InMux
    port map (
            O => \N__4048\,
            I => \N__4038\
        );

    \I__428\ : InMux
    port map (
            O => \N__4045\,
            I => \N__4038\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__4038\,
            I => \U712_REG_SM.N_169_0\
        );

    \I__426\ : InMux
    port map (
            O => \N__4035\,
            I => \N__4029\
        );

    \I__425\ : InMux
    port map (
            O => \N__4034\,
            I => \N__4029\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__4029\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__423\ : CascadeMux
    port map (
            O => \N__4026\,
            I => \U712_REG_SM.N_170_0_cascade_\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__4023\,
            I => \U712_REG_SM.N_174_cascade_\
        );

    \I__421\ : InMux
    port map (
            O => \N__4020\,
            I => \N__4016\
        );

    \I__420\ : InMux
    port map (
            O => \N__4019\,
            I => \N__4013\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__4016\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__4013\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__417\ : InMux
    port map (
            O => \N__4008\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__416\ : InMux
    port map (
            O => \N__4005\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__415\ : InMux
    port map (
            O => \N__4002\,
            I => \N__3998\
        );

    \I__414\ : InMux
    port map (
            O => \N__4001\,
            I => \N__3995\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__3998\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__3995\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__411\ : ClkMux
    port map (
            O => \N__3990\,
            I => \N__3987\
        );

    \I__410\ : GlobalMux
    port map (
            O => \N__3987\,
            I => \N__3984\
        );

    \I__409\ : gio2CtrlBuf
    port map (
            O => \N__3984\,
            I => \C1_c_g\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__3981\,
            I => \N__3977\
        );

    \I__407\ : InMux
    port map (
            O => \N__3980\,
            I => \N__3973\
        );

    \I__406\ : InMux
    port map (
            O => \N__3977\,
            I => \N__3970\
        );

    \I__405\ : InMux
    port map (
            O => \N__3976\,
            I => \N__3967\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__3973\,
            I => \N__3964\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__3970\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3967\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__401\ : Odrv4
    port map (
            O => \N__3964\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__400\ : CascadeMux
    port map (
            O => \N__3957\,
            I => \N__3953\
        );

    \I__399\ : InMux
    port map (
            O => \N__3956\,
            I => \N__3949\
        );

    \I__398\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3945\
        );

    \I__397\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3942\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3949\,
            I => \N__3939\
        );

    \I__395\ : InMux
    port map (
            O => \N__3948\,
            I => \N__3936\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3945\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3942\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__392\ : Odrv4
    port map (
            O => \N__3939\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__3936\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__390\ : CascadeMux
    port map (
            O => \N__3927\,
            I => \U712_REG_SM.N_168_0_cascade_\
        );

    \I__389\ : CascadeMux
    port map (
            O => \N__3924\,
            I => \N__3920\
        );

    \I__388\ : CascadeMux
    port map (
            O => \N__3923\,
            I => \N__3917\
        );

    \I__387\ : InMux
    port map (
            O => \N__3920\,
            I => \N__3909\
        );

    \I__386\ : InMux
    port map (
            O => \N__3917\,
            I => \N__3909\
        );

    \I__385\ : InMux
    port map (
            O => \N__3916\,
            I => \N__3909\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__3909\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__383\ : InMux
    port map (
            O => \N__3906\,
            I => \N__3903\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3903\,
            I => \N__3900\
        );

    \I__381\ : Span4Mux_v
    port map (
            O => \N__3900\,
            I => \N__3897\
        );

    \I__380\ : Sp12to4
    port map (
            O => \N__3897\,
            I => \N__3894\
        );

    \I__379\ : Span12Mux_h
    port map (
            O => \N__3894\,
            I => \N__3891\
        );

    \I__378\ : Odrv12
    port map (
            O => \N__3891\,
            I => \C3_c\
        );

    \I__377\ : CascadeMux
    port map (
            O => \N__3888\,
            I => \U712_CHIP_RAM.REFRESH_r_1_cascade_\
        );

    \I__376\ : InMux
    port map (
            O => \N__3885\,
            I => \N__3882\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__3882\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__374\ : InMux
    port map (
            O => \N__3879\,
            I => \bfn_7_7_0_\
        );

    \I__373\ : InMux
    port map (
            O => \N__3876\,
            I => \N__3873\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3873\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__371\ : InMux
    port map (
            O => \N__3870\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__370\ : InMux
    port map (
            O => \N__3867\,
            I => \N__3863\
        );

    \I__369\ : InMux
    port map (
            O => \N__3866\,
            I => \N__3860\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3863\,
            I => \U712_CHIP_RAM.REFRESH6lto2\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__3860\,
            I => \U712_CHIP_RAM.REFRESH6lto2\
        );

    \I__366\ : InMux
    port map (
            O => \N__3855\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__365\ : InMux
    port map (
            O => \N__3852\,
            I => \N__3848\
        );

    \I__364\ : InMux
    port map (
            O => \N__3851\,
            I => \N__3845\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3848\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__3845\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__361\ : InMux
    port map (
            O => \N__3840\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__360\ : InMux
    port map (
            O => \N__3837\,
            I => \N__3833\
        );

    \I__359\ : InMux
    port map (
            O => \N__3836\,
            I => \N__3830\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3833\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__3830\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__356\ : InMux
    port map (
            O => \N__3825\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__355\ : CascadeMux
    port map (
            O => \N__3822\,
            I => \N__3818\
        );

    \I__354\ : InMux
    port map (
            O => \N__3821\,
            I => \N__3815\
        );

    \I__353\ : InMux
    port map (
            O => \N__3818\,
            I => \N__3812\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__3815\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3812\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__350\ : InMux
    port map (
            O => \N__3807\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__349\ : IoInMux
    port map (
            O => \N__3804\,
            I => \N__3801\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3801\,
            I => \N__3798\
        );

    \I__347\ : Span4Mux_s2_v
    port map (
            O => \N__3798\,
            I => \N__3795\
        );

    \I__346\ : Span4Mux_v
    port map (
            O => \N__3795\,
            I => \N__3792\
        );

    \I__345\ : Odrv4
    port map (
            O => \N__3792\,
            I => \CLK80_OUT_i_i\
        );

    \I__344\ : IoInMux
    port map (
            O => \N__3789\,
            I => \N__3786\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3786\,
            I => \N__3783\
        );

    \I__342\ : Odrv12
    port map (
            O => \N__3783\,
            I => \CLK40_OUT_i_i\
        );

    \I__341\ : InMux
    port map (
            O => \N__3780\,
            I => \N__3777\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__3777\,
            I => \N__3774\
        );

    \I__339\ : Span4Mux_v
    port map (
            O => \N__3774\,
            I => \N__3771\
        );

    \I__338\ : Span4Mux_h
    port map (
            O => \N__3771\,
            I => \N__3768\
        );

    \I__337\ : Sp12to4
    port map (
            O => \N__3768\,
            I => \N__3765\
        );

    \I__336\ : Span12Mux_v
    port map (
            O => \N__3765\,
            I => \N__3762\
        );

    \I__335\ : Odrv12
    port map (
            O => \N__3762\,
            I => \REGSPACEn_c\
        );

    \I__334\ : CascadeMux
    port map (
            O => \N__3759\,
            I => \U712_REG_SM.un6_REG_CYCLE_START_cascade_\
        );

    \I__333\ : InMux
    port map (
            O => \N__3756\,
            I => \N__3752\
        );

    \I__332\ : InMux
    port map (
            O => \N__3755\,
            I => \N__3749\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__3752\,
            I => \U712_REG_SM.REG_CYCLE_GOZ0\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__3749\,
            I => \U712_REG_SM.REG_CYCLE_GOZ0\
        );

    \I__329\ : InMux
    port map (
            O => \N__3744\,
            I => \N__3741\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__3741\,
            I => \N__3737\
        );

    \I__327\ : IoInMux
    port map (
            O => \N__3740\,
            I => \N__3734\
        );

    \I__326\ : Span4Mux_v
    port map (
            O => \N__3737\,
            I => \N__3731\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__3734\,
            I => \N__3728\
        );

    \I__324\ : Sp12to4
    port map (
            O => \N__3731\,
            I => \N__3725\
        );

    \I__323\ : Span4Mux_s3_h
    port map (
            O => \N__3728\,
            I => \N__3722\
        );

    \I__322\ : Span12Mux_h
    port map (
            O => \N__3725\,
            I => \N__3717\
        );

    \I__321\ : Sp12to4
    port map (
            O => \N__3722\,
            I => \N__3717\
        );

    \I__320\ : Span12Mux_v
    port map (
            O => \N__3717\,
            I => \N__3714\
        );

    \I__319\ : Odrv12
    port map (
            O => \N__3714\,
            I => \C1_c\
        );

    \I__318\ : IoInMux
    port map (
            O => \N__3711\,
            I => \N__3708\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__3708\,
            I => \N__3705\
        );

    \I__316\ : IoSpan4Mux
    port map (
            O => \N__3705\,
            I => \N__3702\
        );

    \I__315\ : Span4Mux_s2_v
    port map (
            O => \N__3702\,
            I => \N__3699\
        );

    \I__314\ : Sp12to4
    port map (
            O => \N__3699\,
            I => \N__3696\
        );

    \I__313\ : Span12Mux_v
    port map (
            O => \N__3696\,
            I => \N__3693\
        );

    \I__312\ : Odrv12
    port map (
            O => \N__3693\,
            I => \CLK40_IN_c\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7812\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3740\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9537\,
            lcout => \CLK80_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40C_obuf_RNO_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5076\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3755\,
            in2 => \_gnd_net_\,
            in3 => \N__3952\,
            lcout => OPEN,
            ltout => \U712_REG_SM.un6_REG_CYCLE_START_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__7996\,
            in1 => \N__3780\,
            in2 => \N__3759\,
            in3 => \N__4836\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9524\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_GO_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011101100"
        )
    port map (
            in0 => \N__3976\,
            in1 => \N__3756\,
            in2 => \N__3957\,
            in3 => \N__4673\,
            lcout => \U712_REG_SM.REG_CYCLE_GOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9527\,
            ce => 'H',
            sr => \N__9293\
        );

    \U712_REG_SM.C3_SYNC_1_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4278\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9530\,
            ce => 'H',
            sr => \N__9284\
        );

    \U712_REG_SM.C1_SYNC_0_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3744\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9530\,
            ce => 'H',
            sr => \N__9284\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__3956\,
            in1 => \N__4316\,
            in2 => \N__3981\,
            in3 => \N__4293\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9530\,
            ce => 'H',
            sr => \N__9284\
        );

    \U712_REG_SM.C1_SYNC_2_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4210\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9531\,
            ce => 'H',
            sr => \N__9277\
        );

    \U712_REG_SM.C1_SYNC_1_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4242\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9531\,
            ce => 'H',
            sr => \N__9277\
        );

    \U712_REG_SM.C3_SYNC_0_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3906\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9533\,
            ce => 'H',
            sr => \N__9270\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__3836\,
            in1 => \N__3851\,
            in2 => \N__3822\,
            in3 => \N__3866\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH_r_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__8007\,
            in1 => \N__4001\,
            in2 => \N__3888\,
            in3 => \N__4019\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9510\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3885\,
            in2 => \_gnd_net_\,
            in3 => \N__3879\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__3990\,
            ce => 'H',
            sr => \N__5523\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3876\,
            in2 => \_gnd_net_\,
            in3 => \N__3870\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__3990\,
            ce => 'H',
            sr => \N__5523\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3867\,
            in2 => \_gnd_net_\,
            in3 => \N__3855\,
            lcout => \U712_CHIP_RAM.REFRESH6lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__3990\,
            ce => 'H',
            sr => \N__5523\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3852\,
            in2 => \_gnd_net_\,
            in3 => \N__3840\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__3990\,
            ce => 'H',
            sr => \N__5523\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3837\,
            in2 => \_gnd_net_\,
            in3 => \N__3825\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__3990\,
            ce => 'H',
            sr => \N__5523\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3821\,
            in2 => \_gnd_net_\,
            in3 => \N__3807\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__3990\,
            ce => 'H',
            sr => \N__5523\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4020\,
            in2 => \_gnd_net_\,
            in3 => \N__4008\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__3990\,
            ce => 'H',
            sr => \N__5523\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4002\,
            in2 => \_gnd_net_\,
            in3 => \N__4005\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3990\,
            ce => 'H',
            sr => \N__5523\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3980\,
            in2 => \_gnd_net_\,
            in3 => \N__3948\,
            lcout => \U712_REG_SM.N_171_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__6971\,
            in1 => \N__4277\,
            in2 => \_gnd_net_\,
            in3 => \N__4241\,
            lcout => \U712_REG_SM.DS_EN_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__4672\,
            in1 => \N__7898\,
            in2 => \N__3924\,
            in3 => \N__4049\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_4_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5366\,
            in1 => \N__6593\,
            in2 => \N__6501\,
            in3 => \N__4490\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_168_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__4470\,
            in1 => \N__7900\,
            in2 => \N__3927\,
            in3 => \N__4452\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4050\,
            in3 => \N__3916\,
            lcout => \U712_REG_SM.N_187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5365\,
            in2 => \N__3923\,
            in3 => \N__4048\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_175_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__7899\,
            in1 => \_gnd_net_\,
            in2 => \N__4065\,
            in3 => \N__5349\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9525\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__8002\,
            in1 => \N__4062\,
            in2 => \N__4674\,
            in3 => \N__4035\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9528\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNICU4F1_1_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4510\,
            in1 => \N__4544\,
            in2 => \N__4215\,
            in3 => \N__4238\,
            lcout => \U712_REG_SM.N_194\,
            ltout => \U712_REG_SM.N_194_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4053\,
            in3 => \N__4150\,
            lcout => \U712_REG_SM.N_195\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__4512\,
            in1 => \N__4560\,
            in2 => \_gnd_net_\,
            in3 => \N__4546\,
            lcout => \U712_REG_SM.N_169_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4545\,
            in1 => \N__4034\,
            in2 => \_gnd_net_\,
            in3 => \N__4511\,
            lcout => \U712_REG_SM.N_172_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__4314\,
            in1 => \N__4183\,
            in2 => \N__4522\,
            in3 => \N__4547\,
            lcout => \U712_REG_SM.N_170_0\,
            ltout => \U712_REG_SM.N_170_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5394\,
            in2 => \N__4026\,
            in3 => \N__4151\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_174_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__4315\,
            in1 => \N__8003\,
            in2 => \N__4023\,
            in3 => \N__4169\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9528\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4270\,
            in2 => \_gnd_net_\,
            in3 => \N__4250\,
            lcout => \U712_REG_SM.N_162_0\,
            ltout => \U712_REG_SM.N_162_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__4185\,
            in1 => \_gnd_net_\,
            in2 => \N__4329\,
            in3 => \N__4326\,
            lcout => \U712_REG_SM.N_173_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__4184\,
            in1 => \N__4325\,
            in2 => \N__4317\,
            in3 => \N__4292\,
            lcout => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1\,
            ltout => \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_1_ess_RNO_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4281\,
            in3 => \N__9355\,
            lcout => \U712_REG_SM.N_186_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4269\,
            in1 => \N__4209\,
            in2 => \N__4254\,
            in3 => \N__4239\,
            lcout => \U712_REG_SM.N_157_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4240\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4214\,
            lcout => \U712_REG_SM.N_163_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_1_ess_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4170\,
            in2 => \_gnd_net_\,
            in3 => \N__4155\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9532\,
            ce => \N__4101\,
            sr => \N__9265\
        );

    \TACKn_obuft_RNO_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6801\,
            lcout => \N_510_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7185\,
            in2 => \_gnd_net_\,
            in3 => \N__8298\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6242\,
            in1 => \N__5916\,
            in2 => \N__6162\,
            in3 => \N__5632\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__4751\,
            in1 => \N__9364\,
            in2 => \N__4424\,
            in3 => \N__4341\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_4_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4339\,
            in1 => \N__4416\,
            in2 => \_gnd_net_\,
            in3 => \N__4749\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9365\,
            in2 => \N__4353\,
            in3 => \N__4443\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4442\,
            in1 => \N__4415\,
            in2 => \N__4388\,
            in3 => \N__4748\,
            lcout => \U712_CHIP_RAM.N_43\,
            ltout => \U712_CHIP_RAM.N_43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4350\,
            in3 => \N__5915\,
            lcout => \U712_CHIP_RAM.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__4444\,
            in1 => \N__4347\,
            in2 => \N__9369\,
            in3 => \N__4387\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__4750\,
            in1 => \N__9363\,
            in2 => \_gnd_net_\,
            in3 => \N__4340\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9503\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4898\,
            in1 => \N__6161\,
            in2 => \N__6263\,
            in3 => \N__5735\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5616\,
            in1 => \N__5913\,
            in2 => \_gnd_net_\,
            in3 => \N__4712\,
            lcout => \U712_CHIP_RAM.N_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3EPC1_5_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4445\,
            in1 => \N__4420\,
            in2 => \_gnd_net_\,
            in3 => \N__5615\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__4386\,
            in1 => \N__4446\,
            in2 => \N__4425\,
            in3 => \N__4731\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__6009\,
            in1 => \_gnd_net_\,
            in2 => \N__4398\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000100000"
        )
    port map (
            in0 => \N__5617\,
            in1 => \N__5914\,
            in2 => \N__4395\,
            in3 => \N__6256\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__4869\,
            in1 => \N__7995\,
            in2 => \N__4392\,
            in3 => \N__5095\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9511\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6F3C2_7_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__6238\,
            in1 => \N__4730\,
            in2 => \N__4389\,
            in3 => \N__6008\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_a2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAB4_5_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__4868\,
            in1 => \_gnd_net_\,
            in2 => \N__4362\,
            in3 => \N__4359\,
            lcout => \U712_CHIP_RAM.N_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111001011110000"
        )
    port map (
            in0 => \N__6047\,
            in1 => \N__7010\,
            in2 => \N__5008\,
            in3 => \N__6179\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9514\,
            ce => 'H',
            sr => \N__9301\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__6178\,
            in1 => \N__6046\,
            in2 => \_gnd_net_\,
            in3 => \N__4799\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__5965\,
            in1 => \N__6905\,
            in2 => \N__4611\,
            in3 => \N__8272\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9514\,
            ce => 'H',
            sr => \N__9301\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111100011111010"
        )
    port map (
            in0 => \N__4595\,
            in1 => \N__5072\,
            in2 => \N__5145\,
            in3 => \N__6564\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9521\,
            ce => 'H',
            sr => \N__9285\
        );

    \U712_REG_SM.DS_EN_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100101110"
        )
    port map (
            in0 => \N__7265\,
            in1 => \N__4584\,
            in2 => \N__4575\,
            in3 => \N__4566\,
            lcout => \U712_REG_SM.DS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9522\,
            ce => 'H',
            sr => \N__9278\
        );

    \U712_REG_SM.C3_SYNC_2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4527\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9522\,
            ce => 'H',
            sr => \N__9278\
        );

    \U712_REG_SM.REG_TACK_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010111000"
        )
    port map (
            in0 => \N__4469\,
            in1 => \N__5397\,
            in2 => \N__5118\,
            in3 => \N__4491\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9522\,
            ce => 'H',
            sr => \N__9278\
        );

    \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4489\,
            in1 => \N__6594\,
            in2 => \_gnd_net_\,
            in3 => \N__6500\,
            lcout => \U712_REG_SM.N_167_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4559\,
            in1 => \N__4548\,
            in2 => \_gnd_net_\,
            in3 => \N__4523\,
            lcout => \U712_REG_SM.N_159_0\,
            ltout => \U712_REG_SM.N_159_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI0ULC2_4_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4473\,
            in3 => \N__4468\,
            lcout => \U712_REG_SM.N_165_0\,
            ltout => \U712_REG_SM.N_165_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__7981\,
            in1 => \N__5395\,
            in2 => \N__4683\,
            in3 => \N__4680\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9526\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111001100"
        )
    port map (
            in0 => \N__4632\,
            in1 => \N__7289\,
            in2 => \N__6964\,
            in3 => \N__4671\,
            lcout => \U712_REG_SM.UDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9529\,
            ce => 'H',
            sr => \N__9266\
        );

    \U712_REG_SM.LDS_OUT_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110100010"
        )
    port map (
            in0 => \N__4670\,
            in1 => \N__4638\,
            in2 => \N__6963\,
            in3 => \N__6383\,
            lcout => \U712_REG_SM.LDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9529\,
            ce => 'H',
            sr => \N__9266\
        );

    \U712_REG_SM.LDS_OUT_RNO_0_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5221\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5290\,
            lcout => \U712_REG_SM.LDS_OUT_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_RNO_0_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5291\,
            in1 => \N__5222\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.UDS_OUT_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001000"
        )
    port map (
            in0 => \N__6243\,
            in1 => \N__4899\,
            in2 => \N__6155\,
            in3 => \N__5734\,
            lcout => \U712_CHIP_RAM.N_105\,
            ltout => \U712_CHIP_RAM.N_105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI264TB_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011111111"
        )
    port map (
            in0 => \N__5747\,
            in1 => \N__5670\,
            in2 => \N__4626\,
            in3 => \N__5952\,
            lcout => \U712_CHIP_RAM.N_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100010001"
        )
    port map (
            in0 => \N__5953\,
            in1 => \N__5697\,
            in2 => \N__5681\,
            in3 => \N__4722\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8001\,
            in2 => \N__4623\,
            in3 => \N__4620\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__5496\,
            in1 => \_gnd_net_\,
            in2 => \N__4614\,
            in3 => \N__8640\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9494\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__5634\,
            in1 => \_gnd_net_\,
            in2 => \N__5922\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5918\,
            in2 => \_gnd_net_\,
            in3 => \N__5633\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6233\,
            in1 => \N__6125\,
            in2 => \_gnd_net_\,
            in3 => \N__4711\,
            lcout => \U712_CHIP_RAM.N_50\,
            ltout => \U712_CHIP_RAM.N_50_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__5901\,
            in1 => \_gnd_net_\,
            in2 => \N__4716\,
            in3 => \N__5629\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRB433_2_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101011110"
        )
    port map (
            in0 => \N__5630\,
            in1 => \N__6048\,
            in2 => \N__6257\,
            in3 => \N__5902\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_tz_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIT32E6_3_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011111111"
        )
    port map (
            in0 => \N__6126\,
            in1 => \N__4713\,
            in2 => \N__4695\,
            in3 => \N__5777\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHPUTC_3_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__4785\,
            in1 => \N__8000\,
            in2 => \N__4692\,
            in3 => \N__4764\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__7999\,
            in1 => \N__4689\,
            in2 => \_gnd_net_\,
            in3 => \N__5736\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__6237\,
            in1 => \N__5477\,
            in2 => \_gnd_net_\,
            in3 => \N__5801\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9497\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIMMGI5_2_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__5757\,
            in1 => \N__6241\,
            in2 => \N__6015\,
            in3 => \N__4763\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIP5G8C_2_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011101010"
        )
    port map (
            in0 => \N__4800\,
            in1 => \N__4784\,
            in2 => \N__4773\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIM9IMI_0_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__9362\,
            in1 => \N__5976\,
            in2 => \N__4770\,
            in3 => \N__5954\,
            lcout => \U712_CHIP_RAM.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6239\,
            in1 => \N__5618\,
            in2 => \N__6148\,
            in3 => \N__5693\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_92_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN7BL3_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__5756\,
            in1 => \N__6240\,
            in2 => \N__4767\,
            in3 => \N__5732\,
            lcout => \U712_CHIP_RAM.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_4_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6127\,
            in2 => \_gnd_net_\,
            in3 => \N__4752\,
            lcout => \U712_CHIP_RAM.BANK0_0_sqmuxa_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__5619\,
            in1 => \N__5887\,
            in2 => \_gnd_net_\,
            in3 => \N__5800\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9504\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__5731\,
            in1 => \N__6318\,
            in2 => \_gnd_net_\,
            in3 => \N__6294\,
            lcout => \U712_CHIP_RAM.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5680\,
            in1 => \N__6006\,
            in2 => \N__5917\,
            in3 => \N__5620\,
            lcout => \U712_CHIP_RAM.N_106\,
            ltout => \U712_CHIP_RAM.N_106_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI7Q5U5_0_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4935\,
            in3 => \N__6037\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_3_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__6275\,
            in1 => \N__6258\,
            in2 => \N__4932\,
            in3 => \N__6157\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010110011111100"
        )
    port map (
            in0 => \N__5911\,
            in1 => \N__5413\,
            in2 => \N__4929\,
            in3 => \N__7023\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9512\,
            ce => 'H',
            sr => \N__9294\
        );

    \U712_CHIP_RAM.CLK_EN_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011111110110000"
        )
    port map (
            in0 => \N__6864\,
            in1 => \N__5912\,
            in2 => \N__6081\,
            in3 => \N__4910\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9512\,
            ce => 'H',
            sr => \N__9294\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI72V93_0_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6007\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4894\,
            lcout => \U712_CHIP_RAM.N_70_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__7214\,
            in1 => \N__5966\,
            in2 => \N__4878\,
            in3 => \N__6906\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9512\,
            ce => 'H',
            sr => \N__9294\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJDDI_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5857\,
            in2 => \_gnd_net_\,
            in3 => \N__8239\,
            lcout => \U712_CHIP_RAM.CPU_TACK_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8240\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6070\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un6_CPU_CYCLE_START_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__4857\,
            in1 => \N__7967\,
            in2 => \N__4839\,
            in3 => \N__4832\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9515\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__7963\,
            in1 => \N__5124\,
            in2 => \N__5071\,
            in3 => \N__6818\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7965\,
            in2 => \_gnd_net_\,
            in3 => \N__5031\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__7966\,
            in1 => \_gnd_net_\,
            in2 => \N__5144\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5137\,
            in2 => \_gnd_net_\,
            in3 => \N__5030\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110111"
        )
    port map (
            in0 => \N__5097\,
            in1 => \N__6817\,
            in2 => \N__5117\,
            in3 => \N__6561\,
            lcout => \U712_CYCLE_TERM.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5110\,
            in2 => \_gnd_net_\,
            in3 => \N__5096\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__7962\,
            in1 => \N__6539\,
            in2 => \N__5079\,
            in3 => \N__6816\,
            lcout => \U712_CYCLE_TERM.N_45_0_0_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__6562\,
            in1 => \N__7964\,
            in2 => \_gnd_net_\,
            in3 => \N__5064\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9517\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_0_i_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110010"
        )
    port map (
            in0 => \N__7171\,
            in1 => \N__6972\,
            in2 => \N__7238\,
            in3 => \N__5015\,
            lcout => \DRDDIR_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011011101"
        )
    port map (
            in0 => \N__5466\,
            in1 => \N__7344\,
            in2 => \N__5328\,
            in3 => \N__8324\,
            lcout => \CLMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un3_CLLBEn_1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7233\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5422\,
            lcout => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1\,
            ltout => \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__7378\,
            in1 => \N__5337\,
            in2 => \N__5460\,
            in3 => \N__8323\,
            lcout => \CLLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un3_CUMBEn_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7234\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5423\,
            lcout => \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__5396\,
            in1 => \N__7170\,
            in2 => \N__5373\,
            in3 => \N__5348\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9523\,
            ce => 'H',
            sr => \N__9267\
        );

    \U712_BYTE_ENABLE.LLBE_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100100010"
        )
    port map (
            in0 => \N__5182\,
            in1 => \N__5263\,
            in2 => \N__5234\,
            in3 => \N__5314\,
            lcout => \U712_BYTE_ENABLE.LLBE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LMBE_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000110100010"
        )
    port map (
            in0 => \N__5183\,
            in1 => \N__5264\,
            in2 => \N__5235\,
            in3 => \N__5315\,
            lcout => \U712_BYTE_ENABLE.LMBE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000001100100"
        )
    port map (
            in0 => \N__5190\,
            in1 => \N__5316\,
            in2 => \N__5268\,
            in3 => \N__5232\,
            lcout => \U712_BYTE_ENABLE.UMBE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010010101000"
        )
    port map (
            in0 => \N__5313\,
            in1 => \N__5262\,
            in2 => \N__5233\,
            in3 => \N__5181\,
            lcout => \U712_BYTE_ENABLE.UUBE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100111"
        )
    port map (
            in0 => \N__8615\,
            in1 => \N__8835\,
            in2 => \N__8987\,
            in3 => \N__8537\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__6609\,
            in1 => \N__8616\,
            in2 => \N__8375\,
            in3 => \N__8019\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8346\,
            in1 => \N__5559\,
            in2 => \N__5541\,
            in3 => \N__5538\,
            lcout => \U712_CHIP_RAM.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8834\,
            in1 => \N__8962\,
            in2 => \N__8641\,
            in3 => \N__8535\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7994\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5504\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_78_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000011"
        )
    port map (
            in0 => \N__8536\,
            in1 => \N__5763\,
            in2 => \N__5511\,
            in3 => \N__5495\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5679\,
            in1 => \N__5748\,
            in2 => \_gnd_net_\,
            in3 => \N__7993\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_76_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101100000001"
        )
    port map (
            in0 => \N__5494\,
            in1 => \N__5784\,
            in2 => \N__5508\,
            in3 => \N__8963\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001110111"
        )
    port map (
            in0 => \N__5505\,
            in1 => \N__7992\,
            in2 => \N__8881\,
            in3 => \N__5493\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__6129\,
            in1 => \N__5478\,
            in2 => \N__6264\,
            in3 => \N__5802\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5778\,
            in1 => \N__5614\,
            in2 => \N__5682\,
            in3 => \N__6860\,
            lcout => \U712_CHIP_RAM.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7991\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6010\,
            lcout => \U712_CHIP_RAM.N_99\,
            ltout => \U712_CHIP_RAM.N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__5677\,
            in1 => \_gnd_net_\,
            in2 => \N__5766\,
            in3 => \N__5613\,
            lcout => \U712_CHIP_RAM.N_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6128\,
            in2 => \_gnd_net_\,
            in3 => \N__5611\,
            lcout => \U712_CHIP_RAM.N_93_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8836\,
            in1 => \N__8633\,
            in2 => \_gnd_net_\,
            in3 => \N__8967\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMT791_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001010101"
        )
    port map (
            in0 => \N__5897\,
            in1 => \N__5612\,
            in2 => \_gnd_net_\,
            in3 => \N__5733\,
            lcout => \U712_CHIP_RAM.N_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__5730\,
            in1 => \N__6316\,
            in2 => \_gnd_net_\,
            in3 => \N__6291\,
            lcout => \U712_CHIP_RAM.N_54\,
            ltout => \U712_CHIP_RAM.N_54_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000001"
        )
    port map (
            in0 => \N__5886\,
            in1 => \N__5678\,
            in2 => \N__5637\,
            in3 => \N__5631\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNO_0_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__6333\,
            in1 => \N__6072\,
            in2 => \_gnd_net_\,
            in3 => \N__8357\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH_CYCLE_START_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__7229\,
            in1 => \N__6904\,
            in2 => \N__6321\,
            in3 => \N__7998\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__5961\,
            in1 => \N__6317\,
            in2 => \_gnd_net_\,
            in3 => \N__6292\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH_CYCLE_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__6293\,
            in1 => \N__7997\,
            in2 => \N__6303\,
            in3 => \N__6300\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9498\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__6276\,
            in1 => \N__6259\,
            in2 => \N__6180\,
            in3 => \N__6156\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER53_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__6586\,
            in1 => \N__6894\,
            in2 => \N__6071\,
            in3 => \N__6493\,
            lcout => \U712_CHIP_RAM.N_40\,
            ltout => \U712_CHIP_RAM.N_40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6018\,
            in3 => \N__6011\,
            lcout => \U712_CHIP_RAM.N_59\,
            ltout => \U712_CHIP_RAM.N_59_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101010100"
        )
    port map (
            in0 => \N__9359\,
            in1 => \N__5888\,
            in2 => \N__5970\,
            in3 => \N__5967\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9505\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9357\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5808\,
            lcout => \U712_CYCLE_TERM.N_45_0_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9356\,
            in2 => \_gnd_net_\,
            in3 => \N__6600\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6492\,
            lcout => \U712_REG_SM_DBR_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9516\,
            ce => 'H',
            sr => \N__9271\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010001010000"
        )
    port map (
            in0 => \N__6563\,
            in1 => \N__6830\,
            in2 => \N__6543\,
            in3 => \N__6528\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9516\,
            ce => 'H',
            sr => \N__9271\
        );

    \U712_CHIP_RAM.DBR_SYNC_0_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6522\,
            lcout => \U712_REG_SM_DBR_SYNC_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9518\,
            ce => 'H',
            sr => \N__9268\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__6419\,
            in1 => \N__7386\,
            in2 => \N__8391\,
            in3 => \N__6462\,
            lcout => \CUMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110101"
        )
    port map (
            in0 => \N__8390\,
            in1 => \N__7337\,
            in2 => \N__6432\,
            in3 => \N__6420\,
            lcout => \CUUBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_RNIL31J_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6390\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7277\,
            lcout => \U712_REG_SM_un1_LDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__8890\,
            in1 => \N__9005\,
            in2 => \_gnd_net_\,
            in3 => \N__6639\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9479\,
            ce => \N__9081\,
            sr => \N__9313\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__6765\,
            in1 => \_gnd_net_\,
            in2 => \N__9021\,
            in3 => \N__8891\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9479\,
            ce => \N__9081\,
            sr => \N__9313\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__6747\,
            in1 => \N__6633\,
            in2 => \N__6729\,
            in3 => \N__8345\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__8854\,
            in1 => \_gnd_net_\,
            in2 => \N__6705\,
            in3 => \N__8986\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9482\,
            ce => \N__9064\,
            sr => \N__9310\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__6618\,
            in1 => \N__8343\,
            in2 => \N__8710\,
            in3 => \N__8415\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8344\,
            in1 => \N__6678\,
            in2 => \N__6660\,
            in3 => \N__6657\,
            lcout => \U712_CHIP_RAM.N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__7494\,
            in1 => \N__8377\,
            in2 => \N__6627\,
            in3 => \N__8666\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7487\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9489\,
            ce => \N__7409\,
            sr => \N__9295\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7517\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9489\,
            ce => \N__7409\,
            sr => \N__9295\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8454\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9489\,
            ce => \N__7409\,
            sr => \N__9295\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8055\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9489\,
            ce => \N__7409\,
            sr => \N__9295\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9358\,
            in2 => \_gnd_net_\,
            in3 => \N__6779\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110101"
        )
    port map (
            in0 => \N__7065\,
            in1 => \N__9144\,
            in2 => \N__8378\,
            in3 => \N__8694\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8356\,
            in1 => \N__7059\,
            in2 => \N__7041\,
            in3 => \N__7038\,
            lcout => \U712_CHIP_RAM.N_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7425\,
            in2 => \_gnd_net_\,
            in3 => \N__6895\,
            lcout => \U712_CHIP_RAM.DBENn_7_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__7225\,
            in1 => \N__6896\,
            in2 => \N__6783\,
            in3 => \N__7982\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9499\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__7014\,
            in1 => \N__6962\,
            in2 => \_gnd_net_\,
            in3 => \N__6903\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9506\,
            ce => \N__6843\,
            sr => \N__9272\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__7937\,
            in1 => \N__6834\,
            in2 => \_gnd_net_\,
            in3 => \N__6819\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9513\,
            ce => \N__6789\,
            sr => \N__9269\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNILUVG_1_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7299\,
            in2 => \_gnd_net_\,
            in3 => \N__7310\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7385\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7336\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9519\,
            ce => 'H',
            sr => \N__9264\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7311\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9519\,
            ce => 'H',
            sr => \N__9264\
        );

    \U712_REG_SM.UDS_OUT_RNIUP9B_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__7293\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7278\,
            lcout => \U712_REG_SM_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7239\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7184\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7419\,
            in1 => \N__8373\,
            in2 => \N__8709\,
            in3 => \N__7449\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8374\,
            in1 => \N__7110\,
            in2 => \N__7092\,
            in3 => \N__7089\,
            lcout => \U712_CHIP_RAM.N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9360\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7074\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7518\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9481\,
            ce => \N__8774\,
            sr => \N__9292\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7488\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9481\,
            ce => \N__8774\,
            sr => \N__9292\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000001"
        )
    port map (
            in0 => \N__8897\,
            in1 => \N__9019\,
            in2 => \N__8718\,
            in3 => \N__7443\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9484\,
            ce => \N__9080\,
            sr => \N__9283\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8097\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9487\,
            ce => \N__7410\,
            sr => \N__9276\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9171\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9487\,
            ce => \N__7410\,
            sr => \N__9276\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8126\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9487\,
            ce => \N__7410\,
            sr => \N__9276\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8487\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9487\,
            ce => \N__7410\,
            sr => \N__9276\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8169\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9487\,
            ce => \N__7410\,
            sr => \N__9276\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7392\,
            in1 => \N__8314\,
            in2 => \N__8698\,
            in3 => \N__8460\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7897\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__7698\,
            in1 => \N__8895\,
            in2 => \_gnd_net_\,
            in3 => \N__9018\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9480\,
            ce => \N__9096\,
            sr => \N__9314\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000001"
        )
    port map (
            in0 => \N__9017\,
            in1 => \N__8896\,
            in2 => \N__8714\,
            in3 => \N__7785\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9480\,
            ce => \N__9096\,
            sr => \N__9314\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7755\,
            in1 => \N__8369\,
            in2 => \N__8716\,
            in3 => \N__8064\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8370\,
            in1 => \N__7746\,
            in2 => \N__7725\,
            in3 => \N__7722\,
            lcout => \U712_CHIP_RAM.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__7692\,
            in1 => \N__7635\,
            in2 => \N__8142\,
            in3 => \N__8379\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9485\,
            ce => \N__9091\,
            sr => \N__9302\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__7524\,
            in1 => \N__8901\,
            in2 => \_gnd_net_\,
            in3 => \N__9020\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9490\,
            ce => \N__9095\,
            sr => \N__9296\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__9585\,
            in1 => \N__7634\,
            in2 => \N__7614\,
            in3 => \N__8380\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9490\,
            ce => \N__9095\,
            sr => \N__9296\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__7575\,
            in1 => \N__7554\,
            in2 => \N__7548\,
            in3 => \N__8376\,
            lcout => \U712_CHIP_RAM.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8483\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9500\,
            ce => \N__8765\,
            sr => \N__9279\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8450\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9500\,
            ce => \N__8765\,
            sr => \N__9279\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__8403\,
            in1 => \N__8371\,
            in2 => \N__8715\,
            in3 => \N__8103\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8372\,
            in1 => \N__8202\,
            in2 => \N__8187\,
            in3 => \N__8184\,
            lcout => \U712_CHIP_RAM.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8168\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9491\,
            ce => \N__8775\,
            sr => \N__9311\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8133\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9491\,
            ce => \N__8775\,
            sr => \N__9311\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8093\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9496\,
            ce => \N__8770\,
            sr => \N__9303\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8048\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9496\,
            ce => \N__8770\,
            sr => \N__9303\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9167\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9501\,
            ce => \N__8769\,
            sr => \N__9297\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100011001000"
        )
    port map (
            in0 => \N__8899\,
            in1 => \N__9135\,
            in2 => \N__9030\,
            in3 => \_gnd_net_\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9492\,
            ce => \N__9065\,
            sr => \N__9318\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8898\,
            in1 => \N__8708\,
            in2 => \N__9029\,
            in3 => \N__8550\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9492\,
            ce => \N__9065\,
            sr => \N__9318\
        );

    \U712_CHIP_RAM.WEn_LC_16_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9028\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9483\,
            ce => 'H',
            sr => \N__9321\
        );

    \U712_CHIP_RAM.RASn_LC_16_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8900\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9493\,
            ce => 'H',
            sr => \N__9319\
        );

    \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9361\,
            in1 => \N__9543\,
            in2 => \_gnd_net_\,
            in3 => \N__9554\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_17_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8717\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9486\,
            ce => 'H',
            sr => \N__9322\
        );

    \U712_CHIP_RAM.CRCSn_LC_17_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8549\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9502\,
            ce => 'H',
            sr => \N__9320\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8499\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9581\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9520\,
            ce => 'H',
            sr => \N__9312\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9555\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9520\,
            ce => 'H',
            sr => \N__9312\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 14 2024 11:09:01

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U111_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U111_TOP
entity U111_TOP is
port (
    D_LL_AMIGA : inout std_logic_vector(7 downto 0);
    D_LM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_AMIGA : inout std_logic_vector(7 downto 0);
    D_UM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_040 : inout std_logic_vector(7 downto 0);
    D_LL_040 : inout std_logic_vector(7 downto 0);
    D_LM_040 : inout std_logic_vector(7 downto 0);
    D_UM_040 : inout std_logic_vector(7 downto 0);
    A_AMIGA : out std_logic_vector(1 downto 0);
    A_040 : in std_logic_vector(1 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    TSn : out std_logic;
    RESETn : in std_logic;
    CLKRAMA : out std_logic;
    PORTSIZE : in std_logic;
    CLK40B : out std_logic;
    TBI_CPUn : out std_logic;
    TAn : out std_logic;
    CPUBGn : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CLK80_CPU : out std_logic;
    BUFDIR : out std_logic;
    TCI_CPUn : out std_logic;
    TS_CPUn : in std_logic;
    CLKRAMB : out std_logic;
    CLK40A : out std_logic;
    DMAn : out std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    TACKn : in std_logic;
    BGn : in std_logic);
end U111_TOP;

-- Architecture of U111_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U111_TOP is

signal \N__7858\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3625\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2959\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2875\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2461\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2449\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2222\ : std_logic;
signal \N__2219\ : std_logic;
signal \N__2216\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2198\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \A_040_c_1\ : std_logic;
signal \A_040_c_0\ : std_logic;
signal \A_AMIGA_c_0\ : std_logic;
signal \D_LL_AMIGA_in_2\ : std_logic;
signal \un1_D_LL_AMIGA_2\ : std_logic;
signal \D_LM_AMIGA_in_2\ : std_logic;
signal \un1_D_LM_AMIGA_2\ : std_logic;
signal \D_UM_040_in_1\ : std_logic;
signal \D_LL_040_in_1\ : std_logic;
signal \un1_D_UM_040_1\ : std_logic;
signal \RnW_c_i_0\ : std_logic;
signal \D_LM_AMIGA_in_4\ : std_logic;
signal \un1_D_LM_AMIGA_4\ : std_logic;
signal \D_LM_AMIGA_in_5\ : std_logic;
signal \un1_D_LM_AMIGA_5\ : std_logic;
signal \D_LM_AMIGA_in_6\ : std_logic;
signal \un1_D_LM_AMIGA_6\ : std_logic;
signal \D_UU_040_in_3\ : std_logic;
signal \D_LM_040_in_3\ : std_logic;
signal \un1_D_UU_040_3\ : std_logic;
signal \D_LL_AMIGA_in_0\ : std_logic;
signal \un1_D_LL_AMIGA_0\ : std_logic;
signal \D_LL_AMIGA_in_1\ : std_logic;
signal \un1_D_LL_AMIGA_1\ : std_logic;
signal \D_LM_AMIGA_in_3\ : std_logic;
signal \un1_D_LM_AMIGA_3\ : std_logic;
signal \D_LM_AMIGA_in_7\ : std_logic;
signal \un1_D_LM_AMIGA_7\ : std_logic;
signal \A_AMIGA_c_1\ : std_logic;
signal \D_UM_040_in_7\ : std_logic;
signal \D_LL_040_in_7\ : std_logic;
signal \un1_D_UM_040_7\ : std_logic;
signal \D_LM_040_in_6\ : std_logic;
signal \D_UU_040_in_6\ : std_logic;
signal \un1_D_UU_040_6\ : std_logic;
signal \D_LL_AMIGA_in_3\ : std_logic;
signal \un1_D_LL_AMIGA_3\ : std_logic;
signal \un1_D_UM_AMIGA_0\ : std_logic;
signal \D_UM_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net\ : std_logic;
signal \INVU111_CYCLE_SM.TA_EN_nessC_net\ : std_logic;
signal \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\ : std_logic;
signal \D_LM_040_in_1\ : std_logic;
signal \D_UU_040_in_1\ : std_logic;
signal \un1_D_UU_040_1\ : std_logic;
signal \D_UU_AMIGA_in_6\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\ : std_logic;
signal \un1_D_UU_AMIGA_6\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\ : std_logic;
signal \D_UU_AMIGA_in_4\ : std_logic;
signal \un1_D_UU_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\ : std_logic;
signal \D_UU_AMIGA_in_7\ : std_logic;
signal \un1_D_UU_AMIGA_7\ : std_logic;
signal \D_LL_AMIGA_in_4\ : std_logic;
signal \un1_D_LL_AMIGA_4\ : std_logic;
signal \D_LM_AMIGA_in_0\ : std_logic;
signal \un1_D_LM_AMIGA_0\ : std_logic;
signal \D_LM_AMIGA_in_1\ : std_logic;
signal \un1_D_LM_AMIGA_1\ : std_logic;
signal \INVU111_CYCLE_SM.TSnC_net\ : std_logic;
signal \U111_CYCLE_SM.A_OUTZ0\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLE_r_1_cascade_\ : std_logic;
signal \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\ : std_logic;
signal \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_cascade_\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_0\ : std_logic;
signal \U111_CYCLE_SM.TS_EN10\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLE_STARTZ0\ : std_logic;
signal \INVU111_CYCLE_SM.A_OUTC_net\ : std_logic;
signal \INVU111_CYCLE_SM.CYCLE_STATE_0C_net\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\ : std_logic;
signal \D_UM_AMIGA_in_1\ : std_logic;
signal \un1_D_UM_AMIGA_1\ : std_logic;
signal \D_UU_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\ : std_logic;
signal \un1_D_UU_AMIGA_1\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\ : std_logic;
signal \D_UM_AMIGA_in_4\ : std_logic;
signal \un1_D_UM_AMIGA_4\ : std_logic;
signal \D_UU_040_in_0\ : std_logic;
signal \D_LM_040_in_0\ : std_logic;
signal \un1_D_UU_040_0\ : std_logic;
signal \D_UU_040_in_2\ : std_logic;
signal \D_LM_040_in_2\ : std_logic;
signal \un1_D_UU_040_2\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\ : std_logic;
signal \D_UU_AMIGA_in_0\ : std_logic;
signal \un1_D_UU_AMIGA_0\ : std_logic;
signal \D_LL_AMIGA_in_6\ : std_logic;
signal \un1_D_LL_AMIGA_6\ : std_logic;
signal \D_LL_AMIGA_in_5\ : std_logic;
signal \un1_D_LL_AMIGA_5\ : std_logic;
signal \D_LL_AMIGA_in_7\ : std_logic;
signal \un1_D_LL_AMIGA_7\ : std_logic;
signal \D_UM_040_in_2\ : std_logic;
signal \D_LL_040_in_2\ : std_logic;
signal \un1_D_UM_040_2\ : std_logic;
signal \un1_D_UM_AMIGA_2\ : std_logic;
signal \D_UM_AMIGA_in_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\ : std_logic;
signal \U111_CYCLE_SM.TA_ENZ0\ : std_logic;
signal \TACKn_c\ : std_logic;
signal \TAn_0_i\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\ : std_logic;
signal \TS_CPUn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\ : std_logic;
signal \U111_CYCLE_SM.TS_EN_4\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\ : std_logic;
signal \D_UM_AMIGA_in_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\ : std_logic;
signal \un1_D_UM_AMIGA_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\ : std_logic;
signal \D_UM_AMIGA_in_7\ : std_logic;
signal \un1_D_UM_AMIGA_7\ : std_logic;
signal \D_LL_040_in_4\ : std_logic;
signal \D_UM_040_in_4\ : std_logic;
signal \un1_D_UM_040_4\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\ : std_logic;
signal \D_UU_AMIGA_in_3\ : std_logic;
signal \un1_D_UU_AMIGA_3\ : std_logic;
signal \D_UM_040_in_5\ : std_logic;
signal \D_LL_040_in_5\ : std_logic;
signal \un1_D_UM_040_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\ : std_logic;
signal \D_UU_AMIGA_in_5\ : std_logic;
signal \un1_D_UU_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\ : std_logic;
signal \D_UU_AMIGA_in_2\ : std_logic;
signal \un1_D_UU_AMIGA_2\ : std_logic;
signal \D_UM_AMIGA_in_5\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\ : std_logic;
signal \un1_D_UM_AMIGA_5\ : std_logic;
signal \CLK40\ : std_logic;
signal \GB_BUFFER_CLK40_THRU_CO\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLEZ0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\ : std_logic;
signal \D_UM_AMIGA_in_6\ : std_logic;
signal \un1_D_UM_AMIGA_6\ : std_logic;
signal \CLK80\ : std_logic;
signal \GB_BUFFER_CLK80_THRU_CO\ : std_logic;
signal \D_LM_040_in_5\ : std_logic;
signal \D_UU_040_in_5\ : std_logic;
signal \un1_D_UU_040_5\ : std_logic;
signal \D_LM_040_in_7\ : std_logic;
signal \D_UU_040_in_7\ : std_logic;
signal \un1_D_UU_040_7\ : std_logic;
signal \D_UM_040_in_0\ : std_logic;
signal \D_LL_040_in_0\ : std_logic;
signal \un1_D_UM_040_0\ : std_logic;
signal \D_LL_040_in_6\ : std_logic;
signal \D_UM_040_in_6\ : std_logic;
signal \un1_D_UM_040_6\ : std_logic;
signal \D_LL_040_in_3\ : std_logic;
signal \D_UM_040_in_3\ : std_logic;
signal \un1_D_UM_040_3\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \PORTSIZE_c\ : std_logic;
signal \U111_CYCLE_SM.LW_TRANS_0\ : std_logic;
signal \D_UU_040_in_4\ : std_logic;
signal \U111_CYCLE_SM.FLIP\ : std_logic;
signal \D_LM_040_in_4\ : std_logic;
signal \un1_D_UU_040_4\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \CPUBGn_wire\ : std_logic;
signal \A_040_wire\ : std_logic_vector(1 downto 0);
signal \A_AMIGA_wire\ : std_logic_vector(1 downto 0);
signal \CLK40B_wire\ : std_logic;
signal \TBI_CPUn_wire\ : std_logic;
signal \CLK40A_wire\ : std_logic;
signal \BUFDIR_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \TS_CPUn_wire\ : std_logic;
signal \CLKRAMA_wire\ : std_logic;
signal \TCI_CPUn_wire\ : std_logic;
signal \CLKRAMB_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \TAn_wire\ : std_logic;
signal \DMAn_wire\ : std_logic;
signal \CLK80_CPU_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \pll_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \TACKn_wire\ <= TACKn;
    CPUBGn <= \CPUBGn_wire\;
    \A_040_wire\ <= A_040;
    A_AMIGA <= \A_AMIGA_wire\;
    CLK40B <= \CLK40B_wire\;
    TBI_CPUn <= \TBI_CPUn_wire\;
    CLK40A <= \CLK40A_wire\;
    BUFDIR <= \BUFDIR_wire\;
    \SIZ_wire\ <= SIZ;
    \TS_CPUn_wire\ <= TS_CPUn;
    CLKRAMA <= \CLKRAMA_wire\;
    TCI_CPUn <= \TCI_CPUn_wire\;
    CLKRAMB <= \CLKRAMB_wire\;
    BUFENn <= \BUFENn_wire\;
    \RnW_wire\ <= RnW;
    TAn <= \TAn_wire\;
    DMAn <= \DMAn_wire\;
    CLK80_CPU <= \CLK80_CPU_wire\;
    TSn <= \TSn_wire\;
    \PORTSIZE_wire\ <= PORTSIZE;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    \pll_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_pll\ : PLL40_2F
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            SCLK => '0',
            PLLOUTGLOBALA => \CLK80\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALB => \CLK40\,
            SDI => '0',
            PLLOUTCOREA => OPEN,
            BYPASS => '0',
            RESETB => \N__7030\,
            PLLOUTCOREB => OPEN,
            LOCK => OPEN,
            SDO => OPEN,
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \pll_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__7858\
        );

    \pll_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__7858\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \D_UM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7842\,
            DIN => \N__7841\,
            DOUT => \N__7840\,
            PACKAGEPIN => D_UM_040(3)
        );

    \D_UM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7842\,
            PADOUT => \N__7841\,
            PADIN => \N__7840\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3889\,
            DIN0 => \D_UM_040_in_3\,
            DOUT0 => \N__5078\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7833\,
            DIN => \N__7832\,
            DOUT => \N__7831\,
            PACKAGEPIN => D_LL_AMIGA(1)
        );

    \D_LL_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7833\,
            PADOUT => \N__7832\,
            PADIN => \N__7831\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2822\,
            DIN0 => \D_LL_AMIGA_in_1\,
            DOUT0 => \N__2905\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7824\,
            DIN => \N__7823\,
            DOUT => \N__7822\,
            PACKAGEPIN => D_UU_AMIGA(5)
        );

    \D_UU_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7824\,
            PADOUT => \N__7823\,
            PADIN => \N__7822\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2819\,
            DIN0 => \D_UU_AMIGA_in_5\,
            DOUT0 => \N__6809\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7815\,
            DIN => \N__7814\,
            DOUT => \N__7813\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7815\,
            PADOUT => \N__7814\,
            PADIN => \N__7813\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TACKn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7806\,
            DIN => \N__7805\,
            DOUT => \N__7804\,
            PACKAGEPIN => D_UU_040(6)
        );

    \D_UU_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7806\,
            PADOUT => \N__7805\,
            PADIN => \N__7804\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3936\,
            DIN0 => \D_UU_040_in_6\,
            DOUT0 => \N__3449\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUBGn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7797\,
            DIN => \N__7796\,
            DOUT => \N__7795\,
            PACKAGEPIN => \CPUBGn_wire\
        );

    \CPUBGn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7797\,
            PADOUT => \N__7796\,
            PADIN => \N__7795\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7788\,
            DIN => \N__7787\,
            DOUT => \N__7786\,
            PACKAGEPIN => D_LL_040(7)
        );

    \D_LL_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7788\,
            PADOUT => \N__7787\,
            PADIN => \N__7786\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4003\,
            DIN0 => \D_LL_040_in_7\,
            DOUT0 => \N__4916\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7779\,
            DIN => \N__7778\,
            DOUT => \N__7777\,
            PACKAGEPIN => D_LL_AMIGA(4)
        );

    \D_LL_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7779\,
            PADOUT => \N__7778\,
            PADIN => \N__7777\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2821\,
            DIN0 => \D_LL_AMIGA_in_4\,
            DOUT0 => \N__6031\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7770\,
            DIN => \N__7769\,
            DOUT => \N__7768\,
            PACKAGEPIN => D_UM_AMIGA(3)
        );

    \D_UM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7770\,
            PADOUT => \N__7769\,
            PADIN => \N__7768\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2779\,
            DIN0 => \D_UM_AMIGA_in_3\,
            DOUT0 => \N__6503\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7761\,
            DIN => \N__7760\,
            DOUT => \N__7759\,
            PACKAGEPIN => D_UU_040(3)
        );

    \D_UU_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7761\,
            PADOUT => \N__7760\,
            PADIN => \N__7759\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3931\,
            DIN0 => \D_UU_040_in_3\,
            DOUT0 => \N__5894\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7752\,
            DIN => \N__7751\,
            DOUT => \N__7750\,
            PACKAGEPIN => \A_040_wire\(1)
        );

    \A_040_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7752\,
            PADOUT => \N__7751\,
            PADIN => \N__7750\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7743\,
            DIN => \N__7742\,
            DOUT => \N__7741\,
            PACKAGEPIN => D_LM_AMIGA(3)
        );

    \D_LM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7743\,
            PADOUT => \N__7742\,
            PADIN => \N__7741\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2617\,
            DIN0 => \D_LM_AMIGA_in_3\,
            DOUT0 => \N__2471\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7734\,
            DIN => \N__7733\,
            DOUT => \N__7732\,
            PACKAGEPIN => D_LM_040(0)
        );

    \D_LM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7734\,
            PADOUT => \N__7733\,
            PADIN => \N__7732\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4004\,
            DIN0 => \D_LM_040_in_0\,
            DOUT0 => \N__3704\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7725\,
            DIN => \N__7724\,
            DOUT => \N__7723\,
            PACKAGEPIN => D_UM_AMIGA(6)
        );

    \D_UM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7725\,
            PADOUT => \N__7724\,
            PADIN => \N__7723\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2818\,
            DIN0 => \D_UM_AMIGA_in_6\,
            DOUT0 => \N__6581\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7716\,
            DIN => \N__7715\,
            DOUT => \N__7714\,
            PACKAGEPIN => D_LM_AMIGA(4)
        );

    \D_LM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7716\,
            PADOUT => \N__7715\,
            PADIN => \N__7714\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2674\,
            DIN0 => \D_LM_AMIGA_in_4\,
            DOUT0 => \N__6095\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7707\,
            DIN => \N__7706\,
            DOUT => \N__7705\,
            PACKAGEPIN => \A_AMIGA_wire\(1)
        );

    \A_AMIGA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7707\,
            PADOUT => \N__7706\,
            PADIN => \N__7705\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3205\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7698\,
            DIN => \N__7697\,
            DOUT => \N__7696\,
            PACKAGEPIN => D_LM_040(7)
        );

    \D_LM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7698\,
            PADOUT => \N__7697\,
            PADIN => \N__7696\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3812\,
            DIN0 => \D_LM_040_in_7\,
            DOUT0 => \N__3230\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7689\,
            DIN => \N__7688\,
            DOUT => \N__7687\,
            PACKAGEPIN => D_UM_040(4)
        );

    \D_UM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7689\,
            PADOUT => \N__7688\,
            PADIN => \N__7687\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3932\,
            DIN0 => \D_UM_040_in_4\,
            DOUT0 => \N__4376\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7680\,
            DIN => \N__7679\,
            DOUT => \N__7678\,
            PACKAGEPIN => \CLK40B_wire\
        );

    \CLK40B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7680\,
            PADOUT => \N__7679\,
            PADIN => \N__7678\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5546\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7671\,
            DIN => \N__7670\,
            DOUT => \N__7669\,
            PACKAGEPIN => D_UU_AMIGA(0)
        );

    \D_UU_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7671\,
            PADOUT => \N__7670\,
            PADIN => \N__7669\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2834\,
            DIN0 => \D_UU_AMIGA_in_0\,
            DOUT0 => \N__4292\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7662\,
            DIN => \N__7661\,
            DOUT => \N__7660\,
            PACKAGEPIN => \A_040_wire\(0)
        );

    \A_040_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7662\,
            PADOUT => \N__7661\,
            PADIN => \N__7660\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7653\,
            DIN => \N__7652\,
            DOUT => \N__7651\,
            PACKAGEPIN => D_LM_AMIGA(0)
        );

    \D_LM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7653\,
            PADOUT => \N__7652\,
            PADIN => \N__7651\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2783\,
            DIN0 => \D_LM_AMIGA_in_0\,
            DOUT0 => \N__4334\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7644\,
            DIN => \N__7643\,
            DOUT => \N__7642\,
            PACKAGEPIN => D_UM_040(1)
        );

    \D_UM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7644\,
            PADOUT => \N__7643\,
            PADIN => \N__7642\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3887\,
            DIN0 => \D_UM_040_in_1\,
            DOUT0 => \N__4520\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7635\,
            DIN => \N__7634\,
            DOUT => \N__7633\,
            PACKAGEPIN => \TBI_CPUn_wire\
        );

    \TBI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7635\,
            PADOUT => \N__7634\,
            PADIN => \N__7633\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7626\,
            DIN => \N__7625\,
            DOUT => \N__7624\,
            PACKAGEPIN => \CLK40A_wire\
        );

    \CLK40A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7626\,
            PADOUT => \N__7625\,
            PADIN => \N__7624\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5545\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7617\,
            DIN => \N__7616\,
            DOUT => \N__7615\,
            PACKAGEPIN => D_LM_040(3)
        );

    \D_LM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7617\,
            PADOUT => \N__7616\,
            PADIN => \N__7615\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3923\,
            DIN0 => \D_LM_040_in_3\,
            DOUT0 => \N__2324\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7608\,
            DIN => \N__7607\,
            DOUT => \N__7606\,
            PACKAGEPIN => D_LL_040(4)
        );

    \D_LL_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7608\,
            PADOUT => \N__7607\,
            PADIN => \N__7606\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4020\,
            DIN0 => \D_LL_040_in_4\,
            DOUT0 => \N__3266\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7599\,
            DIN => \N__7598\,
            DOUT => \N__7597\,
            PACKAGEPIN => D_LL_AMIGA(7)
        );

    \D_LL_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7599\,
            PADOUT => \N__7598\,
            PADIN => \N__7597\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2782\,
            DIN0 => \D_LL_AMIGA_in_7\,
            DOUT0 => \N__3173\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7590\,
            DIN => \N__7589\,
            DOUT => \N__7588\,
            PACKAGEPIN => D_UU_AMIGA(7)
        );

    \D_UU_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7590\,
            PADOUT => \N__7589\,
            PADIN => \N__7588\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2836\,
            DIN0 => \D_UU_AMIGA_in_7\,
            DOUT0 => \N__6734\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7581\,
            DIN => \N__7580\,
            DOUT => \N__7579\,
            PACKAGEPIN => \BUFDIR_wire\
        );

    \BUFDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7581\,
            PADOUT => \N__7580\,
            PADIN => \N__7579\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4002\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7572\,
            DIN => \N__7571\,
            DOUT => \N__7570\,
            PACKAGEPIN => D_LM_AMIGA(5)
        );

    \D_LM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7572\,
            PADOUT => \N__7571\,
            PADIN => \N__7570\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2710\,
            DIN0 => \D_LM_AMIGA_in_5\,
            DOUT0 => \N__6878\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7563\,
            DIN => \N__7562\,
            DOUT => \N__7561\,
            PACKAGEPIN => D_UU_040(4)
        );

    \D_UU_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7563\,
            PADOUT => \N__7562\,
            PADIN => \N__7561\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3970\,
            DIN0 => \D_UU_040_in_4\,
            DOUT0 => \N__3374\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7554\,
            DIN => \N__7553\,
            DOUT => \N__7552\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7554\,
            PADOUT => \N__7553\,
            PADIN => \N__7552\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7545\,
            DIN => \N__7544\,
            DOUT => \N__7543\,
            PACKAGEPIN => D_LM_040(6)
        );

    \D_LM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7545\,
            PADOUT => \N__7544\,
            PADIN => \N__7543\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3792\,
            DIN0 => \D_LM_040_in_6\,
            DOUT0 => \N__2516\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7536\,
            DIN => \N__7535\,
            DOUT => \N__7534\,
            PACKAGEPIN => D_UM_040(5)
        );

    \D_UM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7536\,
            PADOUT => \N__7535\,
            PADIN => \N__7534\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3933\,
            DIN0 => \D_UM_040_in_5\,
            DOUT0 => \N__5591\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TS_CPUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7527\,
            DIN => \N__7526\,
            DOUT => \N__7525\,
            PACKAGEPIN => \TS_CPUn_wire\
        );

    \TS_CPUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7527\,
            PADOUT => \N__7526\,
            PADIN => \N__7525\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TS_CPUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7518\,
            DIN => \N__7517\,
            DOUT => \N__7516\,
            PACKAGEPIN => D_LL_040(1)
        );

    \D_LL_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7518\,
            PADOUT => \N__7517\,
            PADIN => \N__7516\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4019\,
            DIN0 => \D_LL_040_in_1\,
            DOUT0 => \N__2363\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7509\,
            DIN => \N__7508\,
            DOUT => \N__7507\,
            PACKAGEPIN => D_LL_AMIGA(3)
        );

    \D_LL_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7509\,
            PADOUT => \N__7508\,
            PADIN => \N__7507\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2838\,
            DIN0 => \D_LL_AMIGA_in_3\,
            DOUT0 => \N__6565\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7500\,
            DIN => \N__7499\,
            DOUT => \N__7498\,
            PACKAGEPIN => D_UM_AMIGA(5)
        );

    \D_UM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7500\,
            PADOUT => \N__7499\,
            PADIN => \N__7498\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2835\,
            DIN0 => \D_UM_AMIGA_in_5\,
            DOUT0 => \N__5807\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7491\,
            DIN => \N__7490\,
            DOUT => \N__7489\,
            PACKAGEPIN => D_UU_040(1)
        );

    \D_UU_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7491\,
            PADOUT => \N__7490\,
            PADIN => \N__7489\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3890\,
            DIN0 => \D_UU_040_in_1\,
            DOUT0 => \N__4454\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7482\,
            DIN => \N__7481\,
            DOUT => \N__7480\,
            PACKAGEPIN => D_UU_AMIGA(3)
        );

    \D_UU_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7482\,
            PADOUT => \N__7481\,
            PADIN => \N__7480\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2820\,
            DIN0 => \D_UU_AMIGA_in_3\,
            DOUT0 => \N__2426\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7473\,
            DIN => \N__7472\,
            DOUT => \N__7471\,
            PACKAGEPIN => D_LM_AMIGA(1)
        );

    \D_LM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7473\,
            PADOUT => \N__7472\,
            PADIN => \N__7471\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2671\,
            DIN0 => \D_LM_AMIGA_in_1\,
            DOUT0 => \N__3580\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7464\,
            DIN => \N__7463\,
            DOUT => \N__7462\,
            PACKAGEPIN => D_LM_040(2)
        );

    \D_LM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7464\,
            PADOUT => \N__7463\,
            PADIN => \N__7462\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3978\,
            DIN0 => \D_LM_040_in_2\,
            DOUT0 => \N__2213\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7455\,
            DIN => \N__7454\,
            DOUT => \N__7453\,
            PACKAGEPIN => D_LL_040(5)
        );

    \D_LL_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7455\,
            PADOUT => \N__7454\,
            PADIN => \N__7453\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4005\,
            DIN0 => \D_LL_040_in_5\,
            DOUT0 => \N__4955\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7446\,
            DIN => \N__7445\,
            DOUT => \N__7444\,
            PACKAGEPIN => D_LL_AMIGA(6)
        );

    \D_LL_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7446\,
            PADOUT => \N__7445\,
            PADIN => \N__7444\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2784\,
            DIN0 => \D_LL_AMIGA_in_6\,
            DOUT0 => \N__6647\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7437\,
            DIN => \N__7436\,
            DOUT => \N__7435\,
            PACKAGEPIN => D_UU_AMIGA(6)
        );

    \D_UU_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7437\,
            PADOUT => \N__7436\,
            PADIN => \N__7435\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2837\,
            DIN0 => \D_UU_AMIGA_in_6\,
            DOUT0 => \N__3050\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7428\,
            DIN => \N__7427\,
            DOUT => \N__7426\,
            PACKAGEPIN => D_UM_AMIGA(1)
        );

    \D_UM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7428\,
            PADOUT => \N__7427\,
            PADIN => \N__7426\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2711\,
            DIN0 => \D_UM_AMIGA_in_1\,
            DOUT0 => \N__2858\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7419\,
            DIN => \N__7418\,
            DOUT => \N__7417\,
            PACKAGEPIN => D_UU_040(5)
        );

    \D_UU_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7419\,
            PADOUT => \N__7418\,
            PADIN => \N__7417\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3934\,
            DIN0 => \D_UU_040_in_5\,
            DOUT0 => \N__5729\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7410\,
            DIN => \N__7409\,
            DOUT => \N__7408\,
            PACKAGEPIN => \CLKRAMA_wire\
        );

    \CLKRAMA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7410\,
            PADOUT => \N__7409\,
            PADIN => \N__7408\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6935\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7401\,
            DIN => \N__7400\,
            DOUT => \N__7399\,
            PACKAGEPIN => D_UM_040(2)
        );

    \D_UM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7401\,
            PADOUT => \N__7400\,
            PADIN => \N__7399\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3833\,
            DIN0 => \D_UM_040_in_2\,
            DOUT0 => \N__4814\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7392\,
            DIN => \N__7391\,
            DOUT => \N__7390\,
            PACKAGEPIN => D_LL_040(2)
        );

    \D_LL_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7392\,
            PADOUT => \N__7391\,
            PADIN => \N__7390\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4007\,
            DIN0 => \D_LL_040_in_2\,
            DOUT0 => \N__2243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7383\,
            DIN => \N__7382\,
            DOUT => \N__7381\,
            PACKAGEPIN => \TCI_CPUn_wire\
        );

    \TCI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7383\,
            PADOUT => \N__7382\,
            PADIN => \N__7381\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7023\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7374\,
            DIN => \N__7373\,
            DOUT => \N__7372\,
            PACKAGEPIN => \CLKRAMB_wire\
        );

    \CLKRAMB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7374\,
            PADOUT => \N__7373\,
            PADIN => \N__7372\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6928\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7365\,
            DIN => \N__7364\,
            DOUT => \N__7363\,
            PACKAGEPIN => D_LL_AMIGA(2)
        );

    \D_LL_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7365\,
            PADOUT => \N__7364\,
            PADIN => \N__7363\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2839\,
            DIN0 => \D_LL_AMIGA_in_2\,
            DOUT0 => \N__4877\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7356\,
            DIN => \N__7355\,
            DOUT => \N__7354\,
            PACKAGEPIN => D_UM_AMIGA(4)
        );

    \D_UM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7356\,
            PADOUT => \N__7355\,
            PADIN => \N__7354\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2781\,
            DIN0 => \D_UM_AMIGA_in_4\,
            DOUT0 => \N__5963\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7347\,
            DIN => \N__7346\,
            DOUT => \N__7345\,
            PACKAGEPIN => D_UU_AMIGA(2)
        );

    \D_UU_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7347\,
            PADOUT => \N__7346\,
            PADIN => \N__7345\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2833\,
            DIN0 => \D_UU_AMIGA_in_2\,
            DOUT0 => \N__4220\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7338\,
            DIN => \N__7337\,
            DOUT => \N__7336\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7338\,
            PADOUT => \N__7337\,
            PADIN => \N__7336\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7329\,
            DIN => \N__7328\,
            DOUT => \N__7327\,
            PACKAGEPIN => D_LM_AMIGA(6)
        );

    \D_LM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7329\,
            PADOUT => \N__7328\,
            PADIN => \N__7327\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2713\,
            DIN0 => \D_LM_AMIGA_in_6\,
            DOUT0 => \N__3110\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7320\,
            DIN => \N__7319\,
            DOUT => \N__7318\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7320\,
            PADOUT => \N__7319\,
            PADIN => \N__7318\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7311\,
            DIN => \N__7310\,
            DOUT => \N__7309\,
            PACKAGEPIN => D_LM_040(5)
        );

    \D_LM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7311\,
            PADOUT => \N__7310\,
            PADIN => \N__7309\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3835\,
            DIN0 => \D_LM_040_in_5\,
            DOUT0 => \N__2549\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7302\,
            DIN => \N__7301\,
            DOUT => \N__7300\,
            PACKAGEPIN => D_UM_040(6)
        );

    \D_UM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7302\,
            PADOUT => \N__7301\,
            PADIN => \N__7300\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3796\,
            DIN0 => \D_UM_040_in_6\,
            DOUT0 => \N__5318\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7293\,
            DIN => \N__7292\,
            DOUT => \N__7291\,
            PACKAGEPIN => \TAn_wire\
        );

    \TAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7293\,
            PADOUT => \N__7292\,
            PADIN => \N__7291\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4634\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMAn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7284\,
            DIN => \N__7283\,
            DOUT => \N__7282\,
            PACKAGEPIN => \DMAn_wire\
        );

    \DMAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7284\,
            PADOUT => \N__7283\,
            PADIN => \N__7282\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7031\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7275\,
            DIN => \N__7274\,
            DOUT => \N__7273\,
            PACKAGEPIN => D_LL_040(6)
        );

    \D_LL_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7275\,
            PADOUT => \N__7274\,
            PADIN => \N__7273\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4006\,
            DIN0 => \D_LL_040_in_6\,
            DOUT0 => \N__4109\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7266\,
            DIN => \N__7265\,
            DOUT => \N__7264\,
            PACKAGEPIN => D_LL_AMIGA(5)
        );

    \D_LL_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7266\,
            PADOUT => \N__7265\,
            PADIN => \N__7264\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2785\,
            DIN0 => \D_LL_AMIGA_in_5\,
            DOUT0 => \N__5849\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7257\,
            DIN => \N__7256\,
            DOUT => \N__7255\,
            PACKAGEPIN => D_UM_AMIGA(0)
        );

    \D_UM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7257\,
            PADOUT => \N__7256\,
            PADIN => \N__7255\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2673\,
            DIN0 => \D_UM_AMIGA_in_0\,
            DOUT0 => \N__6662\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7248\,
            DIN => \N__7247\,
            DOUT => \N__7246\,
            PACKAGEPIN => D_UU_040(2)
        );

    \D_UU_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7248\,
            PADOUT => \N__7247\,
            PADIN => \N__7246\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3969\,
            DIN0 => \D_UU_040_in_2\,
            DOUT0 => \N__5657\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7239\,
            DIN => \N__7238\,
            DOUT => \N__7237\,
            PACKAGEPIN => D_LM_AMIGA(2)
        );

    \D_LM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7239\,
            PADOUT => \N__7238\,
            PADIN => \N__7237\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2672\,
            DIN0 => \D_LM_AMIGA_in_2\,
            DOUT0 => \N__4256\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK80_CPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7230\,
            DIN => \N__7229\,
            DOUT => \N__7228\,
            PACKAGEPIN => \CLK80_CPU_wire\
        );

    \CLK80_CPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7230\,
            PADOUT => \N__7229\,
            PADIN => \N__7228\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6927\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7221\,
            DIN => \N__7220\,
            DOUT => \N__7219\,
            PACKAGEPIN => D_LL_040(3)
        );

    \D_LL_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7221\,
            PADOUT => \N__7220\,
            PADIN => \N__7219\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4027\,
            DIN0 => \D_LL_040_in_3\,
            DOUT0 => \N__3017\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7212\,
            DIN => \N__7211\,
            DOUT => \N__7210\,
            PACKAGEPIN => D_LM_040(1)
        );

    \D_LM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7212\,
            PADOUT => \N__7211\,
            PADIN => \N__7210\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3977\,
            DIN0 => \D_LM_040_in_1\,
            DOUT0 => \N__3668\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7203\,
            DIN => \N__7202\,
            DOUT => \N__7201\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7203\,
            PADOUT => \N__7202\,
            PADIN => \N__7201\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4064\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7194\,
            DIN => \N__7193\,
            DOUT => \N__7192\,
            PACKAGEPIN => D_UM_AMIGA(7)
        );

    \D_UM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7194\,
            PADOUT => \N__7193\,
            PADIN => \N__7192\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2780\,
            DIN0 => \D_UM_AMIGA_in_7\,
            DOUT0 => \N__3128\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7185\,
            DIN => \N__7184\,
            DOUT => \N__7183\,
            PACKAGEPIN => D_LM_AMIGA(7)
        );

    \D_LM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7185\,
            PADOUT => \N__7184\,
            PADIN => \N__7183\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2712\,
            DIN0 => \D_LM_AMIGA_in_7\,
            DOUT0 => \N__6794\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7176\,
            DIN => \N__7175\,
            DOUT => \N__7174\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7176\,
            PADOUT => \N__7175\,
            PADIN => \N__7174\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PORTSIZE_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7167\,
            DIN => \N__7166\,
            DOUT => \N__7165\,
            PACKAGEPIN => \A_AMIGA_wire\(0)
        );

    \A_AMIGA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7167\,
            PADOUT => \N__7166\,
            PADIN => \N__7165\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2273\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7158\,
            DIN => \N__7157\,
            DOUT => \N__7156\,
            PACKAGEPIN => D_LM_040(4)
        );

    \D_LM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7158\,
            PADOUT => \N__7157\,
            PADIN => \N__7156\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3880\,
            DIN0 => \D_LM_040_in_4\,
            DOUT0 => \N__2588\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7149\,
            DIN => \N__7148\,
            DOUT => \N__7147\,
            PACKAGEPIN => D_UM_040(7)
        );

    \D_UM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7149\,
            PADOUT => \N__7148\,
            PADIN => \N__7147\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3888\,
            DIN0 => \D_UM_040_in_7\,
            DOUT0 => \N__4997\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7140\,
            DIN => \N__7139\,
            DOUT => \N__7138\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7140\,
            PADOUT => \N__7139\,
            PADIN => \N__7138\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7131\,
            DIN => \N__7130\,
            DOUT => \N__7129\,
            PACKAGEPIN => D_UU_AMIGA(1)
        );

    \D_UU_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7131\,
            PADOUT => \N__7130\,
            PADIN => \N__7129\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2778\,
            DIN0 => \D_UU_AMIGA_in_1\,
            DOUT0 => \N__3509\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7122\,
            DIN => \N__7121\,
            DOUT => \N__7120\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7122\,
            PADOUT => \N__7121\,
            PADIN => \N__7120\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5544\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7113\,
            DIN => \N__7112\,
            DOUT => \N__7111\,
            PACKAGEPIN => D_UM_040(0)
        );

    \D_UM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7113\,
            PADOUT => \N__7112\,
            PADIN => \N__7111\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3834\,
            DIN0 => \D_UM_040_in_0\,
            DOUT0 => \N__2996\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7104\,
            DIN => \N__7103\,
            DOUT => \N__7102\,
            PACKAGEPIN => D_LL_AMIGA(0)
        );

    \D_LL_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7104\,
            PADOUT => \N__7103\,
            PADIN => \N__7102\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2840\,
            DIN0 => \D_LL_AMIGA_in_0\,
            DOUT0 => \N__6707\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7095\,
            DIN => \N__7094\,
            DOUT => \N__7093\,
            PACKAGEPIN => D_UU_AMIGA(4)
        );

    \D_UU_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7095\,
            PADOUT => \N__7094\,
            PADIN => \N__7093\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2832\,
            DIN0 => \D_UU_AMIGA_in_4\,
            DOUT0 => \N__6056\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7086\,
            DIN => \N__7085\,
            DOUT => \N__7084\,
            PACKAGEPIN => D_UU_040(7)
        );

    \D_UU_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7086\,
            PADOUT => \N__7085\,
            PADIN => \N__7084\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3935\,
            DIN0 => \D_UU_040_in_7\,
            DOUT0 => \N__3305\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7077\,
            DIN => \N__7076\,
            DOUT => \N__7075\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7077\,
            PADOUT => \N__7076\,
            PADIN => \N__7075\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7068\,
            DIN => \N__7067\,
            DOUT => \N__7066\,
            PACKAGEPIN => D_LL_040(0)
        );

    \D_LL_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7068\,
            PADOUT => \N__7067\,
            PADIN => \N__7066\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4028\,
            DIN0 => \D_LL_040_in_0\,
            DOUT0 => \N__2393\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7059\,
            DIN => \N__7058\,
            DOUT => \N__7057\,
            PACKAGEPIN => D_UM_AMIGA(2)
        );

    \D_UM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7059\,
            PADOUT => \N__7058\,
            PADIN => \N__7057\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2675\,
            DIN0 => \D_UM_AMIGA_in_2\,
            DOUT0 => \N__4835\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7050\,
            DIN => \N__7049\,
            DOUT => \N__7048\,
            PACKAGEPIN => D_UU_040(0)
        );

    \D_UU_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7050\,
            PADOUT => \N__7049\,
            PADIN => \N__7048\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3871\,
            DIN0 => \D_UU_040_in_0\,
            DOUT0 => \N__4148\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1804\ : IoInMux
    port map (
            O => \N__7031\,
            I => \N__7027\
        );

    \I__1803\ : IoInMux
    port map (
            O => \N__7030\,
            I => \N__7024\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__7027\,
            I => \N__7020\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__7024\,
            I => \N__7017\
        );

    \I__1800\ : IoInMux
    port map (
            O => \N__7023\,
            I => \N__7014\
        );

    \I__1799\ : Span4Mux_s3_v
    port map (
            O => \N__7020\,
            I => \N__7011\
        );

    \I__1798\ : IoSpan4Mux
    port map (
            O => \N__7017\,
            I => \N__7008\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__7014\,
            I => \N__7005\
        );

    \I__1796\ : Span4Mux_h
    port map (
            O => \N__7011\,
            I => \N__7002\
        );

    \I__1795\ : Span4Mux_s1_v
    port map (
            O => \N__7008\,
            I => \N__6999\
        );

    \I__1794\ : Span4Mux_s2_h
    port map (
            O => \N__7005\,
            I => \N__6996\
        );

    \I__1793\ : Sp12to4
    port map (
            O => \N__7002\,
            I => \N__6993\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__6999\,
            I => \N__6990\
        );

    \I__1791\ : Span4Mux_h
    port map (
            O => \N__6996\,
            I => \N__6987\
        );

    \I__1790\ : Span12Mux_h
    port map (
            O => \N__6993\,
            I => \N__6984\
        );

    \I__1789\ : Span4Mux_v
    port map (
            O => \N__6990\,
            I => \N__6979\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__6987\,
            I => \N__6979\
        );

    \I__1787\ : Odrv12
    port map (
            O => \N__6984\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1786\ : Odrv4
    port map (
            O => \N__6979\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1785\ : InMux
    port map (
            O => \N__6974\,
            I => \N__6971\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__6971\,
            I => \N__6960\
        );

    \I__1783\ : ClkMux
    port map (
            O => \N__6970\,
            I => \N__6938\
        );

    \I__1782\ : ClkMux
    port map (
            O => \N__6969\,
            I => \N__6938\
        );

    \I__1781\ : ClkMux
    port map (
            O => \N__6968\,
            I => \N__6938\
        );

    \I__1780\ : ClkMux
    port map (
            O => \N__6967\,
            I => \N__6938\
        );

    \I__1779\ : ClkMux
    port map (
            O => \N__6966\,
            I => \N__6938\
        );

    \I__1778\ : ClkMux
    port map (
            O => \N__6965\,
            I => \N__6938\
        );

    \I__1777\ : ClkMux
    port map (
            O => \N__6964\,
            I => \N__6938\
        );

    \I__1776\ : ClkMux
    port map (
            O => \N__6963\,
            I => \N__6938\
        );

    \I__1775\ : Glb2LocalMux
    port map (
            O => \N__6960\,
            I => \N__6938\
        );

    \I__1774\ : ClkMux
    port map (
            O => \N__6959\,
            I => \N__6938\
        );

    \I__1773\ : GlobalMux
    port map (
            O => \N__6938\,
            I => \CLK80\
        );

    \I__1772\ : IoInMux
    port map (
            O => \N__6935\,
            I => \N__6932\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__6932\,
            I => \N__6929\
        );

    \I__1770\ : IoSpan4Mux
    port map (
            O => \N__6929\,
            I => \N__6924\
        );

    \I__1769\ : IoInMux
    port map (
            O => \N__6928\,
            I => \N__6921\
        );

    \I__1768\ : IoInMux
    port map (
            O => \N__6927\,
            I => \N__6918\
        );

    \I__1767\ : IoSpan4Mux
    port map (
            O => \N__6924\,
            I => \N__6915\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__6921\,
            I => \N__6912\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__6918\,
            I => \N__6909\
        );

    \I__1764\ : Span4Mux_s3_v
    port map (
            O => \N__6915\,
            I => \N__6904\
        );

    \I__1763\ : Span4Mux_s3_v
    port map (
            O => \N__6912\,
            I => \N__6904\
        );

    \I__1762\ : IoSpan4Mux
    port map (
            O => \N__6909\,
            I => \N__6901\
        );

    \I__1761\ : Span4Mux_v
    port map (
            O => \N__6904\,
            I => \N__6898\
        );

    \I__1760\ : Span4Mux_s3_h
    port map (
            O => \N__6901\,
            I => \N__6895\
        );

    \I__1759\ : Span4Mux_v
    port map (
            O => \N__6898\,
            I => \N__6892\
        );

    \I__1758\ : Span4Mux_h
    port map (
            O => \N__6895\,
            I => \N__6889\
        );

    \I__1757\ : Span4Mux_v
    port map (
            O => \N__6892\,
            I => \N__6886\
        );

    \I__1756\ : Sp12to4
    port map (
            O => \N__6889\,
            I => \N__6883\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__6886\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1754\ : Odrv12
    port map (
            O => \N__6883\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1753\ : IoInMux
    port map (
            O => \N__6878\,
            I => \N__6875\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__6875\,
            I => \N__6872\
        );

    \I__1751\ : IoSpan4Mux
    port map (
            O => \N__6872\,
            I => \N__6868\
        );

    \I__1750\ : InMux
    port map (
            O => \N__6871\,
            I => \N__6865\
        );

    \I__1749\ : Span4Mux_s2_h
    port map (
            O => \N__6868\,
            I => \N__6862\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__6865\,
            I => \N__6859\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__6862\,
            I => \N__6856\
        );

    \I__1746\ : Span4Mux_v
    port map (
            O => \N__6859\,
            I => \N__6853\
        );

    \I__1745\ : Sp12to4
    port map (
            O => \N__6856\,
            I => \N__6850\
        );

    \I__1744\ : Sp12to4
    port map (
            O => \N__6853\,
            I => \N__6847\
        );

    \I__1743\ : Span12Mux_s9_h
    port map (
            O => \N__6850\,
            I => \N__6844\
        );

    \I__1742\ : Span12Mux_h
    port map (
            O => \N__6847\,
            I => \N__6841\
        );

    \I__1741\ : Span12Mux_h
    port map (
            O => \N__6844\,
            I => \N__6838\
        );

    \I__1740\ : Span12Mux_v
    port map (
            O => \N__6841\,
            I => \N__6835\
        );

    \I__1739\ : Odrv12
    port map (
            O => \N__6838\,
            I => \D_LM_040_in_5\
        );

    \I__1738\ : Odrv12
    port map (
            O => \N__6835\,
            I => \D_LM_040_in_5\
        );

    \I__1737\ : InMux
    port map (
            O => \N__6830\,
            I => \N__6827\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__6827\,
            I => \N__6824\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__6824\,
            I => \N__6821\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__6821\,
            I => \N__6818\
        );

    \I__1733\ : Sp12to4
    port map (
            O => \N__6818\,
            I => \N__6815\
        );

    \I__1732\ : Span12Mux_h
    port map (
            O => \N__6815\,
            I => \N__6812\
        );

    \I__1731\ : Odrv12
    port map (
            O => \N__6812\,
            I => \D_UU_040_in_5\
        );

    \I__1730\ : IoInMux
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__6806\,
            I => \N__6803\
        );

    \I__1728\ : Span12Mux_s3_h
    port map (
            O => \N__6803\,
            I => \N__6800\
        );

    \I__1727\ : Span12Mux_h
    port map (
            O => \N__6800\,
            I => \N__6797\
        );

    \I__1726\ : Odrv12
    port map (
            O => \N__6797\,
            I => \un1_D_UU_040_5\
        );

    \I__1725\ : IoInMux
    port map (
            O => \N__6794\,
            I => \N__6791\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__6791\,
            I => \N__6788\
        );

    \I__1723\ : Span4Mux_s1_h
    port map (
            O => \N__6788\,
            I => \N__6784\
        );

    \I__1722\ : InMux
    port map (
            O => \N__6787\,
            I => \N__6781\
        );

    \I__1721\ : Sp12to4
    port map (
            O => \N__6784\,
            I => \N__6778\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__6781\,
            I => \N__6775\
        );

    \I__1719\ : Span12Mux_s9_v
    port map (
            O => \N__6778\,
            I => \N__6772\
        );

    \I__1718\ : Span4Mux_v
    port map (
            O => \N__6775\,
            I => \N__6769\
        );

    \I__1717\ : Span12Mux_h
    port map (
            O => \N__6772\,
            I => \N__6766\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__6769\,
            I => \N__6763\
        );

    \I__1715\ : Span12Mux_h
    port map (
            O => \N__6766\,
            I => \N__6760\
        );

    \I__1714\ : Sp12to4
    port map (
            O => \N__6763\,
            I => \N__6757\
        );

    \I__1713\ : Odrv12
    port map (
            O => \N__6760\,
            I => \D_LM_040_in_7\
        );

    \I__1712\ : Odrv12
    port map (
            O => \N__6757\,
            I => \D_LM_040_in_7\
        );

    \I__1711\ : InMux
    port map (
            O => \N__6752\,
            I => \N__6749\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__6749\,
            I => \N__6746\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__6746\,
            I => \N__6743\
        );

    \I__1708\ : Sp12to4
    port map (
            O => \N__6743\,
            I => \N__6740\
        );

    \I__1707\ : Span12Mux_h
    port map (
            O => \N__6740\,
            I => \N__6737\
        );

    \I__1706\ : Odrv12
    port map (
            O => \N__6737\,
            I => \D_UU_040_in_7\
        );

    \I__1705\ : IoInMux
    port map (
            O => \N__6734\,
            I => \N__6731\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__6731\,
            I => \N__6728\
        );

    \I__1703\ : Span12Mux_s11_v
    port map (
            O => \N__6728\,
            I => \N__6725\
        );

    \I__1702\ : Span12Mux_h
    port map (
            O => \N__6725\,
            I => \N__6722\
        );

    \I__1701\ : Odrv12
    port map (
            O => \N__6722\,
            I => \un1_D_UU_040_7\
        );

    \I__1700\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6716\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__6716\,
            I => \N__6713\
        );

    \I__1698\ : Span12Mux_h
    port map (
            O => \N__6713\,
            I => \N__6710\
        );

    \I__1697\ : Odrv12
    port map (
            O => \N__6710\,
            I => \D_UM_040_in_0\
        );

    \I__1696\ : IoInMux
    port map (
            O => \N__6707\,
            I => \N__6704\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__6704\,
            I => \N__6700\
        );

    \I__1694\ : InMux
    port map (
            O => \N__6703\,
            I => \N__6697\
        );

    \I__1693\ : IoSpan4Mux
    port map (
            O => \N__6700\,
            I => \N__6694\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__6697\,
            I => \N__6691\
        );

    \I__1691\ : Span4Mux_s2_h
    port map (
            O => \N__6694\,
            I => \N__6688\
        );

    \I__1690\ : Span4Mux_v
    port map (
            O => \N__6691\,
            I => \N__6685\
        );

    \I__1689\ : Sp12to4
    port map (
            O => \N__6688\,
            I => \N__6682\
        );

    \I__1688\ : Sp12to4
    port map (
            O => \N__6685\,
            I => \N__6679\
        );

    \I__1687\ : Span12Mux_h
    port map (
            O => \N__6682\,
            I => \N__6676\
        );

    \I__1686\ : Span12Mux_v
    port map (
            O => \N__6679\,
            I => \N__6673\
        );

    \I__1685\ : Span12Mux_h
    port map (
            O => \N__6676\,
            I => \N__6670\
        );

    \I__1684\ : Span12Mux_h
    port map (
            O => \N__6673\,
            I => \N__6667\
        );

    \I__1683\ : Odrv12
    port map (
            O => \N__6670\,
            I => \D_LL_040_in_0\
        );

    \I__1682\ : Odrv12
    port map (
            O => \N__6667\,
            I => \D_LL_040_in_0\
        );

    \I__1681\ : IoInMux
    port map (
            O => \N__6662\,
            I => \N__6659\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__6659\,
            I => \N__6656\
        );

    \I__1679\ : Span12Mux_s4_h
    port map (
            O => \N__6656\,
            I => \N__6653\
        );

    \I__1678\ : Span12Mux_h
    port map (
            O => \N__6653\,
            I => \N__6650\
        );

    \I__1677\ : Odrv12
    port map (
            O => \N__6650\,
            I => \un1_D_UM_040_0\
        );

    \I__1676\ : IoInMux
    port map (
            O => \N__6647\,
            I => \N__6644\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__6644\,
            I => \N__6641\
        );

    \I__1674\ : IoSpan4Mux
    port map (
            O => \N__6641\,
            I => \N__6637\
        );

    \I__1673\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6634\
        );

    \I__1672\ : IoSpan4Mux
    port map (
            O => \N__6637\,
            I => \N__6631\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__6634\,
            I => \N__6628\
        );

    \I__1670\ : Span4Mux_s2_h
    port map (
            O => \N__6631\,
            I => \N__6625\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__6628\,
            I => \N__6622\
        );

    \I__1668\ : Sp12to4
    port map (
            O => \N__6625\,
            I => \N__6619\
        );

    \I__1667\ : Sp12to4
    port map (
            O => \N__6622\,
            I => \N__6616\
        );

    \I__1666\ : Span12Mux_h
    port map (
            O => \N__6619\,
            I => \N__6613\
        );

    \I__1665\ : Span12Mux_v
    port map (
            O => \N__6616\,
            I => \N__6610\
        );

    \I__1664\ : Span12Mux_h
    port map (
            O => \N__6613\,
            I => \N__6607\
        );

    \I__1663\ : Span12Mux_h
    port map (
            O => \N__6610\,
            I => \N__6604\
        );

    \I__1662\ : Odrv12
    port map (
            O => \N__6607\,
            I => \D_LL_040_in_6\
        );

    \I__1661\ : Odrv12
    port map (
            O => \N__6604\,
            I => \D_LL_040_in_6\
        );

    \I__1660\ : InMux
    port map (
            O => \N__6599\,
            I => \N__6596\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__6596\,
            I => \N__6593\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__6593\,
            I => \N__6590\
        );

    \I__1657\ : Sp12to4
    port map (
            O => \N__6590\,
            I => \N__6587\
        );

    \I__1656\ : Span12Mux_h
    port map (
            O => \N__6587\,
            I => \N__6584\
        );

    \I__1655\ : Odrv12
    port map (
            O => \N__6584\,
            I => \D_UM_040_in_6\
        );

    \I__1654\ : IoInMux
    port map (
            O => \N__6581\,
            I => \N__6578\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__6578\,
            I => \N__6575\
        );

    \I__1652\ : Span12Mux_s6_h
    port map (
            O => \N__6575\,
            I => \N__6572\
        );

    \I__1651\ : Span12Mux_v
    port map (
            O => \N__6572\,
            I => \N__6569\
        );

    \I__1650\ : Odrv12
    port map (
            O => \N__6569\,
            I => \un1_D_UM_040_6\
        );

    \I__1649\ : InMux
    port map (
            O => \N__6566\,
            I => \N__6562\
        );

    \I__1648\ : IoInMux
    port map (
            O => \N__6565\,
            I => \N__6559\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__6562\,
            I => \N__6556\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__6559\,
            I => \N__6553\
        );

    \I__1645\ : Span4Mux_v
    port map (
            O => \N__6556\,
            I => \N__6550\
        );

    \I__1644\ : Span4Mux_s3_h
    port map (
            O => \N__6553\,
            I => \N__6547\
        );

    \I__1643\ : Sp12to4
    port map (
            O => \N__6550\,
            I => \N__6544\
        );

    \I__1642\ : Sp12to4
    port map (
            O => \N__6547\,
            I => \N__6541\
        );

    \I__1641\ : Span12Mux_h
    port map (
            O => \N__6544\,
            I => \N__6538\
        );

    \I__1640\ : Span12Mux_v
    port map (
            O => \N__6541\,
            I => \N__6535\
        );

    \I__1639\ : Span12Mux_v
    port map (
            O => \N__6538\,
            I => \N__6532\
        );

    \I__1638\ : Span12Mux_h
    port map (
            O => \N__6535\,
            I => \N__6529\
        );

    \I__1637\ : Span12Mux_v
    port map (
            O => \N__6532\,
            I => \N__6524\
        );

    \I__1636\ : Span12Mux_h
    port map (
            O => \N__6529\,
            I => \N__6524\
        );

    \I__1635\ : Odrv12
    port map (
            O => \N__6524\,
            I => \D_LL_040_in_3\
        );

    \I__1634\ : InMux
    port map (
            O => \N__6521\,
            I => \N__6518\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__6518\,
            I => \N__6515\
        );

    \I__1632\ : Sp12to4
    port map (
            O => \N__6515\,
            I => \N__6512\
        );

    \I__1631\ : Span12Mux_v
    port map (
            O => \N__6512\,
            I => \N__6509\
        );

    \I__1630\ : Span12Mux_h
    port map (
            O => \N__6509\,
            I => \N__6506\
        );

    \I__1629\ : Odrv12
    port map (
            O => \N__6506\,
            I => \D_UM_040_in_3\
        );

    \I__1628\ : IoInMux
    port map (
            O => \N__6503\,
            I => \N__6500\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__6500\,
            I => \N__6497\
        );

    \I__1626\ : IoSpan4Mux
    port map (
            O => \N__6497\,
            I => \N__6494\
        );

    \I__1625\ : Span4Mux_s3_h
    port map (
            O => \N__6494\,
            I => \N__6491\
        );

    \I__1624\ : Sp12to4
    port map (
            O => \N__6491\,
            I => \N__6488\
        );

    \I__1623\ : Span12Mux_h
    port map (
            O => \N__6488\,
            I => \N__6485\
        );

    \I__1622\ : Odrv12
    port map (
            O => \N__6485\,
            I => \un1_D_UM_040_3\
        );

    \I__1621\ : InMux
    port map (
            O => \N__6482\,
            I => \N__6479\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__6479\,
            I => \N__6476\
        );

    \I__1619\ : Span4Mux_v
    port map (
            O => \N__6476\,
            I => \N__6473\
        );

    \I__1618\ : Sp12to4
    port map (
            O => \N__6473\,
            I => \N__6470\
        );

    \I__1617\ : Span12Mux_h
    port map (
            O => \N__6470\,
            I => \N__6467\
        );

    \I__1616\ : Odrv12
    port map (
            O => \N__6467\,
            I => \SIZ_c_0\
        );

    \I__1615\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6461\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__6461\,
            I => \N__6458\
        );

    \I__1613\ : Span4Mux_v
    port map (
            O => \N__6458\,
            I => \N__6455\
        );

    \I__1612\ : Sp12to4
    port map (
            O => \N__6455\,
            I => \N__6452\
        );

    \I__1611\ : Span12Mux_h
    port map (
            O => \N__6452\,
            I => \N__6449\
        );

    \I__1610\ : Odrv12
    port map (
            O => \N__6449\,
            I => \SIZ_c_1\
        );

    \I__1609\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6443\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__6443\,
            I => \N__6439\
        );

    \I__1607\ : InMux
    port map (
            O => \N__6442\,
            I => \N__6436\
        );

    \I__1606\ : Span4Mux_v
    port map (
            O => \N__6439\,
            I => \N__6433\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__6436\,
            I => \N__6430\
        );

    \I__1604\ : Span4Mux_v
    port map (
            O => \N__6433\,
            I => \N__6427\
        );

    \I__1603\ : Span4Mux_v
    port map (
            O => \N__6430\,
            I => \N__6424\
        );

    \I__1602\ : Sp12to4
    port map (
            O => \N__6427\,
            I => \N__6419\
        );

    \I__1601\ : Sp12to4
    port map (
            O => \N__6424\,
            I => \N__6419\
        );

    \I__1600\ : Span12Mux_h
    port map (
            O => \N__6419\,
            I => \N__6416\
        );

    \I__1599\ : Span12Mux_v
    port map (
            O => \N__6416\,
            I => \N__6413\
        );

    \I__1598\ : Odrv12
    port map (
            O => \N__6413\,
            I => \PORTSIZE_c\
        );

    \I__1597\ : InMux
    port map (
            O => \N__6410\,
            I => \N__6407\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__6407\,
            I => \N__6404\
        );

    \I__1595\ : Span4Mux_h
    port map (
            O => \N__6404\,
            I => \N__6400\
        );

    \I__1594\ : InMux
    port map (
            O => \N__6403\,
            I => \N__6397\
        );

    \I__1593\ : Sp12to4
    port map (
            O => \N__6400\,
            I => \N__6392\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__6397\,
            I => \N__6392\
        );

    \I__1591\ : Span12Mux_v
    port map (
            O => \N__6392\,
            I => \N__6389\
        );

    \I__1590\ : Odrv12
    port map (
            O => \N__6389\,
            I => \U111_CYCLE_SM.LW_TRANS_0\
        );

    \I__1589\ : InMux
    port map (
            O => \N__6386\,
            I => \N__6383\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__6383\,
            I => \N__6380\
        );

    \I__1587\ : Span4Mux_v
    port map (
            O => \N__6380\,
            I => \N__6377\
        );

    \I__1586\ : Span4Mux_h
    port map (
            O => \N__6377\,
            I => \N__6374\
        );

    \I__1585\ : Span4Mux_h
    port map (
            O => \N__6374\,
            I => \N__6371\
        );

    \I__1584\ : Odrv4
    port map (
            O => \N__6371\,
            I => \D_UU_040_in_4\
        );

    \I__1583\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6358\
        );

    \I__1582\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6355\
        );

    \I__1581\ : InMux
    port map (
            O => \N__6366\,
            I => \N__6350\
        );

    \I__1580\ : InMux
    port map (
            O => \N__6365\,
            I => \N__6350\
        );

    \I__1579\ : InMux
    port map (
            O => \N__6364\,
            I => \N__6347\
        );

    \I__1578\ : InMux
    port map (
            O => \N__6363\,
            I => \N__6342\
        );

    \I__1577\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6342\
        );

    \I__1576\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6338\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__6358\,
            I => \N__6335\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__6355\,
            I => \N__6330\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__6350\,
            I => \N__6330\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__6347\,
            I => \N__6321\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__6342\,
            I => \N__6321\
        );

    \I__1570\ : InMux
    port map (
            O => \N__6341\,
            I => \N__6318\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__6338\,
            I => \N__6311\
        );

    \I__1568\ : Span4Mux_v
    port map (
            O => \N__6335\,
            I => \N__6306\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__6330\,
            I => \N__6306\
        );

    \I__1566\ : InMux
    port map (
            O => \N__6329\,
            I => \N__6303\
        );

    \I__1565\ : InMux
    port map (
            O => \N__6328\,
            I => \N__6300\
        );

    \I__1564\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6294\
        );

    \I__1563\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6291\
        );

    \I__1562\ : Span4Mux_v
    port map (
            O => \N__6321\,
            I => \N__6284\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__6318\,
            I => \N__6284\
        );

    \I__1560\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6281\
        );

    \I__1559\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6276\
        );

    \I__1558\ : InMux
    port map (
            O => \N__6315\,
            I => \N__6273\
        );

    \I__1557\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6270\
        );

    \I__1556\ : Span4Mux_v
    port map (
            O => \N__6311\,
            I => \N__6262\
        );

    \I__1555\ : Span4Mux_h
    port map (
            O => \N__6306\,
            I => \N__6262\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__6303\,
            I => \N__6262\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__6300\,
            I => \N__6259\
        );

    \I__1552\ : InMux
    port map (
            O => \N__6299\,
            I => \N__6256\
        );

    \I__1551\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6253\
        );

    \I__1550\ : InMux
    port map (
            O => \N__6297\,
            I => \N__6250\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__6294\,
            I => \N__6244\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__6291\,
            I => \N__6241\
        );

    \I__1547\ : InMux
    port map (
            O => \N__6290\,
            I => \N__6238\
        );

    \I__1546\ : InMux
    port map (
            O => \N__6289\,
            I => \N__6235\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__6284\,
            I => \N__6229\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__6281\,
            I => \N__6226\
        );

    \I__1543\ : InMux
    port map (
            O => \N__6280\,
            I => \N__6223\
        );

    \I__1542\ : InMux
    port map (
            O => \N__6279\,
            I => \N__6220\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__6276\,
            I => \N__6217\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__6273\,
            I => \N__6214\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__6270\,
            I => \N__6211\
        );

    \I__1538\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6208\
        );

    \I__1537\ : Span4Mux_v
    port map (
            O => \N__6262\,
            I => \N__6197\
        );

    \I__1536\ : Span4Mux_h
    port map (
            O => \N__6259\,
            I => \N__6197\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__6256\,
            I => \N__6197\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__6253\,
            I => \N__6197\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__6250\,
            I => \N__6197\
        );

    \I__1532\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6194\
        );

    \I__1531\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6191\
        );

    \I__1530\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6188\
        );

    \I__1529\ : Span4Mux_h
    port map (
            O => \N__6244\,
            I => \N__6179\
        );

    \I__1528\ : Span4Mux_v
    port map (
            O => \N__6241\,
            I => \N__6179\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__6238\,
            I => \N__6179\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__6235\,
            I => \N__6179\
        );

    \I__1525\ : InMux
    port map (
            O => \N__6234\,
            I => \N__6174\
        );

    \I__1524\ : InMux
    port map (
            O => \N__6233\,
            I => \N__6174\
        );

    \I__1523\ : InMux
    port map (
            O => \N__6232\,
            I => \N__6171\
        );

    \I__1522\ : Span4Mux_h
    port map (
            O => \N__6229\,
            I => \N__6165\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__6226\,
            I => \N__6165\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__6223\,
            I => \N__6160\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__6220\,
            I => \N__6160\
        );

    \I__1518\ : Span4Mux_v
    port map (
            O => \N__6217\,
            I => \N__6157\
        );

    \I__1517\ : Span4Mux_v
    port map (
            O => \N__6214\,
            I => \N__6152\
        );

    \I__1516\ : Span4Mux_v
    port map (
            O => \N__6211\,
            I => \N__6152\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__6208\,
            I => \N__6149\
        );

    \I__1514\ : Span4Mux_v
    port map (
            O => \N__6197\,
            I => \N__6144\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__6194\,
            I => \N__6144\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__6191\,
            I => \N__6139\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__6188\,
            I => \N__6139\
        );

    \I__1510\ : Span4Mux_h
    port map (
            O => \N__6179\,
            I => \N__6134\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6134\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__6171\,
            I => \N__6131\
        );

    \I__1507\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6128\
        );

    \I__1506\ : Span4Mux_v
    port map (
            O => \N__6165\,
            I => \N__6125\
        );

    \I__1505\ : Span12Mux_v
    port map (
            O => \N__6160\,
            I => \N__6122\
        );

    \I__1504\ : Span4Mux_h
    port map (
            O => \N__6157\,
            I => \N__6115\
        );

    \I__1503\ : Span4Mux_h
    port map (
            O => \N__6152\,
            I => \N__6115\
        );

    \I__1502\ : Span4Mux_v
    port map (
            O => \N__6149\,
            I => \N__6115\
        );

    \I__1501\ : Span4Mux_v
    port map (
            O => \N__6144\,
            I => \N__6104\
        );

    \I__1500\ : Span4Mux_v
    port map (
            O => \N__6139\,
            I => \N__6104\
        );

    \I__1499\ : Span4Mux_v
    port map (
            O => \N__6134\,
            I => \N__6104\
        );

    \I__1498\ : Span4Mux_h
    port map (
            O => \N__6131\,
            I => \N__6104\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__6128\,
            I => \N__6104\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__6125\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1495\ : Odrv12
    port map (
            O => \N__6122\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1494\ : Odrv4
    port map (
            O => \N__6115\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__6104\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__1492\ : IoInMux
    port map (
            O => \N__6095\,
            I => \N__6092\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__6092\,
            I => \N__6089\
        );

    \I__1490\ : Span4Mux_s1_h
    port map (
            O => \N__6089\,
            I => \N__6086\
        );

    \I__1489\ : Sp12to4
    port map (
            O => \N__6086\,
            I => \N__6082\
        );

    \I__1488\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6079\
        );

    \I__1487\ : Span12Mux_v
    port map (
            O => \N__6082\,
            I => \N__6076\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__6079\,
            I => \N__6073\
        );

    \I__1485\ : Span12Mux_h
    port map (
            O => \N__6076\,
            I => \N__6070\
        );

    \I__1484\ : Span12Mux_h
    port map (
            O => \N__6073\,
            I => \N__6067\
        );

    \I__1483\ : Span12Mux_h
    port map (
            O => \N__6070\,
            I => \N__6064\
        );

    \I__1482\ : Span12Mux_v
    port map (
            O => \N__6067\,
            I => \N__6061\
        );

    \I__1481\ : Odrv12
    port map (
            O => \N__6064\,
            I => \D_LM_040_in_4\
        );

    \I__1480\ : Odrv12
    port map (
            O => \N__6061\,
            I => \D_LM_040_in_4\
        );

    \I__1479\ : IoInMux
    port map (
            O => \N__6056\,
            I => \N__6053\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__6053\,
            I => \N__6050\
        );

    \I__1477\ : IoSpan4Mux
    port map (
            O => \N__6050\,
            I => \N__6047\
        );

    \I__1476\ : IoSpan4Mux
    port map (
            O => \N__6047\,
            I => \N__6044\
        );

    \I__1475\ : Span4Mux_s2_v
    port map (
            O => \N__6044\,
            I => \N__6041\
        );

    \I__1474\ : Span4Mux_v
    port map (
            O => \N__6041\,
            I => \N__6038\
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__6038\,
            I => \un1_D_UU_040_4\
        );

    \I__1472\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6032\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__6032\,
            I => \N__6028\
        );

    \I__1470\ : IoInMux
    port map (
            O => \N__6031\,
            I => \N__6025\
        );

    \I__1469\ : Span4Mux_v
    port map (
            O => \N__6028\,
            I => \N__6022\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__6025\,
            I => \N__6019\
        );

    \I__1467\ : Span4Mux_h
    port map (
            O => \N__6022\,
            I => \N__6016\
        );

    \I__1466\ : Span4Mux_s2_h
    port map (
            O => \N__6019\,
            I => \N__6013\
        );

    \I__1465\ : Sp12to4
    port map (
            O => \N__6016\,
            I => \N__6010\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__6013\,
            I => \N__6007\
        );

    \I__1463\ : Span12Mux_h
    port map (
            O => \N__6010\,
            I => \N__6004\
        );

    \I__1462\ : Sp12to4
    port map (
            O => \N__6007\,
            I => \N__6001\
        );

    \I__1461\ : Span12Mux_v
    port map (
            O => \N__6004\,
            I => \N__5998\
        );

    \I__1460\ : Span12Mux_h
    port map (
            O => \N__6001\,
            I => \N__5995\
        );

    \I__1459\ : Span12Mux_v
    port map (
            O => \N__5998\,
            I => \N__5992\
        );

    \I__1458\ : Span12Mux_h
    port map (
            O => \N__5995\,
            I => \N__5989\
        );

    \I__1457\ : Odrv12
    port map (
            O => \N__5992\,
            I => \D_LL_040_in_4\
        );

    \I__1456\ : Odrv12
    port map (
            O => \N__5989\,
            I => \D_LL_040_in_4\
        );

    \I__1455\ : InMux
    port map (
            O => \N__5984\,
            I => \N__5981\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__5981\,
            I => \N__5978\
        );

    \I__1453\ : Span4Mux_v
    port map (
            O => \N__5978\,
            I => \N__5975\
        );

    \I__1452\ : Span4Mux_h
    port map (
            O => \N__5975\,
            I => \N__5972\
        );

    \I__1451\ : Sp12to4
    port map (
            O => \N__5972\,
            I => \N__5969\
        );

    \I__1450\ : Span12Mux_h
    port map (
            O => \N__5969\,
            I => \N__5966\
        );

    \I__1449\ : Odrv12
    port map (
            O => \N__5966\,
            I => \D_UM_040_in_4\
        );

    \I__1448\ : IoInMux
    port map (
            O => \N__5963\,
            I => \N__5960\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__5960\,
            I => \N__5957\
        );

    \I__1446\ : Span4Mux_s2_h
    port map (
            O => \N__5957\,
            I => \N__5954\
        );

    \I__1445\ : Span4Mux_h
    port map (
            O => \N__5954\,
            I => \N__5951\
        );

    \I__1444\ : Span4Mux_h
    port map (
            O => \N__5951\,
            I => \N__5948\
        );

    \I__1443\ : Span4Mux_h
    port map (
            O => \N__5948\,
            I => \N__5945\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__5945\,
            I => \un1_D_UM_040_4\
        );

    \I__1441\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5939\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__5939\,
            I => \N__5936\
        );

    \I__1439\ : Odrv12
    port map (
            O => \N__5936\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__1438\ : InMux
    port map (
            O => \N__5933\,
            I => \N__5930\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__5930\,
            I => \N__5927\
        );

    \I__1436\ : Span4Mux_v
    port map (
            O => \N__5927\,
            I => \N__5922\
        );

    \I__1435\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5919\
        );

    \I__1434\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5916\
        );

    \I__1433\ : Sp12to4
    port map (
            O => \N__5922\,
            I => \N__5913\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__5919\,
            I => \N__5908\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__5916\,
            I => \N__5908\
        );

    \I__1430\ : Span12Mux_h
    port map (
            O => \N__5913\,
            I => \N__5905\
        );

    \I__1429\ : Span12Mux_v
    port map (
            O => \N__5908\,
            I => \N__5902\
        );

    \I__1428\ : Span12Mux_v
    port map (
            O => \N__5905\,
            I => \N__5897\
        );

    \I__1427\ : Span12Mux_h
    port map (
            O => \N__5902\,
            I => \N__5897\
        );

    \I__1426\ : Odrv12
    port map (
            O => \N__5897\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__1425\ : IoInMux
    port map (
            O => \N__5894\,
            I => \N__5891\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__5891\,
            I => \N__5888\
        );

    \I__1423\ : Span4Mux_s3_v
    port map (
            O => \N__5888\,
            I => \N__5885\
        );

    \I__1422\ : Span4Mux_h
    port map (
            O => \N__5885\,
            I => \N__5882\
        );

    \I__1421\ : Span4Mux_h
    port map (
            O => \N__5882\,
            I => \N__5879\
        );

    \I__1420\ : Span4Mux_h
    port map (
            O => \N__5879\,
            I => \N__5876\
        );

    \I__1419\ : Span4Mux_h
    port map (
            O => \N__5876\,
            I => \N__5873\
        );

    \I__1418\ : Odrv4
    port map (
            O => \N__5873\,
            I => \un1_D_UU_AMIGA_3\
        );

    \I__1417\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5867\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__5867\,
            I => \N__5864\
        );

    \I__1415\ : Span4Mux_v
    port map (
            O => \N__5864\,
            I => \N__5861\
        );

    \I__1414\ : Span4Mux_h
    port map (
            O => \N__5861\,
            I => \N__5858\
        );

    \I__1413\ : Sp12to4
    port map (
            O => \N__5858\,
            I => \N__5855\
        );

    \I__1412\ : Span12Mux_h
    port map (
            O => \N__5855\,
            I => \N__5852\
        );

    \I__1411\ : Odrv12
    port map (
            O => \N__5852\,
            I => \D_UM_040_in_5\
        );

    \I__1410\ : IoInMux
    port map (
            O => \N__5849\,
            I => \N__5846\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__5846\,
            I => \N__5842\
        );

    \I__1408\ : InMux
    port map (
            O => \N__5845\,
            I => \N__5839\
        );

    \I__1407\ : IoSpan4Mux
    port map (
            O => \N__5842\,
            I => \N__5836\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__5839\,
            I => \N__5833\
        );

    \I__1405\ : Span4Mux_s3_h
    port map (
            O => \N__5836\,
            I => \N__5830\
        );

    \I__1404\ : Sp12to4
    port map (
            O => \N__5833\,
            I => \N__5827\
        );

    \I__1403\ : Sp12to4
    port map (
            O => \N__5830\,
            I => \N__5824\
        );

    \I__1402\ : Span12Mux_v
    port map (
            O => \N__5827\,
            I => \N__5821\
        );

    \I__1401\ : Span12Mux_v
    port map (
            O => \N__5824\,
            I => \N__5818\
        );

    \I__1400\ : Span12Mux_v
    port map (
            O => \N__5821\,
            I => \N__5813\
        );

    \I__1399\ : Span12Mux_h
    port map (
            O => \N__5818\,
            I => \N__5813\
        );

    \I__1398\ : Span12Mux_h
    port map (
            O => \N__5813\,
            I => \N__5810\
        );

    \I__1397\ : Odrv12
    port map (
            O => \N__5810\,
            I => \D_LL_040_in_5\
        );

    \I__1396\ : IoInMux
    port map (
            O => \N__5807\,
            I => \N__5804\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__1394\ : IoSpan4Mux
    port map (
            O => \N__5801\,
            I => \N__5798\
        );

    \I__1393\ : IoSpan4Mux
    port map (
            O => \N__5798\,
            I => \N__5795\
        );

    \I__1392\ : Span4Mux_s2_v
    port map (
            O => \N__5795\,
            I => \N__5792\
        );

    \I__1391\ : Span4Mux_v
    port map (
            O => \N__5792\,
            I => \N__5789\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__5789\,
            I => \un1_D_UM_040_5\
        );

    \I__1389\ : InMux
    port map (
            O => \N__5786\,
            I => \N__5783\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__5783\,
            I => \N__5780\
        );

    \I__1387\ : Span4Mux_v
    port map (
            O => \N__5780\,
            I => \N__5777\
        );

    \I__1386\ : Odrv4
    port map (
            O => \N__5777\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__1385\ : InMux
    port map (
            O => \N__5774\,
            I => \N__5771\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__5771\,
            I => \N__5768\
        );

    \I__1383\ : Span4Mux_v
    port map (
            O => \N__5768\,
            I => \N__5764\
        );

    \I__1382\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5761\
        );

    \I__1381\ : Span4Mux_v
    port map (
            O => \N__5764\,
            I => \N__5756\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__5761\,
            I => \N__5756\
        );

    \I__1379\ : Span4Mux_h
    port map (
            O => \N__5756\,
            I => \N__5752\
        );

    \I__1378\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5749\
        );

    \I__1377\ : Span4Mux_v
    port map (
            O => \N__5752\,
            I => \N__5746\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__5749\,
            I => \N__5743\
        );

    \I__1375\ : Span4Mux_h
    port map (
            O => \N__5746\,
            I => \N__5740\
        );

    \I__1374\ : Span12Mux_v
    port map (
            O => \N__5743\,
            I => \N__5737\
        );

    \I__1373\ : Span4Mux_h
    port map (
            O => \N__5740\,
            I => \N__5734\
        );

    \I__1372\ : Odrv12
    port map (
            O => \N__5737\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1371\ : Odrv4
    port map (
            O => \N__5734\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1370\ : IoInMux
    port map (
            O => \N__5729\,
            I => \N__5726\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__5726\,
            I => \N__5723\
        );

    \I__1368\ : Span12Mux_s6_v
    port map (
            O => \N__5723\,
            I => \N__5720\
        );

    \I__1367\ : Span12Mux_h
    port map (
            O => \N__5720\,
            I => \N__5717\
        );

    \I__1366\ : Odrv12
    port map (
            O => \N__5717\,
            I => \un1_D_UU_AMIGA_5\
        );

    \I__1365\ : InMux
    port map (
            O => \N__5714\,
            I => \N__5711\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__5711\,
            I => \N__5708\
        );

    \I__1363\ : Odrv12
    port map (
            O => \N__5708\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__1362\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5702\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__5702\,
            I => \N__5698\
        );

    \I__1360\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5694\
        );

    \I__1359\ : Span4Mux_v
    port map (
            O => \N__5698\,
            I => \N__5691\
        );

    \I__1358\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5688\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__5694\,
            I => \N__5685\
        );

    \I__1356\ : Span4Mux_v
    port map (
            O => \N__5691\,
            I => \N__5680\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__5688\,
            I => \N__5680\
        );

    \I__1354\ : Span4Mux_v
    port map (
            O => \N__5685\,
            I => \N__5677\
        );

    \I__1353\ : Span4Mux_v
    port map (
            O => \N__5680\,
            I => \N__5674\
        );

    \I__1352\ : Span4Mux_h
    port map (
            O => \N__5677\,
            I => \N__5671\
        );

    \I__1351\ : Sp12to4
    port map (
            O => \N__5674\,
            I => \N__5668\
        );

    \I__1350\ : Sp12to4
    port map (
            O => \N__5671\,
            I => \N__5665\
        );

    \I__1349\ : Span12Mux_h
    port map (
            O => \N__5668\,
            I => \N__5662\
        );

    \I__1348\ : Odrv12
    port map (
            O => \N__5665\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__1347\ : Odrv12
    port map (
            O => \N__5662\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__1346\ : IoInMux
    port map (
            O => \N__5657\,
            I => \N__5654\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__5654\,
            I => \N__5651\
        );

    \I__1344\ : Span12Mux_s0_v
    port map (
            O => \N__5651\,
            I => \N__5648\
        );

    \I__1343\ : Span12Mux_h
    port map (
            O => \N__5648\,
            I => \N__5645\
        );

    \I__1342\ : Odrv12
    port map (
            O => \N__5645\,
            I => \un1_D_UU_AMIGA_2\
        );

    \I__1341\ : InMux
    port map (
            O => \N__5642\,
            I => \N__5639\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__1339\ : Span4Mux_v
    port map (
            O => \N__5636\,
            I => \N__5632\
        );

    \I__1338\ : InMux
    port map (
            O => \N__5635\,
            I => \N__5629\
        );

    \I__1337\ : Span4Mux_v
    port map (
            O => \N__5632\,
            I => \N__5624\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__5629\,
            I => \N__5624\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__5624\,
            I => \N__5620\
        );

    \I__1334\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5617\
        );

    \I__1333\ : Span4Mux_v
    port map (
            O => \N__5620\,
            I => \N__5612\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__5617\,
            I => \N__5612\
        );

    \I__1331\ : Span4Mux_v
    port map (
            O => \N__5612\,
            I => \N__5609\
        );

    \I__1330\ : Sp12to4
    port map (
            O => \N__5609\,
            I => \N__5606\
        );

    \I__1329\ : Span12Mux_h
    port map (
            O => \N__5606\,
            I => \N__5603\
        );

    \I__1328\ : Odrv12
    port map (
            O => \N__5603\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1327\ : InMux
    port map (
            O => \N__5600\,
            I => \N__5597\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__1325\ : Odrv12
    port map (
            O => \N__5594\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__1324\ : IoInMux
    port map (
            O => \N__5591\,
            I => \N__5588\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__5588\,
            I => \N__5585\
        );

    \I__1322\ : Span4Mux_s2_v
    port map (
            O => \N__5585\,
            I => \N__5582\
        );

    \I__1321\ : Span4Mux_h
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__1320\ : Span4Mux_v
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__1319\ : Sp12to4
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__1318\ : Odrv12
    port map (
            O => \N__5573\,
            I => \un1_D_UM_AMIGA_5\
        );

    \I__1317\ : InMux
    port map (
            O => \N__5570\,
            I => \N__5566\
        );

    \I__1316\ : InMux
    port map (
            O => \N__5569\,
            I => \N__5563\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__5566\,
            I => \N__5559\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__5563\,
            I => \N__5556\
        );

    \I__1313\ : ClkMux
    port map (
            O => \N__5562\,
            I => \N__5549\
        );

    \I__1312\ : Glb2LocalMux
    port map (
            O => \N__5559\,
            I => \N__5549\
        );

    \I__1311\ : Glb2LocalMux
    port map (
            O => \N__5556\,
            I => \N__5549\
        );

    \I__1310\ : GlobalMux
    port map (
            O => \N__5549\,
            I => \CLK40\
        );

    \I__1309\ : IoInMux
    port map (
            O => \N__5546\,
            I => \N__5541\
        );

    \I__1308\ : IoInMux
    port map (
            O => \N__5545\,
            I => \N__5538\
        );

    \I__1307\ : IoInMux
    port map (
            O => \N__5544\,
            I => \N__5535\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__5541\,
            I => \N__5532\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__5538\,
            I => \N__5529\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5535\,
            I => \N__5526\
        );

    \I__1303\ : Span12Mux_s5_v
    port map (
            O => \N__5532\,
            I => \N__5523\
        );

    \I__1302\ : Span12Mux_s10_h
    port map (
            O => \N__5529\,
            I => \N__5518\
        );

    \I__1301\ : Span12Mux_s9_h
    port map (
            O => \N__5526\,
            I => \N__5518\
        );

    \I__1300\ : Odrv12
    port map (
            O => \N__5523\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__1299\ : Odrv12
    port map (
            O => \N__5518\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5513\,
            I => \N__5507\
        );

    \I__1297\ : InMux
    port map (
            O => \N__5512\,
            I => \N__5507\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__5507\,
            I => \N__5497\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5506\,
            I => \N__5488\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5488\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5488\
        );

    \I__1292\ : InMux
    port map (
            O => \N__5503\,
            I => \N__5488\
        );

    \I__1291\ : InMux
    port map (
            O => \N__5502\,
            I => \N__5481\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5501\,
            I => \N__5478\
        );

    \I__1289\ : InMux
    port map (
            O => \N__5500\,
            I => \N__5473\
        );

    \I__1288\ : Span4Mux_v
    port map (
            O => \N__5497\,
            I => \N__5470\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5488\,
            I => \N__5467\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5487\,
            I => \N__5464\
        );

    \I__1285\ : InMux
    port map (
            O => \N__5486\,
            I => \N__5461\
        );

    \I__1284\ : InMux
    port map (
            O => \N__5485\,
            I => \N__5456\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5484\,
            I => \N__5456\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__5481\,
            I => \N__5451\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__5478\,
            I => \N__5451\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5477\,
            I => \N__5448\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5476\,
            I => \N__5445\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5473\,
            I => \N__5441\
        );

    \I__1277\ : Sp12to4
    port map (
            O => \N__5470\,
            I => \N__5437\
        );

    \I__1276\ : Span4Mux_v
    port map (
            O => \N__5467\,
            I => \N__5430\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5464\,
            I => \N__5430\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5461\,
            I => \N__5430\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__5456\,
            I => \N__5421\
        );

    \I__1272\ : Span4Mux_v
    port map (
            O => \N__5451\,
            I => \N__5421\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__5448\,
            I => \N__5421\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__5445\,
            I => \N__5421\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5418\
        );

    \I__1268\ : Span4Mux_v
    port map (
            O => \N__5441\,
            I => \N__5413\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5440\,
            I => \N__5410\
        );

    \I__1266\ : Span12Mux_h
    port map (
            O => \N__5437\,
            I => \N__5405\
        );

    \I__1265\ : Span4Mux_v
    port map (
            O => \N__5430\,
            I => \N__5402\
        );

    \I__1264\ : Span4Mux_v
    port map (
            O => \N__5421\,
            I => \N__5397\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5418\,
            I => \N__5397\
        );

    \I__1262\ : InMux
    port map (
            O => \N__5417\,
            I => \N__5394\
        );

    \I__1261\ : InMux
    port map (
            O => \N__5416\,
            I => \N__5391\
        );

    \I__1260\ : Span4Mux_v
    port map (
            O => \N__5413\,
            I => \N__5386\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__5410\,
            I => \N__5386\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5409\,
            I => \N__5381\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5381\
        );

    \I__1256\ : Odrv12
    port map (
            O => \N__5405\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__5402\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__5397\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__5394\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__5391\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1251\ : Odrv4
    port map (
            O => \N__5386\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5381\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5363\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__5357\,
            I => \N__5354\
        );

    \I__1245\ : Span4Mux_h
    port map (
            O => \N__5354\,
            I => \N__5350\
        );

    \I__1244\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5347\
        );

    \I__1243\ : Span4Mux_v
    port map (
            O => \N__5350\,
            I => \N__5343\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5347\,
            I => \N__5340\
        );

    \I__1241\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5337\
        );

    \I__1240\ : Span4Mux_h
    port map (
            O => \N__5343\,
            I => \N__5334\
        );

    \I__1239\ : Sp12to4
    port map (
            O => \N__5340\,
            I => \N__5329\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__5337\,
            I => \N__5329\
        );

    \I__1237\ : Sp12to4
    port map (
            O => \N__5334\,
            I => \N__5324\
        );

    \I__1236\ : Span12Mux_h
    port map (
            O => \N__5329\,
            I => \N__5324\
        );

    \I__1235\ : Span12Mux_v
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__1234\ : Odrv12
    port map (
            O => \N__5321\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__1233\ : IoInMux
    port map (
            O => \N__5318\,
            I => \N__5315\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__5315\,
            I => \N__5312\
        );

    \I__1231\ : Span12Mux_s4_h
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__1230\ : Span12Mux_h
    port map (
            O => \N__5309\,
            I => \N__5306\
        );

    \I__1229\ : Odrv12
    port map (
            O => \N__5306\,
            I => \un1_D_UM_AMIGA_6\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__5303\,
            I => \N__5300\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5297\,
            I => \N__5294\
        );

    \I__1225\ : Span12Mux_h
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__1224\ : Span12Mux_v
    port map (
            O => \N__5291\,
            I => \N__5288\
        );

    \I__1223\ : Odrv12
    port map (
            O => \N__5288\,
            I => \TS_CPUn_c\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5285\,
            I => \N__5282\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5282\,
            I => \N__5270\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5265\
        );

    \I__1219\ : InMux
    port map (
            O => \N__5280\,
            I => \N__5265\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5254\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5278\,
            I => \N__5254\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5277\,
            I => \N__5254\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5254\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5254\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5274\,
            I => \N__5249\
        );

    \I__1212\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5249\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__5270\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__5265\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__5254\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__5249\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5237\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__5237\,
            I => \U111_CYCLE_SM.TS_EN_4\
        );

    \I__1205\ : CEMux
    port map (
            O => \N__5234\,
            I => \N__5227\
        );

    \I__1204\ : CEMux
    port map (
            O => \N__5233\,
            I => \N__5224\
        );

    \I__1203\ : CEMux
    port map (
            O => \N__5232\,
            I => \N__5221\
        );

    \I__1202\ : CEMux
    port map (
            O => \N__5231\,
            I => \N__5218\
        );

    \I__1201\ : CEMux
    port map (
            O => \N__5230\,
            I => \N__5215\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5227\,
            I => \N__5210\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5224\,
            I => \N__5210\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5221\,
            I => \N__5205\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5218\,
            I => \N__5205\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5215\,
            I => \N__5202\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__5210\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1194\ : Odrv4
    port map (
            O => \N__5205\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1193\ : Odrv4
    port map (
            O => \N__5202\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1192\ : SRMux
    port map (
            O => \N__5195\,
            I => \N__5190\
        );

    \I__1191\ : SRMux
    port map (
            O => \N__5194\,
            I => \N__5185\
        );

    \I__1190\ : SRMux
    port map (
            O => \N__5193\,
            I => \N__5182\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5190\,
            I => \N__5179\
        );

    \I__1188\ : SRMux
    port map (
            O => \N__5189\,
            I => \N__5176\
        );

    \I__1187\ : SRMux
    port map (
            O => \N__5188\,
            I => \N__5173\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5185\,
            I => \N__5170\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__5182\,
            I => \N__5167\
        );

    \I__1184\ : Span4Mux_h
    port map (
            O => \N__5179\,
            I => \N__5162\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5176\,
            I => \N__5162\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__5173\,
            I => \N__5159\
        );

    \I__1181\ : Span4Mux_h
    port map (
            O => \N__5170\,
            I => \N__5154\
        );

    \I__1180\ : Span4Mux_h
    port map (
            O => \N__5167\,
            I => \N__5154\
        );

    \I__1179\ : Span4Mux_h
    port map (
            O => \N__5162\,
            I => \N__5149\
        );

    \I__1178\ : Span4Mux_h
    port map (
            O => \N__5159\,
            I => \N__5149\
        );

    \I__1177\ : Odrv4
    port map (
            O => \N__5154\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__5149\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5141\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__5141\,
            I => \N__5136\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5140\,
            I => \N__5133\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5139\,
            I => \N__5130\
        );

    \I__1171\ : Span4Mux_v
    port map (
            O => \N__5136\,
            I => \N__5127\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5133\,
            I => \N__5124\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__5130\,
            I => \N__5121\
        );

    \I__1168\ : Span4Mux_v
    port map (
            O => \N__5127\,
            I => \N__5118\
        );

    \I__1167\ : Span4Mux_v
    port map (
            O => \N__5124\,
            I => \N__5115\
        );

    \I__1166\ : Span4Mux_h
    port map (
            O => \N__5121\,
            I => \N__5112\
        );

    \I__1165\ : Sp12to4
    port map (
            O => \N__5118\,
            I => \N__5109\
        );

    \I__1164\ : Span4Mux_v
    port map (
            O => \N__5115\,
            I => \N__5106\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__5112\,
            I => \N__5103\
        );

    \I__1162\ : Span12Mux_h
    port map (
            O => \N__5109\,
            I => \N__5100\
        );

    \I__1161\ : Sp12to4
    port map (
            O => \N__5106\,
            I => \N__5095\
        );

    \I__1160\ : Sp12to4
    port map (
            O => \N__5103\,
            I => \N__5095\
        );

    \I__1159\ : Span12Mux_v
    port map (
            O => \N__5100\,
            I => \N__5090\
        );

    \I__1158\ : Span12Mux_h
    port map (
            O => \N__5095\,
            I => \N__5090\
        );

    \I__1157\ : Odrv12
    port map (
            O => \N__5090\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5084\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__5084\,
            I => \N__5081\
        );

    \I__1154\ : Odrv12
    port map (
            O => \N__5081\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__1153\ : IoInMux
    port map (
            O => \N__5078\,
            I => \N__5075\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5075\,
            I => \N__5072\
        );

    \I__1151\ : Span4Mux_s2_h
    port map (
            O => \N__5072\,
            I => \N__5069\
        );

    \I__1150\ : Span4Mux_h
    port map (
            O => \N__5069\,
            I => \N__5066\
        );

    \I__1149\ : Sp12to4
    port map (
            O => \N__5066\,
            I => \N__5063\
        );

    \I__1148\ : Span12Mux_s9_v
    port map (
            O => \N__5063\,
            I => \N__5060\
        );

    \I__1147\ : Odrv12
    port map (
            O => \N__5060\,
            I => \un1_D_UM_AMIGA_3\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5054\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5054\,
            I => \N__5051\
        );

    \I__1144\ : Odrv12
    port map (
            O => \N__5051\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5048\,
            I => \N__5044\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5041\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5044\,
            I => \N__5037\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5041\,
            I => \N__5034\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5031\
        );

    \I__1138\ : Span4Mux_v
    port map (
            O => \N__5037\,
            I => \N__5028\
        );

    \I__1137\ : Span4Mux_h
    port map (
            O => \N__5034\,
            I => \N__5025\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__5031\,
            I => \N__5022\
        );

    \I__1135\ : Sp12to4
    port map (
            O => \N__5028\,
            I => \N__5019\
        );

    \I__1134\ : Span4Mux_v
    port map (
            O => \N__5025\,
            I => \N__5014\
        );

    \I__1133\ : Span4Mux_h
    port map (
            O => \N__5022\,
            I => \N__5014\
        );

    \I__1132\ : Span12Mux_h
    port map (
            O => \N__5019\,
            I => \N__5011\
        );

    \I__1131\ : Span4Mux_v
    port map (
            O => \N__5014\,
            I => \N__5008\
        );

    \I__1130\ : Span12Mux_v
    port map (
            O => \N__5011\,
            I => \N__5005\
        );

    \I__1129\ : Sp12to4
    port map (
            O => \N__5008\,
            I => \N__5002\
        );

    \I__1128\ : Odrv12
    port map (
            O => \N__5005\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1127\ : Odrv12
    port map (
            O => \N__5002\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1126\ : IoInMux
    port map (
            O => \N__4997\,
            I => \N__4994\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__1124\ : Span4Mux_s1_h
    port map (
            O => \N__4991\,
            I => \N__4988\
        );

    \I__1123\ : Span4Mux_h
    port map (
            O => \N__4988\,
            I => \N__4985\
        );

    \I__1122\ : Sp12to4
    port map (
            O => \N__4985\,
            I => \N__4982\
        );

    \I__1121\ : Span12Mux_s10_v
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__1120\ : Span12Mux_h
    port map (
            O => \N__4979\,
            I => \N__4976\
        );

    \I__1119\ : Odrv12
    port map (
            O => \N__4976\,
            I => \un1_D_UM_AMIGA_7\
        );

    \I__1118\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4970\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__4970\,
            I => \N__4967\
        );

    \I__1116\ : Span4Mux_v
    port map (
            O => \N__4967\,
            I => \N__4964\
        );

    \I__1115\ : Sp12to4
    port map (
            O => \N__4964\,
            I => \N__4961\
        );

    \I__1114\ : Span12Mux_h
    port map (
            O => \N__4961\,
            I => \N__4958\
        );

    \I__1113\ : Odrv12
    port map (
            O => \N__4958\,
            I => \D_LL_AMIGA_in_5\
        );

    \I__1112\ : IoInMux
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__1110\ : IoSpan4Mux
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__1109\ : Span4Mux_s3_h
    port map (
            O => \N__4946\,
            I => \N__4943\
        );

    \I__1108\ : Sp12to4
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__1107\ : Span12Mux_h
    port map (
            O => \N__4940\,
            I => \N__4937\
        );

    \I__1106\ : Odrv12
    port map (
            O => \N__4937\,
            I => \un1_D_LL_AMIGA_5\
        );

    \I__1105\ : InMux
    port map (
            O => \N__4934\,
            I => \N__4931\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__1103\ : Span4Mux_v
    port map (
            O => \N__4928\,
            I => \N__4925\
        );

    \I__1102\ : Sp12to4
    port map (
            O => \N__4925\,
            I => \N__4922\
        );

    \I__1101\ : Span12Mux_h
    port map (
            O => \N__4922\,
            I => \N__4919\
        );

    \I__1100\ : Odrv12
    port map (
            O => \N__4919\,
            I => \D_LL_AMIGA_in_7\
        );

    \I__1099\ : IoInMux
    port map (
            O => \N__4916\,
            I => \N__4913\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__4913\,
            I => \N__4910\
        );

    \I__1097\ : Span4Mux_s2_h
    port map (
            O => \N__4910\,
            I => \N__4907\
        );

    \I__1096\ : Span4Mux_v
    port map (
            O => \N__4907\,
            I => \N__4904\
        );

    \I__1095\ : Span4Mux_v
    port map (
            O => \N__4904\,
            I => \N__4901\
        );

    \I__1094\ : Sp12to4
    port map (
            O => \N__4901\,
            I => \N__4898\
        );

    \I__1093\ : Span12Mux_s9_h
    port map (
            O => \N__4898\,
            I => \N__4895\
        );

    \I__1092\ : Odrv12
    port map (
            O => \N__4895\,
            I => \un1_D_LL_AMIGA_7\
        );

    \I__1091\ : InMux
    port map (
            O => \N__4892\,
            I => \N__4889\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__4889\,
            I => \N__4886\
        );

    \I__1089\ : Sp12to4
    port map (
            O => \N__4886\,
            I => \N__4883\
        );

    \I__1088\ : Span12Mux_h
    port map (
            O => \N__4883\,
            I => \N__4880\
        );

    \I__1087\ : Odrv12
    port map (
            O => \N__4880\,
            I => \D_UM_040_in_2\
        );

    \I__1086\ : IoInMux
    port map (
            O => \N__4877\,
            I => \N__4874\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__4874\,
            I => \N__4870\
        );

    \I__1084\ : InMux
    port map (
            O => \N__4873\,
            I => \N__4867\
        );

    \I__1083\ : IoSpan4Mux
    port map (
            O => \N__4870\,
            I => \N__4864\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__4867\,
            I => \N__4861\
        );

    \I__1081\ : Span4Mux_s2_h
    port map (
            O => \N__4864\,
            I => \N__4858\
        );

    \I__1080\ : Span4Mux_v
    port map (
            O => \N__4861\,
            I => \N__4855\
        );

    \I__1079\ : Sp12to4
    port map (
            O => \N__4858\,
            I => \N__4852\
        );

    \I__1078\ : Sp12to4
    port map (
            O => \N__4855\,
            I => \N__4849\
        );

    \I__1077\ : Span12Mux_h
    port map (
            O => \N__4852\,
            I => \N__4846\
        );

    \I__1076\ : Span12Mux_h
    port map (
            O => \N__4849\,
            I => \N__4843\
        );

    \I__1075\ : Span12Mux_h
    port map (
            O => \N__4846\,
            I => \N__4838\
        );

    \I__1074\ : Span12Mux_v
    port map (
            O => \N__4843\,
            I => \N__4838\
        );

    \I__1073\ : Odrv12
    port map (
            O => \N__4838\,
            I => \D_LL_040_in_2\
        );

    \I__1072\ : IoInMux
    port map (
            O => \N__4835\,
            I => \N__4832\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__1070\ : Span4Mux_s3_h
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__1069\ : Span4Mux_v
    port map (
            O => \N__4826\,
            I => \N__4823\
        );

    \I__1068\ : Sp12to4
    port map (
            O => \N__4823\,
            I => \N__4820\
        );

    \I__1067\ : Span12Mux_s10_h
    port map (
            O => \N__4820\,
            I => \N__4817\
        );

    \I__1066\ : Odrv12
    port map (
            O => \N__4817\,
            I => \un1_D_UM_040_2\
        );

    \I__1065\ : IoInMux
    port map (
            O => \N__4814\,
            I => \N__4811\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__4811\,
            I => \N__4808\
        );

    \I__1063\ : Span12Mux_s5_h
    port map (
            O => \N__4808\,
            I => \N__4805\
        );

    \I__1062\ : Span12Mux_h
    port map (
            O => \N__4805\,
            I => \N__4802\
        );

    \I__1061\ : Odrv12
    port map (
            O => \N__4802\,
            I => \un1_D_UM_AMIGA_2\
        );

    \I__1060\ : InMux
    port map (
            O => \N__4799\,
            I => \N__4794\
        );

    \I__1059\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4791\
        );

    \I__1058\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4788\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__4794\,
            I => \N__4783\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__4791\,
            I => \N__4783\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__4788\,
            I => \N__4780\
        );

    \I__1054\ : Span4Mux_v
    port map (
            O => \N__4783\,
            I => \N__4777\
        );

    \I__1053\ : Sp12to4
    port map (
            O => \N__4780\,
            I => \N__4774\
        );

    \I__1052\ : Sp12to4
    port map (
            O => \N__4777\,
            I => \N__4771\
        );

    \I__1051\ : Span12Mux_v
    port map (
            O => \N__4774\,
            I => \N__4768\
        );

    \I__1050\ : Span12Mux_h
    port map (
            O => \N__4771\,
            I => \N__4765\
        );

    \I__1049\ : Odrv12
    port map (
            O => \N__4768\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1048\ : Odrv12
    port map (
            O => \N__4765\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1047\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__4757\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__4754\,
            I => \N__4749\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__4753\,
            I => \N__4743\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__4752\,
            I => \N__4739\
        );

    \I__1042\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4735\
        );

    \I__1041\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4730\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4747\,
            I => \N__4730\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4746\,
            I => \N__4723\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4723\
        );

    \I__1037\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4723\
        );

    \I__1036\ : InMux
    port map (
            O => \N__4739\,
            I => \N__4720\
        );

    \I__1035\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4717\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__4735\,
            I => \N__4706\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__4730\,
            I => \N__4706\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__4723\,
            I => \N__4706\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4720\,
            I => \N__4706\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__4717\,
            I => \N__4706\
        );

    \I__1029\ : Span4Mux_v
    port map (
            O => \N__4706\,
            I => \N__4703\
        );

    \I__1028\ : Span4Mux_h
    port map (
            O => \N__4703\,
            I => \N__4699\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4696\
        );

    \I__1026\ : Sp12to4
    port map (
            O => \N__4699\,
            I => \N__4693\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__4696\,
            I => \N__4690\
        );

    \I__1024\ : Span12Mux_s11_h
    port map (
            O => \N__4693\,
            I => \N__4685\
        );

    \I__1023\ : Span12Mux_v
    port map (
            O => \N__4690\,
            I => \N__4685\
        );

    \I__1022\ : Span12Mux_v
    port map (
            O => \N__4685\,
            I => \N__4682\
        );

    \I__1021\ : Odrv12
    port map (
            O => \N__4682\,
            I => \RESETn_c\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4676\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__4676\,
            I => \N__4673\
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__4673\,
            I => \U111_CYCLE_SM.TA_ENZ0\
        );

    \I__1017\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4661\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4669\,
            I => \N__4661\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4668\,
            I => \N__4658\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4667\,
            I => \N__4653\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4653\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__4661\,
            I => \N__4648\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4658\,
            I => \N__4648\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4653\,
            I => \N__4645\
        );

    \I__1009\ : Sp12to4
    port map (
            O => \N__4648\,
            I => \N__4640\
        );

    \I__1008\ : Sp12to4
    port map (
            O => \N__4645\,
            I => \N__4640\
        );

    \I__1007\ : Span12Mux_v
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__1006\ : Odrv12
    port map (
            O => \N__4637\,
            I => \TACKn_c\
        );

    \I__1005\ : IoInMux
    port map (
            O => \N__4634\,
            I => \N__4631\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__4631\,
            I => \N__4628\
        );

    \I__1003\ : Span4Mux_s3_v
    port map (
            O => \N__4628\,
            I => \N__4625\
        );

    \I__1002\ : Sp12to4
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__1001\ : Span12Mux_h
    port map (
            O => \N__4622\,
            I => \N__4619\
        );

    \I__1000\ : Odrv12
    port map (
            O => \N__4619\,
            I => \TAn_0_i\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__4616\,
            I => \N__4609\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__4615\,
            I => \N__4606\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__4614\,
            I => \N__4602\
        );

    \I__996\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4598\
        );

    \I__995\ : InMux
    port map (
            O => \N__4612\,
            I => \N__4595\
        );

    \I__994\ : InMux
    port map (
            O => \N__4609\,
            I => \N__4588\
        );

    \I__993\ : InMux
    port map (
            O => \N__4606\,
            I => \N__4588\
        );

    \I__992\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4588\
        );

    \I__991\ : InMux
    port map (
            O => \N__4602\,
            I => \N__4583\
        );

    \I__990\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4583\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4598\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4595\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4588\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__4583\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__985\ : InMux
    port map (
            O => \N__4574\,
            I => \N__4571\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4571\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__983\ : InMux
    port map (
            O => \N__4568\,
            I => \N__4565\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4565\,
            I => \N__4561\
        );

    \I__981\ : InMux
    port map (
            O => \N__4564\,
            I => \N__4558\
        );

    \I__980\ : Span4Mux_v
    port map (
            O => \N__4561\,
            I => \N__4554\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4558\,
            I => \N__4551\
        );

    \I__978\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4548\
        );

    \I__977\ : Sp12to4
    port map (
            O => \N__4554\,
            I => \N__4545\
        );

    \I__976\ : Span4Mux_v
    port map (
            O => \N__4551\,
            I => \N__4542\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__4548\,
            I => \N__4539\
        );

    \I__974\ : Span12Mux_h
    port map (
            O => \N__4545\,
            I => \N__4536\
        );

    \I__973\ : Sp12to4
    port map (
            O => \N__4542\,
            I => \N__4531\
        );

    \I__972\ : Span12Mux_v
    port map (
            O => \N__4539\,
            I => \N__4531\
        );

    \I__971\ : Span12Mux_v
    port map (
            O => \N__4536\,
            I => \N__4528\
        );

    \I__970\ : Span12Mux_h
    port map (
            O => \N__4531\,
            I => \N__4525\
        );

    \I__969\ : Odrv12
    port map (
            O => \N__4528\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__968\ : Odrv12
    port map (
            O => \N__4525\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__967\ : IoInMux
    port map (
            O => \N__4520\,
            I => \N__4517\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__965\ : Span4Mux_s2_h
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__964\ : Sp12to4
    port map (
            O => \N__4511\,
            I => \N__4508\
        );

    \I__963\ : Span12Mux_s11_v
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__962\ : Span12Mux_h
    port map (
            O => \N__4505\,
            I => \N__4502\
        );

    \I__961\ : Odrv12
    port map (
            O => \N__4502\,
            I => \un1_D_UM_AMIGA_1\
        );

    \I__960\ : InMux
    port map (
            O => \N__4499\,
            I => \N__4496\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4496\,
            I => \N__4492\
        );

    \I__958\ : InMux
    port map (
            O => \N__4495\,
            I => \N__4489\
        );

    \I__957\ : Span4Mux_v
    port map (
            O => \N__4492\,
            I => \N__4483\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4489\,
            I => \N__4483\
        );

    \I__955\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4480\
        );

    \I__954\ : Span4Mux_v
    port map (
            O => \N__4483\,
            I => \N__4475\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4480\,
            I => \N__4475\
        );

    \I__952\ : Span4Mux_h
    port map (
            O => \N__4475\,
            I => \N__4472\
        );

    \I__951\ : Span4Mux_v
    port map (
            O => \N__4472\,
            I => \N__4469\
        );

    \I__950\ : Sp12to4
    port map (
            O => \N__4469\,
            I => \N__4466\
        );

    \I__949\ : Odrv12
    port map (
            O => \N__4466\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__948\ : InMux
    port map (
            O => \N__4463\,
            I => \N__4460\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4460\,
            I => \N__4457\
        );

    \I__946\ : Odrv4
    port map (
            O => \N__4457\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__945\ : IoInMux
    port map (
            O => \N__4454\,
            I => \N__4451\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4451\,
            I => \N__4448\
        );

    \I__943\ : IoSpan4Mux
    port map (
            O => \N__4448\,
            I => \N__4445\
        );

    \I__942\ : IoSpan4Mux
    port map (
            O => \N__4445\,
            I => \N__4442\
        );

    \I__941\ : Sp12to4
    port map (
            O => \N__4442\,
            I => \N__4439\
        );

    \I__940\ : Span12Mux_s9_h
    port map (
            O => \N__4439\,
            I => \N__4436\
        );

    \I__939\ : Odrv12
    port map (
            O => \N__4436\,
            I => \un1_D_UU_AMIGA_1\
        );

    \I__938\ : InMux
    port map (
            O => \N__4433\,
            I => \N__4430\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__936\ : Odrv12
    port map (
            O => \N__4427\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__935\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4420\
        );

    \I__934\ : InMux
    port map (
            O => \N__4423\,
            I => \N__4416\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4420\,
            I => \N__4413\
        );

    \I__932\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4410\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4416\,
            I => \N__4407\
        );

    \I__930\ : Span4Mux_h
    port map (
            O => \N__4413\,
            I => \N__4404\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4410\,
            I => \N__4401\
        );

    \I__928\ : Span12Mux_v
    port map (
            O => \N__4407\,
            I => \N__4398\
        );

    \I__927\ : Span4Mux_v
    port map (
            O => \N__4404\,
            I => \N__4393\
        );

    \I__926\ : Span4Mux_h
    port map (
            O => \N__4401\,
            I => \N__4393\
        );

    \I__925\ : Span12Mux_h
    port map (
            O => \N__4398\,
            I => \N__4390\
        );

    \I__924\ : Span4Mux_v
    port map (
            O => \N__4393\,
            I => \N__4387\
        );

    \I__923\ : Span12Mux_v
    port map (
            O => \N__4390\,
            I => \N__4384\
        );

    \I__922\ : Sp12to4
    port map (
            O => \N__4387\,
            I => \N__4381\
        );

    \I__921\ : Odrv12
    port map (
            O => \N__4384\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__920\ : Odrv12
    port map (
            O => \N__4381\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__919\ : IoInMux
    port map (
            O => \N__4376\,
            I => \N__4373\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__917\ : Span4Mux_s0_v
    port map (
            O => \N__4370\,
            I => \N__4367\
        );

    \I__916\ : Span4Mux_v
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__915\ : Span4Mux_v
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__914\ : Sp12to4
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__913\ : Span12Mux_s11_h
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__912\ : Odrv12
    port map (
            O => \N__4355\,
            I => \un1_D_UM_AMIGA_4\
        );

    \I__911\ : InMux
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__909\ : Span4Mux_v
    port map (
            O => \N__4346\,
            I => \N__4343\
        );

    \I__908\ : Sp12to4
    port map (
            O => \N__4343\,
            I => \N__4340\
        );

    \I__907\ : Span12Mux_h
    port map (
            O => \N__4340\,
            I => \N__4337\
        );

    \I__906\ : Odrv12
    port map (
            O => \N__4337\,
            I => \D_UU_040_in_0\
        );

    \I__905\ : IoInMux
    port map (
            O => \N__4334\,
            I => \N__4331\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__4331\,
            I => \N__4328\
        );

    \I__903\ : IoSpan4Mux
    port map (
            O => \N__4328\,
            I => \N__4324\
        );

    \I__902\ : InMux
    port map (
            O => \N__4327\,
            I => \N__4321\
        );

    \I__901\ : IoSpan4Mux
    port map (
            O => \N__4324\,
            I => \N__4318\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4321\,
            I => \N__4315\
        );

    \I__899\ : Span4Mux_s2_h
    port map (
            O => \N__4318\,
            I => \N__4312\
        );

    \I__898\ : Span12Mux_v
    port map (
            O => \N__4315\,
            I => \N__4309\
        );

    \I__897\ : Sp12to4
    port map (
            O => \N__4312\,
            I => \N__4306\
        );

    \I__896\ : Span12Mux_h
    port map (
            O => \N__4309\,
            I => \N__4303\
        );

    \I__895\ : Span12Mux_h
    port map (
            O => \N__4306\,
            I => \N__4300\
        );

    \I__894\ : Span12Mux_v
    port map (
            O => \N__4303\,
            I => \N__4295\
        );

    \I__893\ : Span12Mux_h
    port map (
            O => \N__4300\,
            I => \N__4295\
        );

    \I__892\ : Odrv12
    port map (
            O => \N__4295\,
            I => \D_LM_040_in_0\
        );

    \I__891\ : IoInMux
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4289\,
            I => \N__4286\
        );

    \I__889\ : IoSpan4Mux
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__888\ : Sp12to4
    port map (
            O => \N__4283\,
            I => \N__4280\
        );

    \I__887\ : Span12Mux_s6_v
    port map (
            O => \N__4280\,
            I => \N__4277\
        );

    \I__886\ : Odrv12
    port map (
            O => \N__4277\,
            I => \un1_D_UU_040_0\
        );

    \I__885\ : InMux
    port map (
            O => \N__4274\,
            I => \N__4271\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4271\,
            I => \N__4268\
        );

    \I__883\ : Sp12to4
    port map (
            O => \N__4268\,
            I => \N__4265\
        );

    \I__882\ : Span12Mux_s7_v
    port map (
            O => \N__4265\,
            I => \N__4262\
        );

    \I__881\ : Span12Mux_h
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__880\ : Odrv12
    port map (
            O => \N__4259\,
            I => \D_UU_040_in_2\
        );

    \I__879\ : IoInMux
    port map (
            O => \N__4256\,
            I => \N__4252\
        );

    \I__878\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4249\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__4252\,
            I => \N__4246\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4249\,
            I => \N__4243\
        );

    \I__875\ : Span12Mux_s9_h
    port map (
            O => \N__4246\,
            I => \N__4240\
        );

    \I__874\ : Span12Mux_v
    port map (
            O => \N__4243\,
            I => \N__4237\
        );

    \I__873\ : Span12Mux_v
    port map (
            O => \N__4240\,
            I => \N__4234\
        );

    \I__872\ : Span12Mux_h
    port map (
            O => \N__4237\,
            I => \N__4231\
        );

    \I__871\ : Span12Mux_h
    port map (
            O => \N__4234\,
            I => \N__4228\
        );

    \I__870\ : Span12Mux_v
    port map (
            O => \N__4231\,
            I => \N__4225\
        );

    \I__869\ : Odrv12
    port map (
            O => \N__4228\,
            I => \D_LM_040_in_2\
        );

    \I__868\ : Odrv12
    port map (
            O => \N__4225\,
            I => \D_LM_040_in_2\
        );

    \I__867\ : IoInMux
    port map (
            O => \N__4220\,
            I => \N__4217\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__865\ : IoSpan4Mux
    port map (
            O => \N__4214\,
            I => \N__4211\
        );

    \I__864\ : IoSpan4Mux
    port map (
            O => \N__4211\,
            I => \N__4208\
        );

    \I__863\ : Span4Mux_s3_v
    port map (
            O => \N__4208\,
            I => \N__4205\
        );

    \I__862\ : Odrv4
    port map (
            O => \N__4205\,
            I => \un1_D_UU_040_2\
        );

    \I__861\ : InMux
    port map (
            O => \N__4202\,
            I => \N__4199\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__859\ : Span4Mux_v
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__858\ : Odrv4
    port map (
            O => \N__4193\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__857\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4187\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4187\,
            I => \N__4184\
        );

    \I__855\ : Span4Mux_h
    port map (
            O => \N__4184\,
            I => \N__4180\
        );

    \I__854\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4177\
        );

    \I__853\ : Span4Mux_v
    port map (
            O => \N__4180\,
            I => \N__4172\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4177\,
            I => \N__4172\
        );

    \I__851\ : Span4Mux_v
    port map (
            O => \N__4172\,
            I => \N__4168\
        );

    \I__850\ : InMux
    port map (
            O => \N__4171\,
            I => \N__4165\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__4168\,
            I => \N__4160\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4165\,
            I => \N__4160\
        );

    \I__847\ : Span4Mux_v
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__846\ : Span4Mux_h
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__845\ : Span4Mux_h
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__4151\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__843\ : IoInMux
    port map (
            O => \N__4148\,
            I => \N__4145\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4145\,
            I => \N__4142\
        );

    \I__841\ : IoSpan4Mux
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__840\ : Span4Mux_s2_v
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__839\ : Span4Mux_v
    port map (
            O => \N__4136\,
            I => \N__4133\
        );

    \I__838\ : Sp12to4
    port map (
            O => \N__4133\,
            I => \N__4130\
        );

    \I__837\ : Odrv12
    port map (
            O => \N__4130\,
            I => \un1_D_UU_AMIGA_0\
        );

    \I__836\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4124\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4124\,
            I => \N__4121\
        );

    \I__834\ : Span4Mux_v
    port map (
            O => \N__4121\,
            I => \N__4118\
        );

    \I__833\ : Sp12to4
    port map (
            O => \N__4118\,
            I => \N__4115\
        );

    \I__832\ : Span12Mux_h
    port map (
            O => \N__4115\,
            I => \N__4112\
        );

    \I__831\ : Odrv12
    port map (
            O => \N__4112\,
            I => \D_LL_AMIGA_in_6\
        );

    \I__830\ : IoInMux
    port map (
            O => \N__4109\,
            I => \N__4106\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__828\ : Span4Mux_s2_h
    port map (
            O => \N__4103\,
            I => \N__4100\
        );

    \I__827\ : Span4Mux_v
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__826\ : Span4Mux_v
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__825\ : Sp12to4
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__824\ : Span12Mux_s9_h
    port map (
            O => \N__4091\,
            I => \N__4088\
        );

    \I__823\ : Odrv12
    port map (
            O => \N__4088\,
            I => \un1_D_LL_AMIGA_6\
        );

    \I__822\ : InMux
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4082\,
            I => \U111_CYCLE_SM.TS_EN10\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__819\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4072\
        );

    \I__818\ : InMux
    port map (
            O => \N__4075\,
            I => \N__4069\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4072\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4069\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__815\ : IoInMux
    port map (
            O => \N__4064\,
            I => \N__4061\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__813\ : IoSpan4Mux
    port map (
            O => \N__4058\,
            I => \N__4055\
        );

    \I__812\ : Span4Mux_s2_v
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__811\ : Sp12to4
    port map (
            O => \N__4052\,
            I => \N__4048\
        );

    \I__810\ : InMux
    port map (
            O => \N__4051\,
            I => \N__4045\
        );

    \I__809\ : Odrv12
    port map (
            O => \N__4048\,
            I => \TSn_c\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4045\,
            I => \TSn_c\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__4040\,
            I => \N__4036\
        );

    \I__806\ : InMux
    port map (
            O => \N__4039\,
            I => \N__4031\
        );

    \I__805\ : InMux
    port map (
            O => \N__4036\,
            I => \N__4031\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__4031\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__803\ : IoInMux
    port map (
            O => \N__4028\,
            I => \N__4024\
        );

    \I__802\ : IoInMux
    port map (
            O => \N__4027\,
            I => \N__4021\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4024\,
            I => \N__4014\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4021\,
            I => \N__4014\
        );

    \I__799\ : IoInMux
    port map (
            O => \N__4020\,
            I => \N__4011\
        );

    \I__798\ : IoInMux
    port map (
            O => \N__4019\,
            I => \N__4008\
        );

    \I__797\ : IoSpan4Mux
    port map (
            O => \N__4014\,
            I => \N__3994\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4011\,
            I => \N__3994\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__4008\,
            I => \N__3994\
        );

    \I__794\ : IoInMux
    port map (
            O => \N__4007\,
            I => \N__3991\
        );

    \I__793\ : IoInMux
    port map (
            O => \N__4006\,
            I => \N__3988\
        );

    \I__792\ : IoInMux
    port map (
            O => \N__4005\,
            I => \N__3985\
        );

    \I__791\ : IoInMux
    port map (
            O => \N__4004\,
            I => \N__3982\
        );

    \I__790\ : IoInMux
    port map (
            O => \N__4003\,
            I => \N__3979\
        );

    \I__789\ : IoInMux
    port map (
            O => \N__4002\,
            I => \N__3974\
        );

    \I__788\ : InMux
    port map (
            O => \N__4001\,
            I => \N__3971\
        );

    \I__787\ : IoSpan4Mux
    port map (
            O => \N__3994\,
            I => \N__3956\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__3991\,
            I => \N__3956\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__3988\,
            I => \N__3956\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__3985\,
            I => \N__3956\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__3982\,
            I => \N__3956\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__3979\,
            I => \N__3956\
        );

    \I__781\ : IoInMux
    port map (
            O => \N__3978\,
            I => \N__3953\
        );

    \I__780\ : IoInMux
    port map (
            O => \N__3977\,
            I => \N__3950\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__3974\,
            I => \N__3947\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__3971\,
            I => \N__3944\
        );

    \I__777\ : IoInMux
    port map (
            O => \N__3970\,
            I => \N__3940\
        );

    \I__776\ : IoInMux
    port map (
            O => \N__3969\,
            I => \N__3937\
        );

    \I__775\ : IoSpan4Mux
    port map (
            O => \N__3956\,
            I => \N__3924\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__3953\,
            I => \N__3924\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__3950\,
            I => \N__3924\
        );

    \I__772\ : Span4Mux_s3_v
    port map (
            O => \N__3947\,
            I => \N__3920\
        );

    \I__771\ : Span4Mux_h
    port map (
            O => \N__3944\,
            I => \N__3917\
        );

    \I__770\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3914\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__3940\,
            I => \N__3909\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__3937\,
            I => \N__3909\
        );

    \I__767\ : IoInMux
    port map (
            O => \N__3936\,
            I => \N__3906\
        );

    \I__766\ : IoInMux
    port map (
            O => \N__3935\,
            I => \N__3903\
        );

    \I__765\ : IoInMux
    port map (
            O => \N__3934\,
            I => \N__3900\
        );

    \I__764\ : IoInMux
    port map (
            O => \N__3933\,
            I => \N__3897\
        );

    \I__763\ : IoInMux
    port map (
            O => \N__3932\,
            I => \N__3894\
        );

    \I__762\ : IoInMux
    port map (
            O => \N__3931\,
            I => \N__3891\
        );

    \I__761\ : IoSpan4Mux
    port map (
            O => \N__3924\,
            I => \N__3884\
        );

    \I__760\ : IoInMux
    port map (
            O => \N__3923\,
            I => \N__3881\
        );

    \I__759\ : Span4Mux_v
    port map (
            O => \N__3920\,
            I => \N__3877\
        );

    \I__758\ : Span4Mux_h
    port map (
            O => \N__3917\,
            I => \N__3872\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3914\,
            I => \N__3872\
        );

    \I__756\ : IoSpan4Mux
    port map (
            O => \N__3909\,
            I => \N__3856\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__3906\,
            I => \N__3856\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__3903\,
            I => \N__3856\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__3900\,
            I => \N__3856\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__3897\,
            I => \N__3856\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3894\,
            I => \N__3856\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__3891\,
            I => \N__3856\
        );

    \I__749\ : IoInMux
    port map (
            O => \N__3890\,
            I => \N__3853\
        );

    \I__748\ : IoInMux
    port map (
            O => \N__3889\,
            I => \N__3850\
        );

    \I__747\ : IoInMux
    port map (
            O => \N__3888\,
            I => \N__3847\
        );

    \I__746\ : IoInMux
    port map (
            O => \N__3887\,
            I => \N__3844\
        );

    \I__745\ : IoSpan4Mux
    port map (
            O => \N__3884\,
            I => \N__3839\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__3881\,
            I => \N__3839\
        );

    \I__743\ : IoInMux
    port map (
            O => \N__3880\,
            I => \N__3836\
        );

    \I__742\ : Span4Mux_v
    port map (
            O => \N__3877\,
            I => \N__3830\
        );

    \I__741\ : Span4Mux_v
    port map (
            O => \N__3872\,
            I => \N__3827\
        );

    \I__740\ : IoInMux
    port map (
            O => \N__3871\,
            I => \N__3824\
        );

    \I__739\ : IoSpan4Mux
    port map (
            O => \N__3856\,
            I => \N__3813\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__3853\,
            I => \N__3813\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3850\,
            I => \N__3813\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3847\,
            I => \N__3813\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__3844\,
            I => \N__3813\
        );

    \I__734\ : IoSpan4Mux
    port map (
            O => \N__3839\,
            I => \N__3809\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__3836\,
            I => \N__3806\
        );

    \I__732\ : IoInMux
    port map (
            O => \N__3835\,
            I => \N__3803\
        );

    \I__731\ : IoInMux
    port map (
            O => \N__3834\,
            I => \N__3800\
        );

    \I__730\ : IoInMux
    port map (
            O => \N__3833\,
            I => \N__3797\
        );

    \I__729\ : Sp12to4
    port map (
            O => \N__3830\,
            I => \N__3793\
        );

    \I__728\ : Sp12to4
    port map (
            O => \N__3827\,
            I => \N__3789\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__3824\,
            I => \N__3786\
        );

    \I__726\ : IoSpan4Mux
    port map (
            O => \N__3813\,
            I => \N__3783\
        );

    \I__725\ : IoInMux
    port map (
            O => \N__3812\,
            I => \N__3780\
        );

    \I__724\ : IoSpan4Mux
    port map (
            O => \N__3809\,
            I => \N__3769\
        );

    \I__723\ : IoSpan4Mux
    port map (
            O => \N__3806\,
            I => \N__3769\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__3803\,
            I => \N__3769\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__3800\,
            I => \N__3769\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__3797\,
            I => \N__3769\
        );

    \I__719\ : IoInMux
    port map (
            O => \N__3796\,
            I => \N__3766\
        );

    \I__718\ : Span12Mux_h
    port map (
            O => \N__3793\,
            I => \N__3763\
        );

    \I__717\ : IoInMux
    port map (
            O => \N__3792\,
            I => \N__3760\
        );

    \I__716\ : Span12Mux_h
    port map (
            O => \N__3789\,
            I => \N__3755\
        );

    \I__715\ : Span12Mux_s11_v
    port map (
            O => \N__3786\,
            I => \N__3755\
        );

    \I__714\ : IoSpan4Mux
    port map (
            O => \N__3783\,
            I => \N__3750\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__3780\,
            I => \N__3750\
        );

    \I__712\ : IoSpan4Mux
    port map (
            O => \N__3769\,
            I => \N__3745\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3766\,
            I => \N__3745\
        );

    \I__710\ : Span12Mux_h
    port map (
            O => \N__3763\,
            I => \N__3740\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3760\,
            I => \N__3740\
        );

    \I__708\ : Odrv12
    port map (
            O => \N__3755\,
            I => \RnW_c\
        );

    \I__707\ : Odrv4
    port map (
            O => \N__3750\,
            I => \RnW_c\
        );

    \I__706\ : Odrv4
    port map (
            O => \N__3745\,
            I => \RnW_c\
        );

    \I__705\ : Odrv12
    port map (
            O => \N__3740\,
            I => \RnW_c\
        );

    \I__704\ : CascadeMux
    port map (
            O => \N__3731\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__3728\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_\
        );

    \I__702\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3722\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3722\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\
        );

    \I__700\ : InMux
    port map (
            O => \N__3719\,
            I => \N__3716\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3716\,
            I => \N__3713\
        );

    \I__698\ : Span12Mux_v
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__697\ : Span12Mux_h
    port map (
            O => \N__3710\,
            I => \N__3707\
        );

    \I__696\ : Odrv12
    port map (
            O => \N__3707\,
            I => \D_LM_AMIGA_in_0\
        );

    \I__695\ : IoInMux
    port map (
            O => \N__3704\,
            I => \N__3701\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__3701\,
            I => \N__3698\
        );

    \I__693\ : Span4Mux_s3_h
    port map (
            O => \N__3698\,
            I => \N__3695\
        );

    \I__692\ : Span4Mux_v
    port map (
            O => \N__3695\,
            I => \N__3692\
        );

    \I__691\ : Span4Mux_v
    port map (
            O => \N__3692\,
            I => \N__3689\
        );

    \I__690\ : Span4Mux_h
    port map (
            O => \N__3689\,
            I => \N__3686\
        );

    \I__689\ : Sp12to4
    port map (
            O => \N__3686\,
            I => \N__3683\
        );

    \I__688\ : Odrv12
    port map (
            O => \N__3683\,
            I => \un1_D_LM_AMIGA_0\
        );

    \I__687\ : InMux
    port map (
            O => \N__3680\,
            I => \N__3677\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__3677\,
            I => \N__3674\
        );

    \I__685\ : Span12Mux_h
    port map (
            O => \N__3674\,
            I => \N__3671\
        );

    \I__684\ : Odrv12
    port map (
            O => \N__3671\,
            I => \D_LM_AMIGA_in_1\
        );

    \I__683\ : IoInMux
    port map (
            O => \N__3668\,
            I => \N__3665\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__3665\,
            I => \N__3662\
        );

    \I__681\ : Span4Mux_s0_h
    port map (
            O => \N__3662\,
            I => \N__3659\
        );

    \I__680\ : Span4Mux_h
    port map (
            O => \N__3659\,
            I => \N__3656\
        );

    \I__679\ : Span4Mux_h
    port map (
            O => \N__3656\,
            I => \N__3653\
        );

    \I__678\ : Sp12to4
    port map (
            O => \N__3653\,
            I => \N__3650\
        );

    \I__677\ : Span12Mux_v
    port map (
            O => \N__3650\,
            I => \N__3647\
        );

    \I__676\ : Odrv12
    port map (
            O => \N__3647\,
            I => \un1_D_LM_AMIGA_1\
        );

    \I__675\ : InMux
    port map (
            O => \N__3644\,
            I => \N__3641\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3641\,
            I => \N__3638\
        );

    \I__673\ : Span4Mux_v
    port map (
            O => \N__3638\,
            I => \N__3635\
        );

    \I__672\ : Sp12to4
    port map (
            O => \N__3635\,
            I => \N__3632\
        );

    \I__671\ : Span12Mux_h
    port map (
            O => \N__3632\,
            I => \N__3628\
        );

    \I__670\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3625\
        );

    \I__669\ : Odrv12
    port map (
            O => \N__3628\,
            I => \U111_CYCLE_SM.A_OUTZ0\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3625\,
            I => \U111_CYCLE_SM.A_OUTZ0\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__3620\,
            I => \U111_CYCLE_SM.LW_CYCLE_r_1_cascade_\
        );

    \I__666\ : InMux
    port map (
            O => \N__3617\,
            I => \N__3614\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3614\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__3611\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_cascade_\
        );

    \I__663\ : InMux
    port map (
            O => \N__3608\,
            I => \N__3604\
        );

    \I__662\ : SRMux
    port map (
            O => \N__3607\,
            I => \N__3601\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3604\,
            I => \N__3598\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3601\,
            I => \RESETn_c_i\
        );

    \I__659\ : Odrv12
    port map (
            O => \N__3598\,
            I => \RESETn_c_i\
        );

    \I__658\ : CEMux
    port map (
            O => \N__3593\,
            I => \N__3590\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3590\,
            I => \N__3587\
        );

    \I__656\ : Span4Mux_v
    port map (
            O => \N__3587\,
            I => \N__3584\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__3584\,
            I => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_0\
        );

    \I__654\ : InMux
    port map (
            O => \N__3581\,
            I => \N__3577\
        );

    \I__653\ : IoInMux
    port map (
            O => \N__3580\,
            I => \N__3574\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3577\,
            I => \N__3571\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3574\,
            I => \N__3568\
        );

    \I__650\ : Span4Mux_h
    port map (
            O => \N__3571\,
            I => \N__3565\
        );

    \I__649\ : Span4Mux_s3_h
    port map (
            O => \N__3568\,
            I => \N__3562\
        );

    \I__648\ : Span4Mux_h
    port map (
            O => \N__3565\,
            I => \N__3559\
        );

    \I__647\ : Sp12to4
    port map (
            O => \N__3562\,
            I => \N__3556\
        );

    \I__646\ : Sp12to4
    port map (
            O => \N__3559\,
            I => \N__3553\
        );

    \I__645\ : Span12Mux_v
    port map (
            O => \N__3556\,
            I => \N__3550\
        );

    \I__644\ : Span12Mux_v
    port map (
            O => \N__3553\,
            I => \N__3547\
        );

    \I__643\ : Span12Mux_h
    port map (
            O => \N__3550\,
            I => \N__3544\
        );

    \I__642\ : Span12Mux_v
    port map (
            O => \N__3547\,
            I => \N__3541\
        );

    \I__641\ : Span12Mux_h
    port map (
            O => \N__3544\,
            I => \N__3538\
        );

    \I__640\ : Span12Mux_h
    port map (
            O => \N__3541\,
            I => \N__3535\
        );

    \I__639\ : Odrv12
    port map (
            O => \N__3538\,
            I => \D_LM_040_in_1\
        );

    \I__638\ : Odrv12
    port map (
            O => \N__3535\,
            I => \D_LM_040_in_1\
        );

    \I__637\ : InMux
    port map (
            O => \N__3530\,
            I => \N__3527\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3527\,
            I => \N__3524\
        );

    \I__635\ : Span4Mux_v
    port map (
            O => \N__3524\,
            I => \N__3521\
        );

    \I__634\ : Span4Mux_v
    port map (
            O => \N__3521\,
            I => \N__3518\
        );

    \I__633\ : Sp12to4
    port map (
            O => \N__3518\,
            I => \N__3515\
        );

    \I__632\ : Span12Mux_h
    port map (
            O => \N__3515\,
            I => \N__3512\
        );

    \I__631\ : Odrv12
    port map (
            O => \N__3512\,
            I => \D_UU_040_in_1\
        );

    \I__630\ : IoInMux
    port map (
            O => \N__3509\,
            I => \N__3506\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3506\,
            I => \N__3503\
        );

    \I__628\ : Span4Mux_s3_h
    port map (
            O => \N__3503\,
            I => \N__3500\
        );

    \I__627\ : Sp12to4
    port map (
            O => \N__3500\,
            I => \N__3497\
        );

    \I__626\ : Span12Mux_s8_v
    port map (
            O => \N__3497\,
            I => \N__3494\
        );

    \I__625\ : Odrv12
    port map (
            O => \N__3494\,
            I => \un1_D_UU_040_1\
        );

    \I__624\ : InMux
    port map (
            O => \N__3491\,
            I => \N__3487\
        );

    \I__623\ : InMux
    port map (
            O => \N__3490\,
            I => \N__3484\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3487\,
            I => \N__3481\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3484\,
            I => \N__3478\
        );

    \I__620\ : Span4Mux_v
    port map (
            O => \N__3481\,
            I => \N__3472\
        );

    \I__619\ : Span4Mux_v
    port map (
            O => \N__3478\,
            I => \N__3472\
        );

    \I__618\ : InMux
    port map (
            O => \N__3477\,
            I => \N__3469\
        );

    \I__617\ : Sp12to4
    port map (
            O => \N__3472\,
            I => \N__3464\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__3469\,
            I => \N__3464\
        );

    \I__615\ : Span12Mux_h
    port map (
            O => \N__3464\,
            I => \N__3461\
        );

    \I__614\ : Odrv12
    port map (
            O => \N__3461\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__613\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3455\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3455\,
            I => \N__3452\
        );

    \I__611\ : Odrv12
    port map (
            O => \N__3452\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__610\ : IoInMux
    port map (
            O => \N__3449\,
            I => \N__3446\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3446\,
            I => \N__3443\
        );

    \I__608\ : Span4Mux_s3_v
    port map (
            O => \N__3443\,
            I => \N__3440\
        );

    \I__607\ : Span4Mux_h
    port map (
            O => \N__3440\,
            I => \N__3437\
        );

    \I__606\ : Span4Mux_h
    port map (
            O => \N__3437\,
            I => \N__3434\
        );

    \I__605\ : Span4Mux_h
    port map (
            O => \N__3434\,
            I => \N__3431\
        );

    \I__604\ : Span4Mux_v
    port map (
            O => \N__3431\,
            I => \N__3428\
        );

    \I__603\ : Odrv4
    port map (
            O => \N__3428\,
            I => \un1_D_UU_AMIGA_6\
        );

    \I__602\ : InMux
    port map (
            O => \N__3425\,
            I => \N__3422\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3422\,
            I => \N__3419\
        );

    \I__600\ : Odrv12
    port map (
            O => \N__3419\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__599\ : InMux
    port map (
            O => \N__3416\,
            I => \N__3413\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3413\,
            I => \N__3409\
        );

    \I__597\ : InMux
    port map (
            O => \N__3412\,
            I => \N__3406\
        );

    \I__596\ : Span4Mux_v
    port map (
            O => \N__3409\,
            I => \N__3403\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3406\,
            I => \N__3399\
        );

    \I__594\ : Span4Mux_v
    port map (
            O => \N__3403\,
            I => \N__3396\
        );

    \I__593\ : InMux
    port map (
            O => \N__3402\,
            I => \N__3393\
        );

    \I__592\ : Span4Mux_h
    port map (
            O => \N__3399\,
            I => \N__3390\
        );

    \I__591\ : Sp12to4
    port map (
            O => \N__3396\,
            I => \N__3385\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3393\,
            I => \N__3385\
        );

    \I__589\ : Sp12to4
    port map (
            O => \N__3390\,
            I => \N__3382\
        );

    \I__588\ : Span12Mux_h
    port map (
            O => \N__3385\,
            I => \N__3379\
        );

    \I__587\ : Odrv12
    port map (
            O => \N__3382\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__586\ : Odrv12
    port map (
            O => \N__3379\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__585\ : IoInMux
    port map (
            O => \N__3374\,
            I => \N__3371\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3371\,
            I => \N__3368\
        );

    \I__583\ : Span4Mux_s3_v
    port map (
            O => \N__3368\,
            I => \N__3365\
        );

    \I__582\ : Span4Mux_v
    port map (
            O => \N__3365\,
            I => \N__3362\
        );

    \I__581\ : Sp12to4
    port map (
            O => \N__3362\,
            I => \N__3359\
        );

    \I__580\ : Odrv12
    port map (
            O => \N__3359\,
            I => \un1_D_UU_AMIGA_4\
        );

    \I__579\ : InMux
    port map (
            O => \N__3356\,
            I => \N__3353\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3353\,
            I => \N__3350\
        );

    \I__577\ : Odrv12
    port map (
            O => \N__3350\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__576\ : InMux
    port map (
            O => \N__3347\,
            I => \N__3343\
        );

    \I__575\ : InMux
    port map (
            O => \N__3346\,
            I => \N__3340\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__3343\,
            I => \N__3337\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3340\,
            I => \N__3333\
        );

    \I__572\ : Span4Mux_v
    port map (
            O => \N__3337\,
            I => \N__3330\
        );

    \I__571\ : InMux
    port map (
            O => \N__3336\,
            I => \N__3327\
        );

    \I__570\ : Span4Mux_v
    port map (
            O => \N__3333\,
            I => \N__3324\
        );

    \I__569\ : Sp12to4
    port map (
            O => \N__3330\,
            I => \N__3319\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3327\,
            I => \N__3319\
        );

    \I__567\ : Sp12to4
    port map (
            O => \N__3324\,
            I => \N__3316\
        );

    \I__566\ : Span12Mux_h
    port map (
            O => \N__3319\,
            I => \N__3313\
        );

    \I__565\ : Span12Mux_h
    port map (
            O => \N__3316\,
            I => \N__3310\
        );

    \I__564\ : Odrv12
    port map (
            O => \N__3313\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__563\ : Odrv12
    port map (
            O => \N__3310\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__562\ : IoInMux
    port map (
            O => \N__3305\,
            I => \N__3302\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3302\,
            I => \N__3299\
        );

    \I__560\ : IoSpan4Mux
    port map (
            O => \N__3299\,
            I => \N__3296\
        );

    \I__559\ : Sp12to4
    port map (
            O => \N__3296\,
            I => \N__3293\
        );

    \I__558\ : Span12Mux_s6_v
    port map (
            O => \N__3293\,
            I => \N__3290\
        );

    \I__557\ : Span12Mux_h
    port map (
            O => \N__3290\,
            I => \N__3287\
        );

    \I__556\ : Odrv12
    port map (
            O => \N__3287\,
            I => \un1_D_UU_AMIGA_7\
        );

    \I__555\ : InMux
    port map (
            O => \N__3284\,
            I => \N__3281\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3281\,
            I => \N__3278\
        );

    \I__553\ : Span4Mux_v
    port map (
            O => \N__3278\,
            I => \N__3275\
        );

    \I__552\ : Sp12to4
    port map (
            O => \N__3275\,
            I => \N__3272\
        );

    \I__551\ : Span12Mux_h
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__550\ : Odrv12
    port map (
            O => \N__3269\,
            I => \D_LL_AMIGA_in_4\
        );

    \I__549\ : IoInMux
    port map (
            O => \N__3266\,
            I => \N__3263\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3263\,
            I => \N__3260\
        );

    \I__547\ : IoSpan4Mux
    port map (
            O => \N__3260\,
            I => \N__3257\
        );

    \I__546\ : IoSpan4Mux
    port map (
            O => \N__3257\,
            I => \N__3254\
        );

    \I__545\ : Sp12to4
    port map (
            O => \N__3254\,
            I => \N__3251\
        );

    \I__544\ : Span12Mux_s9_h
    port map (
            O => \N__3251\,
            I => \N__3248\
        );

    \I__543\ : Odrv12
    port map (
            O => \N__3248\,
            I => \un1_D_LL_AMIGA_4\
        );

    \I__542\ : InMux
    port map (
            O => \N__3245\,
            I => \N__3242\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3242\,
            I => \N__3239\
        );

    \I__540\ : Sp12to4
    port map (
            O => \N__3239\,
            I => \N__3236\
        );

    \I__539\ : Span12Mux_v
    port map (
            O => \N__3236\,
            I => \N__3233\
        );

    \I__538\ : Odrv12
    port map (
            O => \N__3233\,
            I => \D_LM_AMIGA_in_7\
        );

    \I__537\ : IoInMux
    port map (
            O => \N__3230\,
            I => \N__3227\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3227\,
            I => \N__3224\
        );

    \I__535\ : IoSpan4Mux
    port map (
            O => \N__3224\,
            I => \N__3221\
        );

    \I__534\ : Span4Mux_s0_h
    port map (
            O => \N__3221\,
            I => \N__3218\
        );

    \I__533\ : Sp12to4
    port map (
            O => \N__3218\,
            I => \N__3215\
        );

    \I__532\ : Span12Mux_h
    port map (
            O => \N__3215\,
            I => \N__3212\
        );

    \I__531\ : Odrv12
    port map (
            O => \N__3212\,
            I => \un1_D_LM_AMIGA_7\
        );

    \I__530\ : InMux
    port map (
            O => \N__3209\,
            I => \N__3206\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3206\,
            I => \N__3202\
        );

    \I__528\ : IoInMux
    port map (
            O => \N__3205\,
            I => \N__3199\
        );

    \I__527\ : Span12Mux_v
    port map (
            O => \N__3202\,
            I => \N__3196\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3199\,
            I => \N__3193\
        );

    \I__525\ : Odrv12
    port map (
            O => \N__3196\,
            I => \A_AMIGA_c_1\
        );

    \I__524\ : Odrv12
    port map (
            O => \N__3193\,
            I => \A_AMIGA_c_1\
        );

    \I__523\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3185\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3185\,
            I => \N__3182\
        );

    \I__521\ : Span12Mux_v
    port map (
            O => \N__3182\,
            I => \N__3179\
        );

    \I__520\ : Span12Mux_h
    port map (
            O => \N__3179\,
            I => \N__3176\
        );

    \I__519\ : Odrv12
    port map (
            O => \N__3176\,
            I => \D_UM_040_in_7\
        );

    \I__518\ : IoInMux
    port map (
            O => \N__3173\,
            I => \N__3170\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3170\,
            I => \N__3167\
        );

    \I__516\ : IoSpan4Mux
    port map (
            O => \N__3167\,
            I => \N__3163\
        );

    \I__515\ : InMux
    port map (
            O => \N__3166\,
            I => \N__3160\
        );

    \I__514\ : Span4Mux_s3_h
    port map (
            O => \N__3163\,
            I => \N__3157\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3160\,
            I => \N__3154\
        );

    \I__512\ : Sp12to4
    port map (
            O => \N__3157\,
            I => \N__3151\
        );

    \I__511\ : Span12Mux_v
    port map (
            O => \N__3154\,
            I => \N__3148\
        );

    \I__510\ : Span12Mux_v
    port map (
            O => \N__3151\,
            I => \N__3145\
        );

    \I__509\ : Span12Mux_v
    port map (
            O => \N__3148\,
            I => \N__3142\
        );

    \I__508\ : Span12Mux_h
    port map (
            O => \N__3145\,
            I => \N__3139\
        );

    \I__507\ : Span12Mux_h
    port map (
            O => \N__3142\,
            I => \N__3136\
        );

    \I__506\ : Span12Mux_h
    port map (
            O => \N__3139\,
            I => \N__3133\
        );

    \I__505\ : Odrv12
    port map (
            O => \N__3136\,
            I => \D_LL_040_in_7\
        );

    \I__504\ : Odrv12
    port map (
            O => \N__3133\,
            I => \D_LL_040_in_7\
        );

    \I__503\ : IoInMux
    port map (
            O => \N__3128\,
            I => \N__3125\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3125\,
            I => \N__3122\
        );

    \I__501\ : Span4Mux_s3_h
    port map (
            O => \N__3122\,
            I => \N__3119\
        );

    \I__500\ : Span4Mux_h
    port map (
            O => \N__3119\,
            I => \N__3116\
        );

    \I__499\ : Span4Mux_h
    port map (
            O => \N__3116\,
            I => \N__3113\
        );

    \I__498\ : Odrv4
    port map (
            O => \N__3113\,
            I => \un1_D_UM_040_7\
        );

    \I__497\ : IoInMux
    port map (
            O => \N__3110\,
            I => \N__3107\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3107\,
            I => \N__3103\
        );

    \I__495\ : InMux
    port map (
            O => \N__3106\,
            I => \N__3100\
        );

    \I__494\ : Span4Mux_s2_h
    port map (
            O => \N__3103\,
            I => \N__3097\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3100\,
            I => \N__3094\
        );

    \I__492\ : Span4Mux_v
    port map (
            O => \N__3097\,
            I => \N__3091\
        );

    \I__491\ : Span4Mux_v
    port map (
            O => \N__3094\,
            I => \N__3088\
        );

    \I__490\ : Sp12to4
    port map (
            O => \N__3091\,
            I => \N__3085\
        );

    \I__489\ : Span4Mux_v
    port map (
            O => \N__3088\,
            I => \N__3082\
        );

    \I__488\ : Span12Mux_h
    port map (
            O => \N__3085\,
            I => \N__3077\
        );

    \I__487\ : Sp12to4
    port map (
            O => \N__3082\,
            I => \N__3077\
        );

    \I__486\ : Span12Mux_h
    port map (
            O => \N__3077\,
            I => \N__3074\
        );

    \I__485\ : Odrv12
    port map (
            O => \N__3074\,
            I => \D_LM_040_in_6\
        );

    \I__484\ : InMux
    port map (
            O => \N__3071\,
            I => \N__3068\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__3068\,
            I => \N__3065\
        );

    \I__482\ : Span4Mux_v
    port map (
            O => \N__3065\,
            I => \N__3062\
        );

    \I__481\ : Span4Mux_h
    port map (
            O => \N__3062\,
            I => \N__3059\
        );

    \I__480\ : Sp12to4
    port map (
            O => \N__3059\,
            I => \N__3056\
        );

    \I__479\ : Span12Mux_h
    port map (
            O => \N__3056\,
            I => \N__3053\
        );

    \I__478\ : Odrv12
    port map (
            O => \N__3053\,
            I => \D_UU_040_in_6\
        );

    \I__477\ : IoInMux
    port map (
            O => \N__3050\,
            I => \N__3047\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3047\,
            I => \N__3044\
        );

    \I__475\ : IoSpan4Mux
    port map (
            O => \N__3044\,
            I => \N__3041\
        );

    \I__474\ : IoSpan4Mux
    port map (
            O => \N__3041\,
            I => \N__3038\
        );

    \I__473\ : Span4Mux_s3_v
    port map (
            O => \N__3038\,
            I => \N__3035\
        );

    \I__472\ : Odrv4
    port map (
            O => \N__3035\,
            I => \un1_D_UU_040_6\
        );

    \I__471\ : InMux
    port map (
            O => \N__3032\,
            I => \N__3029\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3029\,
            I => \N__3026\
        );

    \I__469\ : Span4Mux_v
    port map (
            O => \N__3026\,
            I => \N__3023\
        );

    \I__468\ : Sp12to4
    port map (
            O => \N__3023\,
            I => \N__3020\
        );

    \I__467\ : Odrv12
    port map (
            O => \N__3020\,
            I => \D_LL_AMIGA_in_3\
        );

    \I__466\ : IoInMux
    port map (
            O => \N__3017\,
            I => \N__3014\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3014\,
            I => \N__3011\
        );

    \I__464\ : IoSpan4Mux
    port map (
            O => \N__3011\,
            I => \N__3008\
        );

    \I__463\ : Sp12to4
    port map (
            O => \N__3008\,
            I => \N__3005\
        );

    \I__462\ : Span12Mux_s7_v
    port map (
            O => \N__3005\,
            I => \N__3002\
        );

    \I__461\ : Span12Mux_h
    port map (
            O => \N__3002\,
            I => \N__2999\
        );

    \I__460\ : Odrv12
    port map (
            O => \N__2999\,
            I => \un1_D_LL_AMIGA_3\
        );

    \I__459\ : IoInMux
    port map (
            O => \N__2996\,
            I => \N__2993\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__2993\,
            I => \N__2990\
        );

    \I__457\ : IoSpan4Mux
    port map (
            O => \N__2990\,
            I => \N__2987\
        );

    \I__456\ : Sp12to4
    port map (
            O => \N__2987\,
            I => \N__2984\
        );

    \I__455\ : Span12Mux_s7_h
    port map (
            O => \N__2984\,
            I => \N__2981\
        );

    \I__454\ : Span12Mux_h
    port map (
            O => \N__2981\,
            I => \N__2978\
        );

    \I__453\ : Odrv12
    port map (
            O => \N__2978\,
            I => \un1_D_UM_AMIGA_0\
        );

    \I__452\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2972\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__2972\,
            I => \N__2969\
        );

    \I__450\ : Span4Mux_v
    port map (
            O => \N__2969\,
            I => \N__2965\
        );

    \I__449\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2962\
        );

    \I__448\ : Span4Mux_v
    port map (
            O => \N__2965\,
            I => \N__2959\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2962\,
            I => \N__2956\
        );

    \I__446\ : Span4Mux_v
    port map (
            O => \N__2959\,
            I => \N__2952\
        );

    \I__445\ : Span4Mux_v
    port map (
            O => \N__2956\,
            I => \N__2949\
        );

    \I__444\ : InMux
    port map (
            O => \N__2955\,
            I => \N__2946\
        );

    \I__443\ : Sp12to4
    port map (
            O => \N__2952\,
            I => \N__2939\
        );

    \I__442\ : Sp12to4
    port map (
            O => \N__2949\,
            I => \N__2939\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__2946\,
            I => \N__2939\
        );

    \I__440\ : Span12Mux_h
    port map (
            O => \N__2939\,
            I => \N__2936\
        );

    \I__439\ : Odrv12
    port map (
            O => \N__2936\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__438\ : InMux
    port map (
            O => \N__2933\,
            I => \N__2930\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2930\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__436\ : InMux
    port map (
            O => \N__2927\,
            I => \N__2924\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2924\,
            I => \N__2921\
        );

    \I__434\ : Sp12to4
    port map (
            O => \N__2921\,
            I => \N__2918\
        );

    \I__433\ : Span12Mux_v
    port map (
            O => \N__2918\,
            I => \N__2915\
        );

    \I__432\ : Span12Mux_h
    port map (
            O => \N__2915\,
            I => \N__2912\
        );

    \I__431\ : Odrv12
    port map (
            O => \N__2912\,
            I => \D_UM_040_in_1\
        );

    \I__430\ : InMux
    port map (
            O => \N__2909\,
            I => \N__2906\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2906\,
            I => \N__2902\
        );

    \I__428\ : IoInMux
    port map (
            O => \N__2905\,
            I => \N__2899\
        );

    \I__427\ : Span4Mux_v
    port map (
            O => \N__2902\,
            I => \N__2896\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2899\,
            I => \N__2893\
        );

    \I__425\ : Span4Mux_v
    port map (
            O => \N__2896\,
            I => \N__2890\
        );

    \I__424\ : Span4Mux_s3_h
    port map (
            O => \N__2893\,
            I => \N__2887\
        );

    \I__423\ : Sp12to4
    port map (
            O => \N__2890\,
            I => \N__2884\
        );

    \I__422\ : Sp12to4
    port map (
            O => \N__2887\,
            I => \N__2881\
        );

    \I__421\ : Span12Mux_h
    port map (
            O => \N__2884\,
            I => \N__2878\
        );

    \I__420\ : Span12Mux_v
    port map (
            O => \N__2881\,
            I => \N__2875\
        );

    \I__419\ : Span12Mux_v
    port map (
            O => \N__2878\,
            I => \N__2872\
        );

    \I__418\ : Span12Mux_h
    port map (
            O => \N__2875\,
            I => \N__2869\
        );

    \I__417\ : Span12Mux_h
    port map (
            O => \N__2872\,
            I => \N__2866\
        );

    \I__416\ : Span12Mux_h
    port map (
            O => \N__2869\,
            I => \N__2863\
        );

    \I__415\ : Odrv12
    port map (
            O => \N__2866\,
            I => \D_LL_040_in_1\
        );

    \I__414\ : Odrv12
    port map (
            O => \N__2863\,
            I => \D_LL_040_in_1\
        );

    \I__413\ : IoInMux
    port map (
            O => \N__2858\,
            I => \N__2855\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2855\,
            I => \N__2852\
        );

    \I__411\ : IoSpan4Mux
    port map (
            O => \N__2852\,
            I => \N__2849\
        );

    \I__410\ : Span4Mux_s1_h
    port map (
            O => \N__2849\,
            I => \N__2846\
        );

    \I__409\ : Span4Mux_h
    port map (
            O => \N__2846\,
            I => \N__2843\
        );

    \I__408\ : Odrv4
    port map (
            O => \N__2843\,
            I => \un1_D_UM_040_1\
        );

    \I__407\ : IoInMux
    port map (
            O => \N__2840\,
            I => \N__2829\
        );

    \I__406\ : IoInMux
    port map (
            O => \N__2839\,
            I => \N__2826\
        );

    \I__405\ : IoInMux
    port map (
            O => \N__2838\,
            I => \N__2823\
        );

    \I__404\ : IoInMux
    port map (
            O => \N__2837\,
            I => \N__2815\
        );

    \I__403\ : IoInMux
    port map (
            O => \N__2836\,
            I => \N__2812\
        );

    \I__402\ : IoInMux
    port map (
            O => \N__2835\,
            I => \N__2809\
        );

    \I__401\ : IoInMux
    port map (
            O => \N__2834\,
            I => \N__2806\
        );

    \I__400\ : IoInMux
    port map (
            O => \N__2833\,
            I => \N__2803\
        );

    \I__399\ : IoInMux
    port map (
            O => \N__2832\,
            I => \N__2800\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2829\,
            I => \N__2797\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2826\,
            I => \N__2792\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2823\,
            I => \N__2792\
        );

    \I__395\ : IoInMux
    port map (
            O => \N__2822\,
            I => \N__2789\
        );

    \I__394\ : IoInMux
    port map (
            O => \N__2821\,
            I => \N__2786\
        );

    \I__393\ : IoInMux
    port map (
            O => \N__2820\,
            I => \N__2775\
        );

    \I__392\ : IoInMux
    port map (
            O => \N__2819\,
            I => \N__2772\
        );

    \I__391\ : IoInMux
    port map (
            O => \N__2818\,
            I => \N__2769\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__2815\,
            I => \N__2756\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2812\,
            I => \N__2756\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__2809\,
            I => \N__2756\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2806\,
            I => \N__2756\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2803\,
            I => \N__2756\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2800\,
            I => \N__2756\
        );

    \I__384\ : IoSpan4Mux
    port map (
            O => \N__2797\,
            I => \N__2747\
        );

    \I__383\ : IoSpan4Mux
    port map (
            O => \N__2792\,
            I => \N__2747\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__2789\,
            I => \N__2747\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2786\,
            I => \N__2747\
        );

    \I__380\ : IoInMux
    port map (
            O => \N__2785\,
            I => \N__2744\
        );

    \I__379\ : IoInMux
    port map (
            O => \N__2784\,
            I => \N__2741\
        );

    \I__378\ : IoInMux
    port map (
            O => \N__2783\,
            I => \N__2738\
        );

    \I__377\ : IoInMux
    port map (
            O => \N__2782\,
            I => \N__2735\
        );

    \I__376\ : IoInMux
    port map (
            O => \N__2781\,
            I => \N__2732\
        );

    \I__375\ : IoInMux
    port map (
            O => \N__2780\,
            I => \N__2729\
        );

    \I__374\ : IoInMux
    port map (
            O => \N__2779\,
            I => \N__2726\
        );

    \I__373\ : IoInMux
    port map (
            O => \N__2778\,
            I => \N__2723\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__2775\,
            I => \N__2714\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2772\,
            I => \N__2714\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2769\,
            I => \N__2714\
        );

    \I__369\ : IoSpan4Mux
    port map (
            O => \N__2756\,
            I => \N__2714\
        );

    \I__368\ : IoSpan4Mux
    port map (
            O => \N__2747\,
            I => \N__2699\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2744\,
            I => \N__2699\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2741\,
            I => \N__2699\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__2738\,
            I => \N__2699\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2735\,
            I => \N__2699\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__2732\,
            I => \N__2688\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2729\,
            I => \N__2688\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2726\,
            I => \N__2688\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__2723\,
            I => \N__2688\
        );

    \I__359\ : IoSpan4Mux
    port map (
            O => \N__2714\,
            I => \N__2688\
        );

    \I__358\ : IoInMux
    port map (
            O => \N__2713\,
            I => \N__2685\
        );

    \I__357\ : IoInMux
    port map (
            O => \N__2712\,
            I => \N__2682\
        );

    \I__356\ : IoInMux
    port map (
            O => \N__2711\,
            I => \N__2679\
        );

    \I__355\ : IoInMux
    port map (
            O => \N__2710\,
            I => \N__2676\
        );

    \I__354\ : IoSpan4Mux
    port map (
            O => \N__2699\,
            I => \N__2668\
        );

    \I__353\ : IoSpan4Mux
    port map (
            O => \N__2688\,
            I => \N__2657\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2685\,
            I => \N__2657\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2682\,
            I => \N__2657\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2679\,
            I => \N__2657\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2676\,
            I => \N__2657\
        );

    \I__348\ : IoInMux
    port map (
            O => \N__2675\,
            I => \N__2654\
        );

    \I__347\ : IoInMux
    port map (
            O => \N__2674\,
            I => \N__2651\
        );

    \I__346\ : IoInMux
    port map (
            O => \N__2673\,
            I => \N__2648\
        );

    \I__345\ : IoInMux
    port map (
            O => \N__2672\,
            I => \N__2645\
        );

    \I__344\ : IoInMux
    port map (
            O => \N__2671\,
            I => \N__2642\
        );

    \I__343\ : Span4Mux_s0_h
    port map (
            O => \N__2668\,
            I => \N__2639\
        );

    \I__342\ : IoSpan4Mux
    port map (
            O => \N__2657\,
            I => \N__2628\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2654\,
            I => \N__2628\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2651\,
            I => \N__2628\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2648\,
            I => \N__2628\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2645\,
            I => \N__2628\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2642\,
            I => \N__2625\
        );

    \I__336\ : Span4Mux_v
    port map (
            O => \N__2639\,
            I => \N__2618\
        );

    \I__335\ : IoSpan4Mux
    port map (
            O => \N__2628\,
            I => \N__2618\
        );

    \I__334\ : IoSpan4Mux
    port map (
            O => \N__2625\,
            I => \N__2618\
        );

    \I__333\ : Span4Mux_s0_h
    port map (
            O => \N__2618\,
            I => \N__2614\
        );

    \I__332\ : IoInMux
    port map (
            O => \N__2617\,
            I => \N__2611\
        );

    \I__331\ : Sp12to4
    port map (
            O => \N__2614\,
            I => \N__2606\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2611\,
            I => \N__2606\
        );

    \I__329\ : Odrv12
    port map (
            O => \N__2606\,
            I => \RnW_c_i_0\
        );

    \I__328\ : InMux
    port map (
            O => \N__2603\,
            I => \N__2600\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2600\,
            I => \N__2597\
        );

    \I__326\ : Span4Mux_v
    port map (
            O => \N__2597\,
            I => \N__2594\
        );

    \I__325\ : Sp12to4
    port map (
            O => \N__2594\,
            I => \N__2591\
        );

    \I__324\ : Odrv12
    port map (
            O => \N__2591\,
            I => \D_LM_AMIGA_in_4\
        );

    \I__323\ : IoInMux
    port map (
            O => \N__2588\,
            I => \N__2585\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__2585\,
            I => \N__2582\
        );

    \I__321\ : IoSpan4Mux
    port map (
            O => \N__2582\,
            I => \N__2579\
        );

    \I__320\ : IoSpan4Mux
    port map (
            O => \N__2579\,
            I => \N__2576\
        );

    \I__319\ : Span4Mux_s3_h
    port map (
            O => \N__2576\,
            I => \N__2573\
        );

    \I__318\ : Sp12to4
    port map (
            O => \N__2573\,
            I => \N__2570\
        );

    \I__317\ : Span12Mux_s11_h
    port map (
            O => \N__2570\,
            I => \N__2567\
        );

    \I__316\ : Odrv12
    port map (
            O => \N__2567\,
            I => \un1_D_LM_AMIGA_4\
        );

    \I__315\ : InMux
    port map (
            O => \N__2564\,
            I => \N__2561\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2561\,
            I => \N__2558\
        );

    \I__313\ : Span4Mux_v
    port map (
            O => \N__2558\,
            I => \N__2555\
        );

    \I__312\ : Sp12to4
    port map (
            O => \N__2555\,
            I => \N__2552\
        );

    \I__311\ : Odrv12
    port map (
            O => \N__2552\,
            I => \D_LM_AMIGA_in_5\
        );

    \I__310\ : IoInMux
    port map (
            O => \N__2549\,
            I => \N__2546\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2546\,
            I => \N__2543\
        );

    \I__308\ : Span4Mux_s3_h
    port map (
            O => \N__2543\,
            I => \N__2540\
        );

    \I__307\ : Sp12to4
    port map (
            O => \N__2540\,
            I => \N__2537\
        );

    \I__306\ : Span12Mux_v
    port map (
            O => \N__2537\,
            I => \N__2534\
        );

    \I__305\ : Span12Mux_h
    port map (
            O => \N__2534\,
            I => \N__2531\
        );

    \I__304\ : Odrv12
    port map (
            O => \N__2531\,
            I => \un1_D_LM_AMIGA_5\
        );

    \I__303\ : InMux
    port map (
            O => \N__2528\,
            I => \N__2525\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2525\,
            I => \N__2522\
        );

    \I__301\ : Span12Mux_v
    port map (
            O => \N__2522\,
            I => \N__2519\
        );

    \I__300\ : Odrv12
    port map (
            O => \N__2519\,
            I => \D_LM_AMIGA_in_6\
        );

    \I__299\ : IoInMux
    port map (
            O => \N__2516\,
            I => \N__2513\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2513\,
            I => \N__2510\
        );

    \I__297\ : IoSpan4Mux
    port map (
            O => \N__2510\,
            I => \N__2507\
        );

    \I__296\ : Span4Mux_s3_h
    port map (
            O => \N__2507\,
            I => \N__2504\
        );

    \I__295\ : Span4Mux_h
    port map (
            O => \N__2504\,
            I => \N__2501\
        );

    \I__294\ : Span4Mux_h
    port map (
            O => \N__2501\,
            I => \N__2498\
        );

    \I__293\ : Sp12to4
    port map (
            O => \N__2498\,
            I => \N__2495\
        );

    \I__292\ : Odrv12
    port map (
            O => \N__2495\,
            I => \un1_D_LM_AMIGA_6\
        );

    \I__291\ : InMux
    port map (
            O => \N__2492\,
            I => \N__2489\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2489\,
            I => \N__2486\
        );

    \I__289\ : Span4Mux_v
    port map (
            O => \N__2486\,
            I => \N__2483\
        );

    \I__288\ : Sp12to4
    port map (
            O => \N__2483\,
            I => \N__2480\
        );

    \I__287\ : Span12Mux_h
    port map (
            O => \N__2480\,
            I => \N__2477\
        );

    \I__286\ : Span12Mux_h
    port map (
            O => \N__2477\,
            I => \N__2474\
        );

    \I__285\ : Odrv12
    port map (
            O => \N__2474\,
            I => \D_UU_040_in_3\
        );

    \I__284\ : IoInMux
    port map (
            O => \N__2471\,
            I => \N__2468\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2468\,
            I => \N__2465\
        );

    \I__282\ : IoSpan4Mux
    port map (
            O => \N__2465\,
            I => \N__2462\
        );

    \I__281\ : IoSpan4Mux
    port map (
            O => \N__2462\,
            I => \N__2458\
        );

    \I__280\ : InMux
    port map (
            O => \N__2461\,
            I => \N__2455\
        );

    \I__279\ : Span4Mux_s2_h
    port map (
            O => \N__2458\,
            I => \N__2452\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2455\,
            I => \N__2449\
        );

    \I__277\ : Sp12to4
    port map (
            O => \N__2452\,
            I => \N__2446\
        );

    \I__276\ : Span12Mux_s10_v
    port map (
            O => \N__2449\,
            I => \N__2443\
        );

    \I__275\ : Span12Mux_h
    port map (
            O => \N__2446\,
            I => \N__2440\
        );

    \I__274\ : Span12Mux_v
    port map (
            O => \N__2443\,
            I => \N__2437\
        );

    \I__273\ : Span12Mux_h
    port map (
            O => \N__2440\,
            I => \N__2434\
        );

    \I__272\ : Span12Mux_h
    port map (
            O => \N__2437\,
            I => \N__2431\
        );

    \I__271\ : Odrv12
    port map (
            O => \N__2434\,
            I => \D_LM_040_in_3\
        );

    \I__270\ : Odrv12
    port map (
            O => \N__2431\,
            I => \D_LM_040_in_3\
        );

    \I__269\ : IoInMux
    port map (
            O => \N__2426\,
            I => \N__2423\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2423\,
            I => \N__2420\
        );

    \I__267\ : IoSpan4Mux
    port map (
            O => \N__2420\,
            I => \N__2417\
        );

    \I__266\ : Span4Mux_s3_v
    port map (
            O => \N__2417\,
            I => \N__2414\
        );

    \I__265\ : Span4Mux_h
    port map (
            O => \N__2414\,
            I => \N__2411\
        );

    \I__264\ : Odrv4
    port map (
            O => \N__2411\,
            I => \un1_D_UU_040_3\
        );

    \I__263\ : InMux
    port map (
            O => \N__2408\,
            I => \N__2405\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__2405\,
            I => \N__2402\
        );

    \I__261\ : Span4Mux_v
    port map (
            O => \N__2402\,
            I => \N__2399\
        );

    \I__260\ : Sp12to4
    port map (
            O => \N__2399\,
            I => \N__2396\
        );

    \I__259\ : Odrv12
    port map (
            O => \N__2396\,
            I => \D_LL_AMIGA_in_0\
        );

    \I__258\ : IoInMux
    port map (
            O => \N__2393\,
            I => \N__2390\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2390\,
            I => \N__2387\
        );

    \I__256\ : Span12Mux_s9_h
    port map (
            O => \N__2387\,
            I => \N__2384\
        );

    \I__255\ : Span12Mux_h
    port map (
            O => \N__2384\,
            I => \N__2381\
        );

    \I__254\ : Odrv12
    port map (
            O => \N__2381\,
            I => \un1_D_LL_AMIGA_0\
        );

    \I__253\ : InMux
    port map (
            O => \N__2378\,
            I => \N__2375\
        );

    \I__252\ : LocalMux
    port map (
            O => \N__2375\,
            I => \N__2372\
        );

    \I__251\ : Span4Mux_v
    port map (
            O => \N__2372\,
            I => \N__2369\
        );

    \I__250\ : Sp12to4
    port map (
            O => \N__2369\,
            I => \N__2366\
        );

    \I__249\ : Odrv12
    port map (
            O => \N__2366\,
            I => \D_LL_AMIGA_in_1\
        );

    \I__248\ : IoInMux
    port map (
            O => \N__2363\,
            I => \N__2360\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__2360\,
            I => \N__2357\
        );

    \I__246\ : IoSpan4Mux
    port map (
            O => \N__2357\,
            I => \N__2354\
        );

    \I__245\ : IoSpan4Mux
    port map (
            O => \N__2354\,
            I => \N__2351\
        );

    \I__244\ : Span4Mux_s2_h
    port map (
            O => \N__2351\,
            I => \N__2348\
        );

    \I__243\ : Sp12to4
    port map (
            O => \N__2348\,
            I => \N__2345\
        );

    \I__242\ : Span12Mux_s9_h
    port map (
            O => \N__2345\,
            I => \N__2342\
        );

    \I__241\ : Span12Mux_h
    port map (
            O => \N__2342\,
            I => \N__2339\
        );

    \I__240\ : Odrv12
    port map (
            O => \N__2339\,
            I => \un1_D_LL_AMIGA_1\
        );

    \I__239\ : InMux
    port map (
            O => \N__2336\,
            I => \N__2333\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2333\,
            I => \N__2330\
        );

    \I__237\ : Span12Mux_h
    port map (
            O => \N__2330\,
            I => \N__2327\
        );

    \I__236\ : Odrv12
    port map (
            O => \N__2327\,
            I => \D_LM_AMIGA_in_3\
        );

    \I__235\ : IoInMux
    port map (
            O => \N__2324\,
            I => \N__2321\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2321\,
            I => \N__2318\
        );

    \I__233\ : IoSpan4Mux
    port map (
            O => \N__2318\,
            I => \N__2315\
        );

    \I__232\ : IoSpan4Mux
    port map (
            O => \N__2315\,
            I => \N__2312\
        );

    \I__231\ : Span4Mux_s0_h
    port map (
            O => \N__2312\,
            I => \N__2309\
        );

    \I__230\ : Sp12to4
    port map (
            O => \N__2309\,
            I => \N__2306\
        );

    \I__229\ : Span12Mux_h
    port map (
            O => \N__2306\,
            I => \N__2303\
        );

    \I__228\ : Odrv12
    port map (
            O => \N__2303\,
            I => \un1_D_LM_AMIGA_3\
        );

    \I__227\ : InMux
    port map (
            O => \N__2300\,
            I => \N__2297\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__2297\,
            I => \N__2294\
        );

    \I__225\ : Span12Mux_h
    port map (
            O => \N__2294\,
            I => \N__2291\
        );

    \I__224\ : Odrv12
    port map (
            O => \N__2291\,
            I => \A_040_c_1\
        );

    \I__223\ : InMux
    port map (
            O => \N__2288\,
            I => \N__2285\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__2285\,
            I => \N__2282\
        );

    \I__221\ : Span4Mux_h
    port map (
            O => \N__2282\,
            I => \N__2279\
        );

    \I__220\ : Span4Mux_v
    port map (
            O => \N__2279\,
            I => \N__2276\
        );

    \I__219\ : Odrv4
    port map (
            O => \N__2276\,
            I => \A_040_c_0\
        );

    \I__218\ : IoInMux
    port map (
            O => \N__2273\,
            I => \N__2270\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__2270\,
            I => \N__2267\
        );

    \I__216\ : Span4Mux_s2_v
    port map (
            O => \N__2267\,
            I => \N__2264\
        );

    \I__215\ : Span4Mux_v
    port map (
            O => \N__2264\,
            I => \N__2261\
        );

    \I__214\ : Odrv4
    port map (
            O => \N__2261\,
            I => \A_AMIGA_c_0\
        );

    \I__213\ : InMux
    port map (
            O => \N__2258\,
            I => \N__2255\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__2255\,
            I => \N__2252\
        );

    \I__211\ : Span4Mux_v
    port map (
            O => \N__2252\,
            I => \N__2249\
        );

    \I__210\ : Sp12to4
    port map (
            O => \N__2249\,
            I => \N__2246\
        );

    \I__209\ : Odrv12
    port map (
            O => \N__2246\,
            I => \D_LL_AMIGA_in_2\
        );

    \I__208\ : IoInMux
    port map (
            O => \N__2243\,
            I => \N__2240\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__2240\,
            I => \N__2237\
        );

    \I__206\ : Span4Mux_s3_h
    port map (
            O => \N__2237\,
            I => \N__2234\
        );

    \I__205\ : Sp12to4
    port map (
            O => \N__2234\,
            I => \N__2231\
        );

    \I__204\ : Span12Mux_s8_v
    port map (
            O => \N__2231\,
            I => \N__2228\
        );

    \I__203\ : Span12Mux_h
    port map (
            O => \N__2228\,
            I => \N__2225\
        );

    \I__202\ : Odrv12
    port map (
            O => \N__2225\,
            I => \un1_D_LL_AMIGA_2\
        );

    \I__201\ : InMux
    port map (
            O => \N__2222\,
            I => \N__2219\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__2219\,
            I => \N__2216\
        );

    \I__199\ : Odrv12
    port map (
            O => \N__2216\,
            I => \D_LM_AMIGA_in_2\
        );

    \I__198\ : IoInMux
    port map (
            O => \N__2213\,
            I => \N__2210\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__2210\,
            I => \N__2207\
        );

    \I__196\ : Sp12to4
    port map (
            O => \N__2207\,
            I => \N__2204\
        );

    \I__195\ : Span12Mux_h
    port map (
            O => \N__2204\,
            I => \N__2201\
        );

    \I__194\ : Span12Mux_v
    port map (
            O => \N__2201\,
            I => \N__2198\
        );

    \I__193\ : Odrv12
    port map (
            O => \N__2198\,
            I => \un1_D_LM_AMIGA_2\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            I => \N__6959\
        );

    \INVU111_CYCLE_SM.CYCLE_STATE_1C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\,
            I => \N__6964\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            I => \N__6967\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net\,
            I => \N__6963\
        );

    \INVU111_CYCLE_SM.CYCLE_STATE_0C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.CYCLE_STATE_0C_net\,
            I => \N__6966\
        );

    \INVU111_CYCLE_SM.A_OUTC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.A_OUTC_net\,
            I => \N__6969\
        );

    \INVU111_CYCLE_SM.TSnC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TSnC_net\,
            I => \N__5562\
        );

    \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\,
            I => \N__6965\
        );

    \INVU111_CYCLE_SM.TA_EN_nessC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TA_EN_nessC_net\,
            I => \N__6968\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net\,
            I => \N__6970\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3644\,
            in1 => \N__2300\,
            in2 => \_gnd_net_\,
            in3 => \N__5512\,
            lcout => \A_AMIGA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__2288\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5513\,
            lcout => \A_AMIGA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4797\,
            in1 => \N__2258\,
            in2 => \_gnd_net_\,
            in3 => \N__6327\,
            lcout => \un1_D_LL_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6316\,
            in1 => \N__5701\,
            in2 => \_gnd_net_\,
            in3 => \N__2222\,
            lcout => \un1_D_LM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6328\,
            in1 => \N__2927\,
            in2 => \_gnd_net_\,
            in3 => \N__2909\,
            lcout => \un1_D_UM_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RnW_c_sbtinv_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4001\,
            lcout => \RnW_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2603\,
            in1 => \N__6297\,
            in2 => \_gnd_net_\,
            in3 => \N__3412\,
            lcout => \un1_D_LM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2564\,
            in1 => \N__6299\,
            in2 => \_gnd_net_\,
            in3 => \N__5755\,
            lcout => \un1_D_LM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3477\,
            in1 => \N__6329\,
            in2 => \_gnd_net_\,
            in3 => \N__2528\,
            lcout => \un1_D_LM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2492\,
            in1 => \N__6361\,
            in2 => \_gnd_net_\,
            in3 => \N__2461\,
            lcout => \un1_D_UU_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2408\,
            in1 => \N__6326\,
            in2 => \_gnd_net_\,
            in3 => \N__2975\,
            lcout => \un1_D_LL_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2378\,
            in1 => \N__6289\,
            in2 => \_gnd_net_\,
            in3 => \N__4568\,
            lcout => \un1_D_LL_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2336\,
            in1 => \N__6249\,
            in2 => \_gnd_net_\,
            in3 => \N__5933\,
            lcout => \un1_D_LM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3245\,
            in1 => \N__6298\,
            in2 => \_gnd_net_\,
            in3 => \N__3336\,
            lcout => \un1_D_LM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIM3VM1_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__3209\,
            in1 => \N__6410\,
            in2 => \_gnd_net_\,
            in3 => \N__5500\,
            lcout => \U111_CYCLE_SM.FLIP\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4702\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3188\,
            in1 => \N__6279\,
            in2 => \_gnd_net_\,
            in3 => \N__3166\,
            lcout => \un1_D_UM_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3106\,
            in1 => \N__6280\,
            in2 => \_gnd_net_\,
            in3 => \N__3071\,
            lcout => \un1_D_UU_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3032\,
            in1 => \N__6269\,
            in2 => \_gnd_net_\,
            in3 => \N__5144\,
            lcout => \un1_D_LL_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__2933\,
            in1 => \N__2968\,
            in2 => \_gnd_net_\,
            in3 => \N__5416\,
            lcout => \un1_D_UM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2955\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net\,
            ce => \N__5231\,
            sr => \N__5193\
        );

    \U111_CYCLE_SM.TA_EN_ness_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5285\,
            lcout => \U111_CYCLE_SM.TA_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TA_EN_nessC_net\,
            ce => \N__3593\,
            sr => \N__3607\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3416\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\,
            ce => \N__5232\,
            sr => \N__5189\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3347\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\,
            ce => \N__5232\,
            sr => \N__5189\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3491\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_4C_net\,
            ce => \N__5232\,
            sr => \N__5189\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3581\,
            in1 => \N__6317\,
            in2 => \_gnd_net_\,
            in3 => \N__3530\,
            lcout => \un1_D_UU_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3490\,
            in1 => \N__3458\,
            in2 => \_gnd_net_\,
            in3 => \N__5485\,
            lcout => \un1_D_UU_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__5484\,
            in1 => \N__3425\,
            in2 => \_gnd_net_\,
            in3 => \N__3402\,
            lcout => \un1_D_UU_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__5502\,
            in1 => \N__3356\,
            in2 => \_gnd_net_\,
            in3 => \N__3346\,
            lcout => \un1_D_UU_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_10_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4423\,
            in1 => \N__6290\,
            in2 => \_gnd_net_\,
            in3 => \N__3284\,
            lcout => \un1_D_LL_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4190\,
            in1 => \N__6170\,
            in2 => \_gnd_net_\,
            in3 => \N__3719\,
            lcout => \un1_D_LM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6247\,
            in1 => \N__4499\,
            in2 => \_gnd_net_\,
            in3 => \N__3680\,
            lcout => \un1_D_LM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TSn_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4738\,
            in2 => \_gnd_net_\,
            in3 => \N__4075\,
            lcout => \TSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TSnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__3631\,
            in1 => \N__3617\,
            in2 => \N__4752\,
            in3 => \N__5279\,
            lcout => \U111_CYCLE_SM.A_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.A_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100100000"
        )
    port map (
            in0 => \N__5277\,
            in1 => \N__4668\,
            in2 => \N__4616\,
            in3 => \N__4039\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.LW_CYCLE_r_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100011001000"
        )
    port map (
            in0 => \N__5409\,
            in1 => \N__4742\,
            in2 => \N__3620\,
            in3 => \N__5278\,
            lcout => \U111_CYCLE_SM.LW_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.A_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_0_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__5276\,
            in1 => \_gnd_net_\,
            in2 => \N__4615\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.TS_EN10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_RNIIU7U_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__5408\,
            in1 => \N__4605\,
            in2 => \N__4040\,
            in3 => \N__5275\,
            lcout => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0\,
            ltout => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_ness_RNO_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3611\,
            in3 => \N__3608\,
            lcout => \U111_CYCLE_SM.un1_CYCLE_STATE_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__5240\,
            in1 => \N__4085\,
            in2 => \N__4079\,
            in3 => \N__4746\,
            lcout => \U111_CYCLE_SM.TS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.A_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6403\,
            in1 => \N__4051\,
            in2 => \N__4753\,
            in3 => \N__6442\,
            lcout => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.A_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_0_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__5274\,
            in1 => \N__4669\,
            in2 => \N__4614\,
            in3 => \N__4747\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.CYCLE_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4670\,
            in1 => \N__5273\,
            in2 => \_gnd_net_\,
            in3 => \N__4601\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111111"
        )
    port map (
            in0 => \N__3943\,
            in1 => \_gnd_net_\,
            in2 => \N__3731\,
            in3 => \N__4748\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3728\,
            in3 => \N__3725\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4424\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net\,
            ce => \N__5230\,
            sr => \N__5188\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4564\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net\,
            ce => \N__5230\,
            sr => \N__5188\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4495\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net\,
            ce => \N__5230\,
            sr => \N__5188\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4183\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net\,
            ce => \N__5230\,
            sr => \N__5188\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4574\,
            in1 => \N__5444\,
            in2 => \_gnd_net_\,
            in3 => \N__4557\,
            lcout => \un1_D_UM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4488\,
            in1 => \N__4463\,
            in2 => \_gnd_net_\,
            in3 => \N__5476\,
            lcout => \un1_D_UU_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__5477\,
            in1 => \N__4433\,
            in2 => \_gnd_net_\,
            in3 => \N__4419\,
            lcout => \un1_D_UM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6366\,
            in1 => \N__4352\,
            in2 => \_gnd_net_\,
            in3 => \N__4327\,
            lcout => \un1_D_UU_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__4274\,
            in1 => \N__6365\,
            in2 => \_gnd_net_\,
            in3 => \N__4255\,
            lcout => \un1_D_UU_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4202\,
            in1 => \N__4171\,
            in2 => \_gnd_net_\,
            in3 => \N__5501\,
            lcout => \un1_D_UU_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6234\,
            in1 => \N__5360\,
            in2 => \_gnd_net_\,
            in3 => \N__4127\,
            lcout => \un1_D_LL_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5642\,
            in1 => \N__6233\,
            in2 => \_gnd_net_\,
            in3 => \N__4973\,
            lcout => \un1_D_LL_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5048\,
            in1 => \N__6232\,
            in2 => \_gnd_net_\,
            in3 => \N__4934\,
            lcout => \un1_D_LL_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6248\,
            in1 => \N__4892\,
            in2 => \_gnd_net_\,
            in3 => \N__4873\,
            lcout => \un1_D_UM_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4799\,
            in1 => \N__4760\,
            in2 => \_gnd_net_\,
            in3 => \N__5417\,
            lcout => \un1_D_UM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5346\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            ce => \N__5233\,
            sr => \N__5194\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4798\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            ce => \N__5233\,
            sr => \N__5194\
        );

    \U111_CYCLE_SM.CYCLE_STATE_1_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001000010100000"
        )
    port map (
            in0 => \N__5281\,
            in1 => \N__4666\,
            in2 => \N__4754\,
            in3 => \N__4613\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_ness_RNIPNOD_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4679\,
            in2 => \_gnd_net_\,
            in3 => \N__4667\,
            lcout => \TAn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_1_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000010"
        )
    port map (
            in0 => \N__5569\,
            in1 => \N__4612\,
            in2 => \N__5303\,
            in3 => \N__5280\,
            lcout => \U111_CYCLE_SM.TS_EN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5140\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__5234\,
            sr => \N__5195\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5705\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__5234\,
            sr => \N__5195\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5047\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__5234\,
            sr => \N__5195\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5635\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__5234\,
            sr => \N__5195\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5774\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__5234\,
            sr => \N__5195\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5926\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__5234\,
            sr => \N__5195\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5139\,
            in1 => \N__5087\,
            in2 => \_gnd_net_\,
            in3 => \N__5486\,
            lcout => \un1_D_UM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__5487\,
            in1 => \N__5057\,
            in2 => \_gnd_net_\,
            in3 => \N__5040\,
            lcout => \un1_D_UM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6035\,
            in1 => \N__6368\,
            in2 => \_gnd_net_\,
            in3 => \N__5984\,
            lcout => \un1_D_UM_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__5505\,
            in1 => \N__5942\,
            in2 => \_gnd_net_\,
            in3 => \N__5925\,
            lcout => \un1_D_UU_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6367\,
            in1 => \N__5870\,
            in2 => \_gnd_net_\,
            in3 => \N__5845\,
            lcout => \un1_D_UM_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5786\,
            in1 => \N__5767\,
            in2 => \_gnd_net_\,
            in3 => \N__5506\,
            lcout => \un1_D_UU_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__5504\,
            in1 => \N__5714\,
            in2 => \_gnd_net_\,
            in3 => \N__5697\,
            lcout => \un1_D_UU_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5623\,
            in1 => \N__5600\,
            in2 => \_gnd_net_\,
            in3 => \N__5503\,
            lcout => \un1_D_UM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5570\,
            lcout => \GB_BUFFER_CLK40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__5440\,
            in1 => \N__5366\,
            in2 => \_gnd_net_\,
            in3 => \N__5353\,
            lcout => \un1_D_UM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6974\,
            lcout => \GB_BUFFER_CLK80_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6871\,
            in1 => \N__6362\,
            in2 => \_gnd_net_\,
            in3 => \N__6830\,
            lcout => \un1_D_UU_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6363\,
            in1 => \N__6787\,
            in2 => \_gnd_net_\,
            in3 => \N__6752\,
            lcout => \un1_D_UU_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6314\,
            in1 => \N__6719\,
            in2 => \_gnd_net_\,
            in3 => \N__6703\,
            lcout => \un1_D_UM_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6640\,
            in1 => \N__6315\,
            in2 => \_gnd_net_\,
            in3 => \N__6599\,
            lcout => \un1_D_UM_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6566\,
            in1 => \N__6341\,
            in2 => \_gnd_net_\,
            in3 => \N__6521\,
            lcout => \un1_D_UM_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_TRANS_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__6482\,
            in1 => \N__6464\,
            in2 => \_gnd_net_\,
            in3 => \N__6446\,
            lcout => \U111_CYCLE_SM.LW_TRANS_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6386\,
            in1 => \N__6364\,
            in2 => \_gnd_net_\,
            in3 => \N__6085\,
            lcout => \un1_D_UU_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

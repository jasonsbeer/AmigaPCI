-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 20 2025 20:31:24

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    TM : in std_logic_vector(1 downto 0);
    TT : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(31 downto 1);
    CIACS1n : out std_logic;
    TICK50 : out std_logic;
    RAMSPACEn : out std_logic;
    TICK60 : out std_logic;
    CIACS0n : out std_logic;
    CLK6 : in std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    REGSPACEn : out std_logic;
    CLK_CIA : out std_logic;
    BUFENn : out std_logic;
    TSn : in std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    TACKn : inout std_logic;
    ROMENn : out std_logic;
    PORTSIZE : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__7109\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3123\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2907\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2677\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_17\ : std_logic;
signal \A_c_31\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_25\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_3\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_28\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_27\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_TRANSFER_ACK.N_41_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3Z0Z_2\ : std_logic;
signal \U409_CIA_PORTSIZE_i_a2_0_3\ : std_logic;
signal \A_c_19\ : std_logic;
signal \A_c_18\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \A_c_26\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_11_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_17\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_4\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_11\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_14\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_10\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_17\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_16\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\ : std_logic;
signal \TM_c_0\ : std_logic;
signal \TM_c_1\ : std_logic;
signal \PORTSIZE_i_a2\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_12\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\ : std_logic;
signal \U409_CIA.N_89\ : std_logic;
signal \A_c_22\ : std_logic;
signal \OVL_c\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3Z0Z_4_cascade_\ : std_logic;
signal \N_53_i\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.N_54_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_5_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a3_0_1_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a3_0_1_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_54_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0Z0Z_0\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3Z0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.N_16_i\ : std_logic;
signal \un1_RAMSPACEn_i_i_a3_cascade_\ : std_logic;
signal \N_11_i\ : std_logic;
signal \un1_RAMSPACEn_i_i_a3\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \un1_REGSPACEn_i_i_a3_0_a2_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \N_90\ : std_logic;
signal \A_c_21\ : std_logic;
signal \N_80\ : std_logic;
signal \N_52_i\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_EN_iC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en\ : std_logic;
signal \ROMENn_c\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROMENnC_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \N_76\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_EN_e_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_28_4\ : std_logic;
signal \U409_TRANSFER_ACK.N_28_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_64\ : std_logic;
signal \U409_TRANSFER_ACK.N_63_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.m9_i_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_45\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_73\ : std_logic;
signal \U409_TRANSFER_ACK.N_60\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_65\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_68\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_23\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \CIA_ENABLE\ : std_logic;
signal \CIA_ENABLE_cascade_\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_0C_net\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U409_CIA.N_93_cascade_\ : std_logic;
signal \U409_CIA.VMA_RNOZ0Z_1_cascade_\ : std_logic;
signal \U409_CIA.VMA_3_0_a2_2\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \U409_CIA.N_91_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2\ : std_logic;
signal \U409_CIA.N_91\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_2_1\ : std_logic;
signal \U409_CIA.CLK_CIA_r_1_cascade_\ : std_logic;
signal \U409_CIA.CLK_CIA6_1_0\ : std_logic;
signal \CLK_CIA_c\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \bfn_13_2_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \bfn_13_3_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \U409_CIA.CLK_CIA6_1\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_6\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_6\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_7\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \U409_TICK.TICK603_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \bfn_15_1_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \bfn_15_2_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \TACK_EN_i\ : std_logic;
signal \N_525_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \TM_wire\ : std_logic_vector(1 downto 0);
signal \CLK_CIA_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    \TT_wire\ <= TT;
    \A_wire\ <= A;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    \TM_wire\ <= TM;
    CLK_CIA <= \CLK_CIA_wire\;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    \TSn_wire\ <= TSn;
    BUFENn <= \BUFENn_wire\;
    PORTSIZE <= \PORTSIZE_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TICK60 <= \TICK60_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__4804\,
            RESETB => \N__5026\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__7107\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7109\,
            DIN => \N__7108\,
            DOUT => \N__7107\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7109\,
            PADOUT => \N__7108\,
            PADIN => \N__7107\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__7097\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7099\,
            DIN => \N__7098\,
            DOUT => \N__7097\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7099\,
            PADOUT => \N__7098\,
            PADIN => \N__7097\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7088\,
            DIN => \N__7087\,
            DOUT => \N__7086\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7088\,
            PADOUT => \N__7087\,
            PADIN => \N__7086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7079\,
            DIN => \N__7078\,
            DOUT => \N__7077\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7079\,
            PADOUT => \N__7078\,
            PADIN => \N__7077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7070\,
            DIN => \N__7069\,
            DOUT => \N__7068\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7070\,
            PADOUT => \N__7069\,
            PADIN => \N__7068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7061\,
            DIN => \N__7060\,
            DOUT => \N__7059\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7061\,
            PADOUT => \N__7060\,
            PADIN => \N__7059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4993\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7052\,
            DIN => \N__7051\,
            DOUT => \N__7050\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7052\,
            PADOUT => \N__7051\,
            PADIN => \N__7050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4249\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7043\,
            DIN => \N__7042\,
            DOUT => \N__7041\,
            PACKAGEPIN => \TM_wire\(1)
        );

    \TM_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7043\,
            PADOUT => \N__7042\,
            PADIN => \N__7041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7034\,
            DIN => \N__7033\,
            DOUT => \N__7032\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7034\,
            PADOUT => \N__7033\,
            PADIN => \N__7032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_CIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7025\,
            DIN => \N__7024\,
            DOUT => \N__7023\,
            PACKAGEPIN => \CLK_CIA_wire\
        );

    \CLK_CIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7025\,
            PADOUT => \N__7024\,
            PADIN => \N__7023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5440\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7016\,
            DIN => \N__7015\,
            DOUT => \N__7014\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7016\,
            PADOUT => \N__7015\,
            PADIN => \N__7014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7007\,
            DIN => \N__7006\,
            DOUT => \N__7005\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7007\,
            PADOUT => \N__7006\,
            PADIN => \N__7005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3388\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6998\,
            DIN => \N__6997\,
            DOUT => \N__6996\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6998\,
            PADOUT => \N__6997\,
            PADIN => \N__6996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6643\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__3661\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6989\,
            DIN => \N__6988\,
            DOUT => \N__6987\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6989\,
            PADOUT => \N__6988\,
            PADIN => \N__6987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6980\,
            DIN => \N__6979\,
            DOUT => \N__6978\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6980\,
            PADOUT => \N__6979\,
            PADIN => \N__6978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4150\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6971\,
            DIN => \N__6970\,
            DOUT => \N__6969\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6971\,
            PADOUT => \N__6970\,
            PADIN => \N__6969\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6962\,
            DIN => \N__6961\,
            DOUT => \N__6960\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6962\,
            PADOUT => \N__6961\,
            PADIN => \N__6960\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6953\,
            DIN => \N__6952\,
            DOUT => \N__6951\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6953\,
            PADOUT => \N__6952\,
            PADIN => \N__6951\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3712\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6944\,
            DIN => \N__6943\,
            DOUT => \N__6942\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6944\,
            PADOUT => \N__6943\,
            PADIN => \N__6942\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3295\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6935\,
            DIN => \N__6934\,
            DOUT => \N__6933\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6935\,
            PADOUT => \N__6934\,
            PADIN => \N__6933\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6926\,
            DIN => \N__6925\,
            DOUT => \N__6924\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6926\,
            PADOUT => \N__6925\,
            PADIN => \N__6924\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6917\,
            DIN => \N__6916\,
            DOUT => \N__6915\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6917\,
            PADOUT => \N__6916\,
            PADIN => \N__6915\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6908\,
            DIN => \N__6907\,
            DOUT => \N__6906\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6908\,
            PADOUT => \N__6907\,
            PADIN => \N__6906\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6899\,
            DIN => \N__6898\,
            DOUT => \N__6897\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6899\,
            PADOUT => \N__6898\,
            PADIN => \N__6897\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6890\,
            DIN => \N__6889\,
            DOUT => \N__6888\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6890\,
            PADOUT => \N__6889\,
            PADIN => \N__6888\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6881\,
            DIN => \N__6880\,
            DOUT => \N__6879\,
            PACKAGEPIN => \TM_wire\(0)
        );

    \TM_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6881\,
            PADOUT => \N__6880\,
            PADIN => \N__6879\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6872\,
            DIN => \N__6871\,
            DOUT => \N__6870\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6872\,
            PADOUT => \N__6871\,
            PADIN => \N__6870\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6863\,
            DIN => \N__6862\,
            DOUT => \N__6861\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6863\,
            PADOUT => \N__6862\,
            PADIN => \N__6861\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6854\,
            DIN => \N__6853\,
            DOUT => \N__6852\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6854\,
            PADOUT => \N__6853\,
            PADIN => \N__6852\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6845\,
            DIN => \N__6844\,
            DOUT => \N__6843\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6845\,
            PADOUT => \N__6844\,
            PADIN => \N__6843\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4948\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6836\,
            DIN => \N__6835\,
            DOUT => \N__6834\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6836\,
            PADOUT => \N__6835\,
            PADIN => \N__6834\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5533\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6827\,
            DIN => \N__6826\,
            DOUT => \N__6825\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6827\,
            PADOUT => \N__6826\,
            PADIN => \N__6825\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6818\,
            DIN => \N__6817\,
            DOUT => \N__6816\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6818\,
            PADOUT => \N__6817\,
            PADIN => \N__6816\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6809\,
            DIN => \N__6808\,
            DOUT => \N__6807\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6809\,
            PADOUT => \N__6808\,
            PADIN => \N__6807\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6800\,
            DIN => \N__6799\,
            DOUT => \N__6798\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6800\,
            PADOUT => \N__6799\,
            PADIN => \N__6798\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6791\,
            DIN => \N__6790\,
            DOUT => \N__6789\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6791\,
            PADOUT => \N__6790\,
            PADIN => \N__6789\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6782\,
            DIN => \N__6781\,
            DOUT => \N__6780\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6782\,
            PADOUT => \N__6781\,
            PADIN => \N__6780\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5899\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6773\,
            DIN => \N__6772\,
            DOUT => \N__6771\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6773\,
            PADOUT => \N__6772\,
            PADIN => \N__6771\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6764\,
            DIN => \N__6763\,
            DOUT => \N__6762\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6764\,
            PADOUT => \N__6763\,
            PADIN => \N__6762\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1592\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6741\
        );

    \I__1591\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6738\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__6741\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__6738\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__6733\,
            I => \N__6730\
        );

    \I__1587\ : InMux
    port map (
            O => \N__6730\,
            I => \N__6727\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__6727\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__1585\ : InMux
    port map (
            O => \N__6724\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__1584\ : InMux
    port map (
            O => \N__6721\,
            I => \N__6717\
        );

    \I__1583\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6714\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__6717\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__6714\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__1580\ : InMux
    port map (
            O => \N__6709\,
            I => \N__6706\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__6706\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__1578\ : InMux
    port map (
            O => \N__6703\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__1577\ : InMux
    port map (
            O => \N__6700\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__1576\ : InMux
    port map (
            O => \N__6697\,
            I => \N__6693\
        );

    \I__1575\ : InMux
    port map (
            O => \N__6696\,
            I => \N__6690\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__6693\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__6690\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__1572\ : ClkMux
    port map (
            O => \N__6685\,
            I => \N__6661\
        );

    \I__1571\ : ClkMux
    port map (
            O => \N__6684\,
            I => \N__6661\
        );

    \I__1570\ : ClkMux
    port map (
            O => \N__6683\,
            I => \N__6661\
        );

    \I__1569\ : ClkMux
    port map (
            O => \N__6682\,
            I => \N__6661\
        );

    \I__1568\ : ClkMux
    port map (
            O => \N__6681\,
            I => \N__6661\
        );

    \I__1567\ : ClkMux
    port map (
            O => \N__6680\,
            I => \N__6661\
        );

    \I__1566\ : ClkMux
    port map (
            O => \N__6679\,
            I => \N__6661\
        );

    \I__1565\ : ClkMux
    port map (
            O => \N__6678\,
            I => \N__6661\
        );

    \I__1564\ : GlobalMux
    port map (
            O => \N__6661\,
            I => \N__6658\
        );

    \I__1563\ : gio2CtrlBuf
    port map (
            O => \N__6658\,
            I => \CLK6_c_g\
        );

    \I__1562\ : InMux
    port map (
            O => \N__6655\,
            I => \N__6652\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__6652\,
            I => \N__6649\
        );

    \I__1560\ : Span12Mux_v
    port map (
            O => \N__6649\,
            I => \N__6646\
        );

    \I__1559\ : Odrv12
    port map (
            O => \N__6646\,
            I => \TACK_EN_i\
        );

    \I__1558\ : IoInMux
    port map (
            O => \N__6643\,
            I => \N__6640\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__6640\,
            I => \N__6637\
        );

    \I__1556\ : IoSpan4Mux
    port map (
            O => \N__6637\,
            I => \N__6634\
        );

    \I__1555\ : Span4Mux_s3_v
    port map (
            O => \N__6634\,
            I => \N__6631\
        );

    \I__1554\ : Span4Mux_v
    port map (
            O => \N__6631\,
            I => \N__6628\
        );

    \I__1553\ : Span4Mux_v
    port map (
            O => \N__6628\,
            I => \N__6625\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__6625\,
            I => \N_525_i\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__6622\,
            I => \N__6618\
        );

    \I__1550\ : InMux
    port map (
            O => \N__6621\,
            I => \N__6615\
        );

    \I__1549\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6612\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__6615\,
            I => \N__6609\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__6612\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__6609\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__1545\ : InMux
    port map (
            O => \N__6604\,
            I => \N__6601\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__6601\,
            I => \N__6598\
        );

    \I__1543\ : Odrv4
    port map (
            O => \N__6598\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__1542\ : InMux
    port map (
            O => \N__6595\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__1541\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6588\
        );

    \I__1540\ : InMux
    port map (
            O => \N__6591\,
            I => \N__6585\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__6588\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__6585\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__1537\ : InMux
    port map (
            O => \N__6580\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__1536\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6573\
        );

    \I__1535\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6570\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__6573\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__6570\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__1532\ : InMux
    port map (
            O => \N__6565\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__1531\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6559\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__6559\,
            I => \N__6555\
        );

    \I__1529\ : InMux
    port map (
            O => \N__6558\,
            I => \N__6552\
        );

    \I__1528\ : Odrv4
    port map (
            O => \N__6555\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__6552\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__1526\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6544\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__6544\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__1524\ : InMux
    port map (
            O => \N__6541\,
            I => \bfn_15_2_0_\
        );

    \I__1523\ : InMux
    port map (
            O => \N__6538\,
            I => \N__6535\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__6535\,
            I => \N__6532\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__6532\,
            I => \N__6528\
        );

    \I__1520\ : InMux
    port map (
            O => \N__6531\,
            I => \N__6525\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__6528\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__6525\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__1517\ : InMux
    port map (
            O => \N__6520\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__1516\ : InMux
    port map (
            O => \N__6517\,
            I => \N__6513\
        );

    \I__1515\ : InMux
    port map (
            O => \N__6516\,
            I => \N__6510\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__6513\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__6510\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__1512\ : InMux
    port map (
            O => \N__6505\,
            I => \N__6502\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__6502\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__1510\ : InMux
    port map (
            O => \N__6499\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__1509\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6493\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__6493\,
            I => \N__6490\
        );

    \I__1507\ : Span4Mux_h
    port map (
            O => \N__6490\,
            I => \N__6486\
        );

    \I__1506\ : InMux
    port map (
            O => \N__6489\,
            I => \N__6483\
        );

    \I__1505\ : Odrv4
    port map (
            O => \N__6486\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__6483\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__1503\ : InMux
    port map (
            O => \N__6478\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__1502\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6471\
        );

    \I__1501\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6468\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__6471\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__6468\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__1498\ : CascadeMux
    port map (
            O => \N__6463\,
            I => \N__6460\
        );

    \I__1497\ : InMux
    port map (
            O => \N__6460\,
            I => \N__6457\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__6457\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__1495\ : InMux
    port map (
            O => \N__6454\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__1494\ : InMux
    port map (
            O => \N__6451\,
            I => \N__6447\
        );

    \I__1493\ : InMux
    port map (
            O => \N__6450\,
            I => \N__6444\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__6447\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__6444\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__1490\ : InMux
    port map (
            O => \N__6439\,
            I => \N__6436\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__6436\,
            I => \N__6432\
        );

    \I__1488\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6429\
        );

    \I__1487\ : Odrv4
    port map (
            O => \N__6432\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__6429\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__6424\,
            I => \N__6421\
        );

    \I__1484\ : InMux
    port map (
            O => \N__6421\,
            I => \N__6417\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__6420\,
            I => \N__6414\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__6417\,
            I => \N__6411\
        );

    \I__1481\ : InMux
    port map (
            O => \N__6414\,
            I => \N__6408\
        );

    \I__1480\ : Odrv4
    port map (
            O => \N__6411\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__6408\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__1478\ : InMux
    port map (
            O => \N__6403\,
            I => \N__6399\
        );

    \I__1477\ : InMux
    port map (
            O => \N__6402\,
            I => \N__6396\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__6399\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__6396\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__1474\ : CascadeMux
    port map (
            O => \N__6391\,
            I => \N__6382\
        );

    \I__1473\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6379\
        );

    \I__1472\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6372\
        );

    \I__1471\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6372\
        );

    \I__1470\ : InMux
    port map (
            O => \N__6387\,
            I => \N__6372\
        );

    \I__1469\ : InMux
    port map (
            O => \N__6386\,
            I => \N__6365\
        );

    \I__1468\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6365\
        );

    \I__1467\ : InMux
    port map (
            O => \N__6382\,
            I => \N__6365\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__6379\,
            I => \N__6362\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__6372\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__6365\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__6362\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__6355\,
            I => \N__6352\
        );

    \I__1461\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6343\
        );

    \I__1460\ : InMux
    port map (
            O => \N__6351\,
            I => \N__6340\
        );

    \I__1459\ : InMux
    port map (
            O => \N__6350\,
            I => \N__6337\
        );

    \I__1458\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6328\
        );

    \I__1457\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6328\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6347\,
            I => \N__6328\
        );

    \I__1455\ : InMux
    port map (
            O => \N__6346\,
            I => \N__6328\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__6343\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__6340\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__6337\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__6328\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__6319\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__1449\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__6313\,
            I => \N__6308\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__6312\,
            I => \N__6304\
        );

    \I__1446\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6301\
        );

    \I__1445\ : Span4Mux_h
    port map (
            O => \N__6308\,
            I => \N__6298\
        );

    \I__1444\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6295\
        );

    \I__1443\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6292\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__6301\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1441\ : Odrv4
    port map (
            O => \N__6298\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__6295\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__6292\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1438\ : InMux
    port map (
            O => \N__6283\,
            I => \N__6279\
        );

    \I__1437\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6276\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__6279\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__6276\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6271\,
            I => \N__6267\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6264\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__6267\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__6264\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__6259\,
            I => \N__6256\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6256\,
            I => \N__6253\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__6253\,
            I => \N__6249\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6252\,
            I => \N__6246\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__6249\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__6246\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1424\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6237\
        );

    \I__1423\ : InMux
    port map (
            O => \N__6240\,
            I => \N__6234\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__6237\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__6234\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6229\,
            I => \N__6219\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6228\,
            I => \N__6212\
        );

    \I__1418\ : InMux
    port map (
            O => \N__6227\,
            I => \N__6212\
        );

    \I__1417\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6212\
        );

    \I__1416\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6203\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6224\,
            I => \N__6203\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6223\,
            I => \N__6203\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6222\,
            I => \N__6203\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6219\,
            I => \N__6200\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6212\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__6203\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1409\ : Odrv4
    port map (
            O => \N__6200\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1408\ : CascadeMux
    port map (
            O => \N__6193\,
            I => \N__6189\
        );

    \I__1407\ : InMux
    port map (
            O => \N__6192\,
            I => \N__6183\
        );

    \I__1406\ : InMux
    port map (
            O => \N__6189\,
            I => \N__6183\
        );

    \I__1405\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6180\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__6183\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__6180\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__6175\,
            I => \N__6171\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__6174\,
            I => \N__6166\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6161\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6161\
        );

    \I__1398\ : InMux
    port map (
            O => \N__6169\,
            I => \N__6158\
        );

    \I__1397\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6155\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__6161\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__6158\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6155\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__1393\ : InMux
    port map (
            O => \N__6148\,
            I => \N__6144\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6141\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6144\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6141\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__1389\ : InMux
    port map (
            O => \N__6136\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__1388\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6130\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__6130\,
            I => \N__6126\
        );

    \I__1386\ : InMux
    port map (
            O => \N__6129\,
            I => \N__6123\
        );

    \I__1385\ : Odrv4
    port map (
            O => \N__6126\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__6123\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6118\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__6115\,
            I => \N__6112\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6112\,
            I => \N__6108\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6105\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6108\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6105\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6100\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6093\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6096\,
            I => \N__6090\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__6093\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__6090\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__1372\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6082\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6082\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__1370\ : InMux
    port map (
            O => \N__6079\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6072\
        );

    \I__1368\ : InMux
    port map (
            O => \N__6075\,
            I => \N__6069\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__6072\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__6069\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6064\,
            I => \N__6060\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6063\,
            I => \N__6057\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__6060\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__6057\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__1361\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6049\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__6049\,
            I => \U409_TICK.TICK603_11\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__6046\,
            I => \U409_TICK.TICK603_8_cascade_\
        );

    \I__1358\ : InMux
    port map (
            O => \N__6043\,
            I => \N__6039\
        );

    \I__1357\ : InMux
    port map (
            O => \N__6042\,
            I => \N__6036\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__6039\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__6036\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__6031\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__1353\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6025\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__6025\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6022\,
            I => \N__6018\
        );

    \I__1350\ : InMux
    port map (
            O => \N__6021\,
            I => \N__6015\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6018\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__6015\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6010\,
            I => \N__5998\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6009\,
            I => \N__5998\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6008\,
            I => \N__5993\
        );

    \I__1344\ : InMux
    port map (
            O => \N__6007\,
            I => \N__5993\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6006\,
            I => \N__5984\
        );

    \I__1342\ : InMux
    port map (
            O => \N__6005\,
            I => \N__5984\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6004\,
            I => \N__5984\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6003\,
            I => \N__5984\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__5998\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__5993\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__5984\,
            I => \U409_TICK.TICK503_10\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__5977\,
            I => \N__5973\
        );

    \I__1335\ : InMux
    port map (
            O => \N__5976\,
            I => \N__5964\
        );

    \I__1334\ : InMux
    port map (
            O => \N__5973\,
            I => \N__5961\
        );

    \I__1333\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5958\
        );

    \I__1332\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5947\
        );

    \I__1331\ : InMux
    port map (
            O => \N__5970\,
            I => \N__5947\
        );

    \I__1330\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5947\
        );

    \I__1329\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5947\
        );

    \I__1328\ : InMux
    port map (
            O => \N__5967\,
            I => \N__5947\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__5964\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__5961\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__5958\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__5947\,
            I => \U409_TICK.TICK503_14\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__5938\,
            I => \N__5931\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__5937\,
            I => \N__5928\
        );

    \I__1321\ : InMux
    port map (
            O => \N__5936\,
            I => \N__5920\
        );

    \I__1320\ : InMux
    port map (
            O => \N__5935\,
            I => \N__5920\
        );

    \I__1319\ : InMux
    port map (
            O => \N__5934\,
            I => \N__5909\
        );

    \I__1318\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5909\
        );

    \I__1317\ : InMux
    port map (
            O => \N__5928\,
            I => \N__5909\
        );

    \I__1316\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5909\
        );

    \I__1315\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5909\
        );

    \I__1314\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5906\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5920\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__5909\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__5906\,
            I => \U409_TICK.TICK503_9\
        );

    \I__1310\ : IoInMux
    port map (
            O => \N__5899\,
            I => \N__5896\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__5896\,
            I => \N__5893\
        );

    \I__1308\ : IoSpan4Mux
    port map (
            O => \N__5893\,
            I => \N__5890\
        );

    \I__1307\ : Span4Mux_s3_v
    port map (
            O => \N__5890\,
            I => \N__5887\
        );

    \I__1306\ : Span4Mux_v
    port map (
            O => \N__5887\,
            I => \N__5883\
        );

    \I__1305\ : InMux
    port map (
            O => \N__5886\,
            I => \N__5880\
        );

    \I__1304\ : Odrv4
    port map (
            O => \N__5883\,
            I => \TICK60_c\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__5880\,
            I => \TICK60_c\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__5875\,
            I => \N__5872\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5869\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__5869\,
            I => \N__5866\
        );

    \I__1299\ : Odrv4
    port map (
            O => \N__5866\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5863\,
            I => \N__5860\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__5860\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__5857\,
            I => \N__5854\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5854\,
            I => \N__5851\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__5851\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5848\,
            I => \N__5845\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5845\,
            I => \U409_TICK.TICK503_11\
        );

    \I__1291\ : CascadeMux
    port map (
            O => \N__5842\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5835\
        );

    \I__1289\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5832\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__5835\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5832\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5827\,
            I => \N__5823\
        );

    \I__1285\ : InMux
    port map (
            O => \N__5826\,
            I => \N__5820\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__5823\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__5820\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__5815\,
            I => \N__5811\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5814\,
            I => \N__5807\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5811\,
            I => \N__5804\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5810\,
            I => \N__5801\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5807\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5804\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__5801\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1275\ : InMux
    port map (
            O => \N__5794\,
            I => \N__5790\
        );

    \I__1274\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5787\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__5790\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__5787\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__5782\,
            I => \N__5779\
        );

    \I__1270\ : InMux
    port map (
            O => \N__5779\,
            I => \N__5776\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__5776\,
            I => \N__5773\
        );

    \I__1268\ : Odrv4
    port map (
            O => \N__5773\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5765\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5769\,
            I => \N__5760\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5768\,
            I => \N__5760\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5765\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5760\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1262\ : InMux
    port map (
            O => \N__5755\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__1261\ : InMux
    port map (
            O => \N__5752\,
            I => \N__5747\
        );

    \I__1260\ : InMux
    port map (
            O => \N__5751\,
            I => \N__5742\
        );

    \I__1259\ : InMux
    port map (
            O => \N__5750\,
            I => \N__5742\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__5747\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5742\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5737\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5727\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5724\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5732\,
            I => \N__5717\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5717\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5730\,
            I => \N__5717\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5727\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5724\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5717\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5710\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5707\,
            I => \N__5701\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5701\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5701\,
            I => \U409_CIA.CIA_CLK_COUNT11\
        );

    \I__1243\ : InMux
    port map (
            O => \N__5698\,
            I => \N__5693\
        );

    \I__1242\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5688\
        );

    \I__1241\ : InMux
    port map (
            O => \N__5696\,
            I => \N__5688\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__5693\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__5688\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5683\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5680\,
            I => \N__5675\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5679\,
            I => \N__5672\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5669\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5675\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__5672\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__5669\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5662\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\
        );

    \I__1230\ : InMux
    port map (
            O => \N__5659\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__5656\,
            I => \N__5652\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5655\,
            I => \N__5648\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5652\,
            I => \N__5645\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5642\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__5648\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5645\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5642\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__5635\,
            I => \N__5628\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5622\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5633\,
            I => \N__5622\
        );

    \I__1219\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5619\
        );

    \I__1218\ : InMux
    port map (
            O => \N__5631\,
            I => \N__5612\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5612\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5627\,
            I => \N__5612\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__5622\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__5619\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5612\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1212\ : ClkMux
    port map (
            O => \N__5605\,
            I => \N__5596\
        );

    \I__1211\ : ClkMux
    port map (
            O => \N__5604\,
            I => \N__5596\
        );

    \I__1210\ : ClkMux
    port map (
            O => \N__5603\,
            I => \N__5596\
        );

    \I__1209\ : GlobalMux
    port map (
            O => \N__5596\,
            I => \N__5593\
        );

    \I__1208\ : gio2CtrlBuf
    port map (
            O => \N__5593\,
            I => \CLK28_IN_c_g\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5590\,
            I => \bfn_13_3_0_\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5587\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5584\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5581\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5578\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5575\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5572\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5569\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5559\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5565\,
            I => \N__5552\
        );

    \I__1197\ : InMux
    port map (
            O => \N__5564\,
            I => \N__5552\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5552\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5549\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5559\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5552\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5549\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5542\,
            I => \N__5539\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__5539\,
            I => \U409_CIA.CLK_CIA6_1\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__5536\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__1188\ : IoInMux
    port map (
            O => \N__5533\,
            I => \N__5530\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5530\,
            I => \N__5527\
        );

    \I__1186\ : Span4Mux_s2_v
    port map (
            O => \N__5527\,
            I => \N__5524\
        );

    \I__1185\ : Span4Mux_v
    port map (
            O => \N__5524\,
            I => \N__5521\
        );

    \I__1184\ : Span4Mux_h
    port map (
            O => \N__5521\,
            I => \N__5517\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5514\
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__5517\,
            I => \TICK50_c\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5514\,
            I => \TICK50_c\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5509\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5506\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5503\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5500\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5497\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5494\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__5491\,
            I => \N__5488\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5485\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__5485\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5482\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5479\,
            I => \N__5476\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__5476\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5473\,
            I => \N__5469\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5472\,
            I => \N__5466\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5469\,
            I => \U409_CIA.N_91\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5466\,
            I => \U409_CIA.N_91\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5458\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5458\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_2_1\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__5455\,
            I => \U409_CIA.CLK_CIA_r_1_cascade_\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5452\,
            I => \N__5448\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5451\,
            I => \N__5445\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5448\,
            I => \U409_CIA.CLK_CIA6_1_0\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5445\,
            I => \U409_CIA.CLK_CIA6_1_0\
        );

    \I__1157\ : IoInMux
    port map (
            O => \N__5440\,
            I => \N__5437\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5437\,
            I => \N__5434\
        );

    \I__1155\ : Span4Mux_s2_v
    port map (
            O => \N__5434\,
            I => \N__5431\
        );

    \I__1154\ : Span4Mux_h
    port map (
            O => \N__5431\,
            I => \N__5428\
        );

    \I__1153\ : Span4Mux_v
    port map (
            O => \N__5428\,
            I => \N__5423\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5427\,
            I => \N__5420\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__5426\,
            I => \N__5416\
        );

    \I__1150\ : Sp12to4
    port map (
            O => \N__5423\,
            I => \N__5411\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5420\,
            I => \N__5411\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5419\,
            I => \N__5406\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5416\,
            I => \N__5406\
        );

    \I__1146\ : Odrv12
    port map (
            O => \N__5411\,
            I => \CLK_CIA_c\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5406\,
            I => \CLK_CIA_c\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__5401\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__5398\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5388\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5394\,
            I => \N__5385\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5378\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5392\,
            I => \N__5378\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5391\,
            I => \N__5378\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5388\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__5385\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5378\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__5368\,
            I => \N__5359\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5367\,
            I => \N__5356\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5353\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5350\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__5364\,
            I => \N__5345\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__5363\,
            I => \N__5342\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__5362\,
            I => \N__5339\
        );

    \I__1126\ : Span4Mux_h
    port map (
            O => \N__5359\,
            I => \N__5334\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__5356\,
            I => \N__5334\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5353\,
            I => \N__5329\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__5350\,
            I => \N__5329\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5326\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5319\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5319\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5319\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5316\
        );

    \I__1117\ : Span4Mux_v
    port map (
            O => \N__5334\,
            I => \N__5312\
        );

    \I__1116\ : Span4Mux_h
    port map (
            O => \N__5329\,
            I => \N__5309\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__5326\,
            I => \N__5302\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__5319\,
            I => \N__5302\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__5316\,
            I => \N__5302\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__5315\,
            I => \N__5298\
        );

    \I__1111\ : Span4Mux_h
    port map (
            O => \N__5312\,
            I => \N__5290\
        );

    \I__1110\ : Span4Mux_v
    port map (
            O => \N__5309\,
            I => \N__5290\
        );

    \I__1109\ : Span4Mux_h
    port map (
            O => \N__5302\,
            I => \N__5290\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5301\,
            I => \N__5287\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5298\,
            I => \N__5282\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5297\,
            I => \N__5282\
        );

    \I__1105\ : Span4Mux_v
    port map (
            O => \N__5290\,
            I => \N__5277\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5287\,
            I => \N__5274\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5282\,
            I => \N__5271\
        );

    \I__1102\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5268\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5280\,
            I => \N__5265\
        );

    \I__1100\ : Sp12to4
    port map (
            O => \N__5277\,
            I => \N__5254\
        );

    \I__1099\ : Span12Mux_v
    port map (
            O => \N__5274\,
            I => \N__5254\
        );

    \I__1098\ : Sp12to4
    port map (
            O => \N__5271\,
            I => \N__5254\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5268\,
            I => \N__5254\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5265\,
            I => \N__5254\
        );

    \I__1095\ : Span12Mux_v
    port map (
            O => \N__5254\,
            I => \N__5251\
        );

    \I__1094\ : Span12Mux_h
    port map (
            O => \N__5251\,
            I => \N__5248\
        );

    \I__1093\ : Odrv12
    port map (
            O => \N__5248\,
            I => \RESETn_c\
        );

    \I__1092\ : SRMux
    port map (
            O => \N__5245\,
            I => \N__5240\
        );

    \I__1091\ : SRMux
    port map (
            O => \N__5244\,
            I => \N__5234\
        );

    \I__1090\ : SRMux
    port map (
            O => \N__5243\,
            I => \N__5231\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5240\,
            I => \N__5227\
        );

    \I__1088\ : SRMux
    port map (
            O => \N__5239\,
            I => \N__5224\
        );

    \I__1087\ : SRMux
    port map (
            O => \N__5238\,
            I => \N__5221\
        );

    \I__1086\ : SRMux
    port map (
            O => \N__5237\,
            I => \N__5218\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5234\,
            I => \N__5215\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__5231\,
            I => \N__5212\
        );

    \I__1083\ : SRMux
    port map (
            O => \N__5230\,
            I => \N__5209\
        );

    \I__1082\ : Span4Mux_h
    port map (
            O => \N__5227\,
            I => \N__5204\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__5224\,
            I => \N__5204\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__5221\,
            I => \N__5201\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5218\,
            I => \N__5196\
        );

    \I__1078\ : Span4Mux_h
    port map (
            O => \N__5215\,
            I => \N__5196\
        );

    \I__1077\ : Span4Mux_v
    port map (
            O => \N__5212\,
            I => \N__5193\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5209\,
            I => \N__5188\
        );

    \I__1075\ : Sp12to4
    port map (
            O => \N__5204\,
            I => \N__5188\
        );

    \I__1074\ : Span4Mux_v
    port map (
            O => \N__5201\,
            I => \N__5183\
        );

    \I__1073\ : Span4Mux_v
    port map (
            O => \N__5196\,
            I => \N__5183\
        );

    \I__1072\ : Odrv4
    port map (
            O => \N__5193\,
            I => \RESETn_c_i\
        );

    \I__1071\ : Odrv12
    port map (
            O => \N__5188\,
            I => \RESETn_c_i\
        );

    \I__1070\ : Odrv4
    port map (
            O => \N__5183\,
            I => \RESETn_c_i\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__5176\,
            I => \U409_CIA.N_93_cascade_\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__5173\,
            I => \U409_CIA.VMA_RNOZ0Z_1_cascade_\
        );

    \I__1067\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5167\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__1065\ : Span4Mux_v
    port map (
            O => \N__5164\,
            I => \N__5161\
        );

    \I__1064\ : Odrv4
    port map (
            O => \N__5161\,
            I => \U409_CIA.VMA_3_0_a2_2\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5154\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5151\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5154\,
            I => \N__5145\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__5151\,
            I => \N__5145\
        );

    \I__1059\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5142\
        );

    \I__1058\ : Odrv12
    port map (
            O => \N__5145\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__5142\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__5137\,
            I => \U409_CIA.N_91_cascade_\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5124\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5124\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5117\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5131\,
            I => \N__5117\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5130\,
            I => \N__5117\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5114\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5124\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5117\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5114\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__5107\,
            I => \N__5102\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__5106\,
            I => \N__5099\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__5105\,
            I => \N__5095\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5085\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5085\
        );

    \I__1041\ : InMux
    port map (
            O => \N__5098\,
            I => \N__5085\
        );

    \I__1040\ : InMux
    port map (
            O => \N__5095\,
            I => \N__5078\
        );

    \I__1039\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5078\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5093\,
            I => \N__5078\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5092\,
            I => \N__5075\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5085\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5078\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5075\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5068\,
            I => \N__5065\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5065\,
            I => \N__5056\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5064\,
            I => \N__5049\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5049\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5049\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5044\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5060\,
            I => \N__5044\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5059\,
            I => \N__5041\
        );

    \I__1025\ : Odrv4
    port map (
            O => \N__5056\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__5049\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5044\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__5041\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5032\,
            I => \N__5029\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5029\,
            I => \U409_TRANSFER_ACK.N_23\
        );

    \I__1019\ : IoInMux
    port map (
            O => \N__5026\,
            I => \N__5023\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5023\,
            I => \N__5020\
        );

    \I__1017\ : Span4Mux_s2_v
    port map (
            O => \N__5020\,
            I => \N__5017\
        );

    \I__1016\ : Span4Mux_v
    port map (
            O => \N__5017\,
            I => \N__5014\
        );

    \I__1015\ : Odrv4
    port map (
            O => \N__5014\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5011\,
            I => \N__5008\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5008\,
            I => \N__5005\
        );

    \I__1012\ : Span4Mux_v
    port map (
            O => \N__5005\,
            I => \N__5002\
        );

    \I__1011\ : Sp12to4
    port map (
            O => \N__5002\,
            I => \N__4999\
        );

    \I__1010\ : Span12Mux_h
    port map (
            O => \N__4999\,
            I => \N__4996\
        );

    \I__1009\ : Odrv12
    port map (
            O => \N__4996\,
            I => \A_c_13\
        );

    \I__1008\ : IoInMux
    port map (
            O => \N__4993\,
            I => \N__4990\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4990\,
            I => \N__4987\
        );

    \I__1006\ : IoSpan4Mux
    port map (
            O => \N__4987\,
            I => \N__4984\
        );

    \I__1005\ : Span4Mux_s2_h
    port map (
            O => \N__4984\,
            I => \N__4981\
        );

    \I__1004\ : Sp12to4
    port map (
            O => \N__4981\,
            I => \N__4978\
        );

    \I__1003\ : Span12Mux_h
    port map (
            O => \N__4978\,
            I => \N__4975\
        );

    \I__1002\ : Odrv12
    port map (
            O => \N__4975\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4969\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4969\,
            I => \CIA_ENABLE\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__4966\,
            I => \CIA_ENABLE_cascade_\
        );

    \I__998\ : InMux
    port map (
            O => \N__4963\,
            I => \N__4960\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__4960\,
            I => \N__4957\
        );

    \I__996\ : Span12Mux_s10_v
    port map (
            O => \N__4957\,
            I => \N__4954\
        );

    \I__995\ : Span12Mux_h
    port map (
            O => \N__4954\,
            I => \N__4951\
        );

    \I__994\ : Odrv12
    port map (
            O => \N__4951\,
            I => \A_c_12\
        );

    \I__993\ : IoInMux
    port map (
            O => \N__4948\,
            I => \N__4945\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__4945\,
            I => \N__4942\
        );

    \I__991\ : IoSpan4Mux
    port map (
            O => \N__4942\,
            I => \N__4939\
        );

    \I__990\ : IoSpan4Mux
    port map (
            O => \N__4939\,
            I => \N__4936\
        );

    \I__989\ : Sp12to4
    port map (
            O => \N__4936\,
            I => \N__4933\
        );

    \I__988\ : Span12Mux_s7_h
    port map (
            O => \N__4933\,
            I => \N__4930\
        );

    \I__987\ : Odrv12
    port map (
            O => \N__4930\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__986\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4922\
        );

    \I__985\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4917\
        );

    \I__984\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4917\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4922\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4917\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__4912\,
            I => \N__4909\
        );

    \I__980\ : InMux
    port map (
            O => \N__4909\,
            I => \N__4903\
        );

    \I__979\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4903\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4903\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__4900\,
            I => \N__4894\
        );

    \I__976\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4891\
        );

    \I__975\ : InMux
    port map (
            O => \N__4898\,
            I => \N__4884\
        );

    \I__974\ : InMux
    port map (
            O => \N__4897\,
            I => \N__4884\
        );

    \I__973\ : InMux
    port map (
            O => \N__4894\,
            I => \N__4884\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4891\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4884\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__970\ : InMux
    port map (
            O => \N__4879\,
            I => \N__4876\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4876\,
            I => \U409_TRANSFER_ACK.N_64\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__4873\,
            I => \U409_TRANSFER_ACK.N_63_cascade_\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__4870\,
            I => \U409_TRANSFER_ACK.m9_i_1_cascade_\
        );

    \I__966\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4861\
        );

    \I__965\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4861\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__4861\,
            I => \U409_TRANSFER_ACK.N_45\
        );

    \I__963\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4853\
        );

    \I__962\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4848\
        );

    \I__961\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4848\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4853\,
            I => \U409_TRANSFER_ACK.N_73\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4848\,
            I => \U409_TRANSFER_ACK.N_73\
        );

    \I__958\ : InMux
    port map (
            O => \N__4843\,
            I => \N__4840\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4840\,
            I => \U409_TRANSFER_ACK.N_60\
        );

    \I__956\ : InMux
    port map (
            O => \N__4837\,
            I => \N__4830\
        );

    \I__955\ : InMux
    port map (
            O => \N__4836\,
            I => \N__4821\
        );

    \I__954\ : InMux
    port map (
            O => \N__4835\,
            I => \N__4821\
        );

    \I__953\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4821\
        );

    \I__952\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4821\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4830\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__4821\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__949\ : CascadeMux
    port map (
            O => \N__4816\,
            I => \U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_\
        );

    \I__948\ : InMux
    port map (
            O => \N__4813\,
            I => \N__4810\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4810\,
            I => \U409_TRANSFER_ACK.N_65\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__4807\,
            I => \N__4800\
        );

    \I__945\ : CascadeMux
    port map (
            O => \N__4806\,
            I => \N__4797\
        );

    \I__944\ : CascadeMux
    port map (
            O => \N__4805\,
            I => \N__4794\
        );

    \I__943\ : IoInMux
    port map (
            O => \N__4804\,
            I => \N__4791\
        );

    \I__942\ : InMux
    port map (
            O => \N__4803\,
            I => \N__4788\
        );

    \I__941\ : InMux
    port map (
            O => \N__4800\,
            I => \N__4785\
        );

    \I__940\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4782\
        );

    \I__939\ : InMux
    port map (
            O => \N__4794\,
            I => \N__4779\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4791\,
            I => \N__4775\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4788\,
            I => \N__4770\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4785\,
            I => \N__4767\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4782\,
            I => \N__4764\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4779\,
            I => \N__4761\
        );

    \I__933\ : InMux
    port map (
            O => \N__4778\,
            I => \N__4758\
        );

    \I__932\ : IoSpan4Mux
    port map (
            O => \N__4775\,
            I => \N__4755\
        );

    \I__931\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4752\
        );

    \I__930\ : InMux
    port map (
            O => \N__4773\,
            I => \N__4749\
        );

    \I__929\ : Span4Mux_v
    port map (
            O => \N__4770\,
            I => \N__4744\
        );

    \I__928\ : Span4Mux_h
    port map (
            O => \N__4767\,
            I => \N__4744\
        );

    \I__927\ : Span4Mux_v
    port map (
            O => \N__4764\,
            I => \N__4737\
        );

    \I__926\ : Span4Mux_h
    port map (
            O => \N__4761\,
            I => \N__4737\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4758\,
            I => \N__4737\
        );

    \I__924\ : Span4Mux_s0_v
    port map (
            O => \N__4755\,
            I => \N__4734\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4752\,
            I => \N__4731\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__4749\,
            I => \N__4728\
        );

    \I__921\ : Span4Mux_v
    port map (
            O => \N__4744\,
            I => \N__4723\
        );

    \I__920\ : Span4Mux_h
    port map (
            O => \N__4737\,
            I => \N__4723\
        );

    \I__919\ : Sp12to4
    port map (
            O => \N__4734\,
            I => \N__4720\
        );

    \I__918\ : Span4Mux_h
    port map (
            O => \N__4731\,
            I => \N__4715\
        );

    \I__917\ : Span4Mux_h
    port map (
            O => \N__4728\,
            I => \N__4715\
        );

    \I__916\ : Span4Mux_v
    port map (
            O => \N__4723\,
            I => \N__4712\
        );

    \I__915\ : Span12Mux_v
    port map (
            O => \N__4720\,
            I => \N__4709\
        );

    \I__914\ : Sp12to4
    port map (
            O => \N__4715\,
            I => \N__4706\
        );

    \I__913\ : Span4Mux_v
    port map (
            O => \N__4712\,
            I => \N__4703\
        );

    \I__912\ : Span12Mux_v
    port map (
            O => \N__4709\,
            I => \N__4700\
        );

    \I__911\ : Span12Mux_v
    port map (
            O => \N__4706\,
            I => \N__4697\
        );

    \I__910\ : Span4Mux_v
    port map (
            O => \N__4703\,
            I => \N__4694\
        );

    \I__909\ : Odrv12
    port map (
            O => \N__4700\,
            I => \CLK40_IN_c\
        );

    \I__908\ : Odrv12
    port map (
            O => \N__4697\,
            I => \CLK40_IN_c\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__4694\,
            I => \CLK40_IN_c\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__4687\,
            I => \N__4682\
        );

    \I__905\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4676\
        );

    \I__904\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4673\
        );

    \I__903\ : InMux
    port map (
            O => \N__4682\,
            I => \N__4664\
        );

    \I__902\ : InMux
    port map (
            O => \N__4681\,
            I => \N__4664\
        );

    \I__901\ : InMux
    port map (
            O => \N__4680\,
            I => \N__4664\
        );

    \I__900\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4664\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4676\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4673\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4664\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__896\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4654\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4654\,
            I => \U409_TRANSFER_ACK.N_68\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__4651\,
            I => \N__4647\
        );

    \I__893\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4644\
        );

    \I__892\ : InMux
    port map (
            O => \N__4647\,
            I => \N__4641\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__4644\,
            I => \N__4638\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4641\,
            I => \N__4635\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__4638\,
            I => \N__4631\
        );

    \I__888\ : Span4Mux_v
    port map (
            O => \N__4635\,
            I => \N__4628\
        );

    \I__887\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4625\
        );

    \I__886\ : Sp12to4
    port map (
            O => \N__4631\,
            I => \N__4618\
        );

    \I__885\ : Sp12to4
    port map (
            O => \N__4628\,
            I => \N__4618\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4625\,
            I => \N__4618\
        );

    \I__883\ : Span12Mux_h
    port map (
            O => \N__4618\,
            I => \N__4615\
        );

    \I__882\ : Span12Mux_v
    port map (
            O => \N__4615\,
            I => \N__4612\
        );

    \I__881\ : Odrv12
    port map (
            O => \N__4612\,
            I => \TSn_c\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__4609\,
            I => \N__4606\
        );

    \I__879\ : InMux
    port map (
            O => \N__4606\,
            I => \N__4601\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__4605\,
            I => \N__4597\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__4604\,
            I => \N__4594\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4601\,
            I => \N__4591\
        );

    \I__875\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4588\
        );

    \I__874\ : InMux
    port map (
            O => \N__4597\,
            I => \N__4585\
        );

    \I__873\ : InMux
    port map (
            O => \N__4594\,
            I => \N__4582\
        );

    \I__872\ : Span4Mux_h
    port map (
            O => \N__4591\,
            I => \N__4575\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4588\,
            I => \N__4575\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4585\,
            I => \N__4575\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4582\,
            I => \N__4572\
        );

    \I__868\ : Span4Mux_v
    port map (
            O => \N__4575\,
            I => \N__4569\
        );

    \I__867\ : Span12Mux_v
    port map (
            O => \N__4572\,
            I => \N__4566\
        );

    \I__866\ : Span4Mux_h
    port map (
            O => \N__4569\,
            I => \N__4563\
        );

    \I__865\ : Odrv12
    port map (
            O => \N__4566\,
            I => \N_76\
        );

    \I__864\ : Odrv4
    port map (
            O => \N__4563\,
            I => \N_76\
        );

    \I__863\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4555\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4555\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\
        );

    \I__861\ : CascadeMux
    port map (
            O => \N__4552\,
            I => \N__4549\
        );

    \I__860\ : InMux
    port map (
            O => \N__4549\,
            I => \N__4546\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4546\,
            I => \U409_TRANSFER_ACK.ROM_TACK_EN_e_1\
        );

    \I__858\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4539\
        );

    \I__857\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4536\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4539\,
            I => \U409_TRANSFER_ACK.N_28_4\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4536\,
            I => \U409_TRANSFER_ACK.N_28_4\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__4531\,
            I => \N__4527\
        );

    \I__853\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4524\
        );

    \I__852\ : InMux
    port map (
            O => \N__4527\,
            I => \N__4521\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4524\,
            I => \N__4516\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4521\,
            I => \N__4516\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__4516\,
            I => \N__4513\
        );

    \I__848\ : Odrv4
    port map (
            O => \N__4513\,
            I => \U409_TRANSFER_ACK.N_28_3\
        );

    \I__847\ : InMux
    port map (
            O => \N__4510\,
            I => \N__4505\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__4509\,
            I => \N__4499\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__4508\,
            I => \N__4495\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4505\,
            I => \N__4492\
        );

    \I__843\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4483\
        );

    \I__842\ : InMux
    port map (
            O => \N__4503\,
            I => \N__4483\
        );

    \I__841\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4483\
        );

    \I__840\ : InMux
    port map (
            O => \N__4499\,
            I => \N__4483\
        );

    \I__839\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4478\
        );

    \I__838\ : InMux
    port map (
            O => \N__4495\,
            I => \N__4478\
        );

    \I__837\ : Odrv4
    port map (
            O => \N__4492\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4483\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4478\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__834\ : InMux
    port map (
            O => \N__4471\,
            I => \N__4468\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4468\,
            I => \un1_RAMSPACEn_i_i_a3\
        );

    \I__832\ : InMux
    port map (
            O => \N__4465\,
            I => \N__4462\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4462\,
            I => \N__4459\
        );

    \I__830\ : Span12Mux_h
    port map (
            O => \N__4459\,
            I => \N__4456\
        );

    \I__829\ : Span12Mux_h
    port map (
            O => \N__4456\,
            I => \N__4453\
        );

    \I__828\ : Span12Mux_v
    port map (
            O => \N__4453\,
            I => \N__4450\
        );

    \I__827\ : Odrv12
    port map (
            O => \N__4450\,
            I => \TACKn_in\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__4447\,
            I => \un1_REGSPACEn_i_i_a3_0_a2_cascade_\
        );

    \I__825\ : SRMux
    port map (
            O => \N__4444\,
            I => \N__4440\
        );

    \I__824\ : SRMux
    port map (
            O => \N__4443\,
            I => \N__4435\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__4440\,
            I => \N__4432\
        );

    \I__822\ : SRMux
    port map (
            O => \N__4439\,
            I => \N__4429\
        );

    \I__821\ : SRMux
    port map (
            O => \N__4438\,
            I => \N__4426\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4435\,
            I => \N__4422\
        );

    \I__819\ : Span4Mux_v
    port map (
            O => \N__4432\,
            I => \N__4419\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4429\,
            I => \N__4416\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4426\,
            I => \N__4413\
        );

    \I__816\ : SRMux
    port map (
            O => \N__4425\,
            I => \N__4410\
        );

    \I__815\ : Span4Mux_v
    port map (
            O => \N__4422\,
            I => \N__4399\
        );

    \I__814\ : Span4Mux_v
    port map (
            O => \N__4419\,
            I => \N__4399\
        );

    \I__813\ : Span4Mux_h
    port map (
            O => \N__4416\,
            I => \N__4399\
        );

    \I__812\ : Span4Mux_v
    port map (
            O => \N__4413\,
            I => \N__4399\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4410\,
            I => \N__4399\
        );

    \I__810\ : Span4Mux_h
    port map (
            O => \N__4399\,
            I => \N__4396\
        );

    \I__809\ : Odrv4
    port map (
            O => \N__4396\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__808\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4389\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__4392\,
            I => \N__4384\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4389\,
            I => \N__4381\
        );

    \I__805\ : InMux
    port map (
            O => \N__4388\,
            I => \N__4376\
        );

    \I__804\ : InMux
    port map (
            O => \N__4387\,
            I => \N__4376\
        );

    \I__803\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4373\
        );

    \I__802\ : Span4Mux_v
    port map (
            O => \N__4381\,
            I => \N__4367\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4376\,
            I => \N__4367\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4373\,
            I => \N__4364\
        );

    \I__799\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4361\
        );

    \I__798\ : Odrv4
    port map (
            O => \N__4367\,
            I => \N_90\
        );

    \I__797\ : Odrv4
    port map (
            O => \N__4364\,
            I => \N_90\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4361\,
            I => \N_90\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__4354\,
            I => \N__4348\
        );

    \I__794\ : InMux
    port map (
            O => \N__4353\,
            I => \N__4343\
        );

    \I__793\ : InMux
    port map (
            O => \N__4352\,
            I => \N__4343\
        );

    \I__792\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4338\
        );

    \I__791\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4338\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4343\,
            I => \N__4333\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__4338\,
            I => \N__4330\
        );

    \I__788\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4323\
        );

    \I__787\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4323\
        );

    \I__786\ : Span4Mux_v
    port map (
            O => \N__4333\,
            I => \N__4318\
        );

    \I__785\ : Span4Mux_v
    port map (
            O => \N__4330\,
            I => \N__4318\
        );

    \I__784\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4315\
        );

    \I__783\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4312\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__4323\,
            I => \N__4309\
        );

    \I__781\ : Span4Mux_h
    port map (
            O => \N__4318\,
            I => \N__4305\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4315\,
            I => \N__4300\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4312\,
            I => \N__4300\
        );

    \I__778\ : Span4Mux_v
    port map (
            O => \N__4309\,
            I => \N__4297\
        );

    \I__777\ : InMux
    port map (
            O => \N__4308\,
            I => \N__4294\
        );

    \I__776\ : Sp12to4
    port map (
            O => \N__4305\,
            I => \N__4285\
        );

    \I__775\ : Span12Mux_h
    port map (
            O => \N__4300\,
            I => \N__4285\
        );

    \I__774\ : Sp12to4
    port map (
            O => \N__4297\,
            I => \N__4285\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4294\,
            I => \N__4285\
        );

    \I__772\ : Odrv12
    port map (
            O => \N__4285\,
            I => \A_c_21\
        );

    \I__771\ : InMux
    port map (
            O => \N__4282\,
            I => \N__4277\
        );

    \I__770\ : InMux
    port map (
            O => \N__4281\,
            I => \N__4272\
        );

    \I__769\ : InMux
    port map (
            O => \N__4280\,
            I => \N__4272\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__4277\,
            I => \N__4269\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4272\,
            I => \N__4266\
        );

    \I__766\ : Span4Mux_h
    port map (
            O => \N__4269\,
            I => \N__4262\
        );

    \I__765\ : Span4Mux_h
    port map (
            O => \N__4266\,
            I => \N__4259\
        );

    \I__764\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4256\
        );

    \I__763\ : Odrv4
    port map (
            O => \N__4262\,
            I => \N_80\
        );

    \I__762\ : Odrv4
    port map (
            O => \N__4259\,
            I => \N_80\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4256\,
            I => \N_80\
        );

    \I__760\ : IoInMux
    port map (
            O => \N__4249\,
            I => \N__4246\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4246\,
            I => \N__4243\
        );

    \I__758\ : IoSpan4Mux
    port map (
            O => \N__4243\,
            I => \N__4240\
        );

    \I__757\ : IoSpan4Mux
    port map (
            O => \N__4240\,
            I => \N__4237\
        );

    \I__756\ : Span4Mux_s0_v
    port map (
            O => \N__4237\,
            I => \N__4234\
        );

    \I__755\ : Sp12to4
    port map (
            O => \N__4234\,
            I => \N__4231\
        );

    \I__754\ : Span12Mux_v
    port map (
            O => \N__4231\,
            I => \N__4228\
        );

    \I__753\ : Odrv12
    port map (
            O => \N__4228\,
            I => \N_52_i\
        );

    \I__752\ : InMux
    port map (
            O => \N__4225\,
            I => \N__4221\
        );

    \I__751\ : InMux
    port map (
            O => \N__4224\,
            I => \N__4218\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__4221\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4218\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__748\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4206\
        );

    \I__747\ : InMux
    port map (
            O => \N__4212\,
            I => \N__4197\
        );

    \I__746\ : InMux
    port map (
            O => \N__4211\,
            I => \N__4197\
        );

    \I__745\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4197\
        );

    \I__744\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4197\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__4206\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4197\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__741\ : InMux
    port map (
            O => \N__4192\,
            I => \N__4185\
        );

    \I__740\ : InMux
    port map (
            O => \N__4191\,
            I => \N__4176\
        );

    \I__739\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4176\
        );

    \I__738\ : InMux
    port map (
            O => \N__4189\,
            I => \N__4176\
        );

    \I__737\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4176\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4185\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__4176\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__734\ : InMux
    port map (
            O => \N__4171\,
            I => \N__4166\
        );

    \I__733\ : InMux
    port map (
            O => \N__4170\,
            I => \N__4161\
        );

    \I__732\ : InMux
    port map (
            O => \N__4169\,
            I => \N__4161\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4166\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4161\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__729\ : CEMux
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4153\,
            I => \U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en\
        );

    \I__727\ : IoInMux
    port map (
            O => \N__4150\,
            I => \N__4147\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4147\,
            I => \N__4144\
        );

    \I__725\ : IoSpan4Mux
    port map (
            O => \N__4144\,
            I => \N__4141\
        );

    \I__724\ : Span4Mux_s2_v
    port map (
            O => \N__4141\,
            I => \N__4138\
        );

    \I__723\ : Span4Mux_v
    port map (
            O => \N__4138\,
            I => \N__4135\
        );

    \I__722\ : Sp12to4
    port map (
            O => \N__4135\,
            I => \N__4131\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__4134\,
            I => \N__4128\
        );

    \I__720\ : Span12Mux_v
    port map (
            O => \N__4131\,
            I => \N__4125\
        );

    \I__719\ : InMux
    port map (
            O => \N__4128\,
            I => \N__4122\
        );

    \I__718\ : Odrv12
    port map (
            O => \N__4125\,
            I => \ROMENn_c\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4122\,
            I => \ROMENn_c\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__4117\,
            I => \N__4113\
        );

    \I__715\ : InMux
    port map (
            O => \N__4116\,
            I => \N__4110\
        );

    \I__714\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4107\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__4110\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4107\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__711\ : InMux
    port map (
            O => \N__4102\,
            I => \N__4099\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4099\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_0\
        );

    \I__709\ : InMux
    port map (
            O => \N__4096\,
            I => \N__4091\
        );

    \I__708\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4088\
        );

    \I__707\ : InMux
    port map (
            O => \N__4094\,
            I => \N__4085\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4091\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4088\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__4085\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__703\ : InMux
    port map (
            O => \N__4078\,
            I => \N__4072\
        );

    \I__702\ : InMux
    port map (
            O => \N__4077\,
            I => \N__4068\
        );

    \I__701\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4065\
        );

    \I__700\ : InMux
    port map (
            O => \N__4075\,
            I => \N__4062\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__4072\,
            I => \N__4059\
        );

    \I__698\ : InMux
    port map (
            O => \N__4071\,
            I => \N__4056\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4068\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__4065\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4062\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__694\ : Odrv4
    port map (
            O => \N__4059\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4056\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__4045\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__4042\,
            I => \N__4039\
        );

    \I__690\ : InMux
    port map (
            O => \N__4039\,
            I => \N__4031\
        );

    \I__689\ : InMux
    port map (
            O => \N__4038\,
            I => \N__4028\
        );

    \I__688\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4025\
        );

    \I__687\ : InMux
    port map (
            O => \N__4036\,
            I => \N__4022\
        );

    \I__686\ : InMux
    port map (
            O => \N__4035\,
            I => \N__4017\
        );

    \I__685\ : InMux
    port map (
            O => \N__4034\,
            I => \N__4017\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__4031\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4028\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__4025\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4022\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4017\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__4006\,
            I => \U409_TRANSFER_ACK.N_54_4_cascade_\
        );

    \I__678\ : InMux
    port map (
            O => \N__4003\,
            I => \N__4000\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4000\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_5\
        );

    \I__676\ : CascadeMux
    port map (
            O => \N__3997\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_5_cascade_\
        );

    \I__675\ : InMux
    port map (
            O => \N__3994\,
            I => \N__3991\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3991\,
            I => \N__3988\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__3988\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out\
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__3985\,
            I => \N__3982\
        );

    \I__671\ : InMux
    port map (
            O => \N__3982\,
            I => \N__3979\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3979\,
            I => \N__3974\
        );

    \I__669\ : InMux
    port map (
            O => \N__3978\,
            I => \N__3971\
        );

    \I__668\ : InMux
    port map (
            O => \N__3977\,
            I => \N__3968\
        );

    \I__667\ : Odrv4
    port map (
            O => \N__3974\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__3971\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3968\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__3961\,
            I => \N__3955\
        );

    \I__663\ : InMux
    port map (
            O => \N__3960\,
            I => \N__3951\
        );

    \I__662\ : InMux
    port map (
            O => \N__3959\,
            I => \N__3948\
        );

    \I__661\ : InMux
    port map (
            O => \N__3958\,
            I => \N__3945\
        );

    \I__660\ : InMux
    port map (
            O => \N__3955\,
            I => \N__3940\
        );

    \I__659\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3940\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3951\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3948\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3945\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__3940\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__3931\,
            I => \N__3928\
        );

    \I__653\ : InMux
    port map (
            O => \N__3928\,
            I => \N__3921\
        );

    \I__652\ : InMux
    port map (
            O => \N__3927\,
            I => \N__3918\
        );

    \I__651\ : InMux
    port map (
            O => \N__3926\,
            I => \N__3915\
        );

    \I__650\ : InMux
    port map (
            O => \N__3925\,
            I => \N__3910\
        );

    \I__649\ : InMux
    port map (
            O => \N__3924\,
            I => \N__3910\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__3921\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3918\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3915\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3910\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__644\ : InMux
    port map (
            O => \N__3901\,
            I => \N__3896\
        );

    \I__643\ : InMux
    port map (
            O => \N__3900\,
            I => \N__3888\
        );

    \I__642\ : InMux
    port map (
            O => \N__3899\,
            I => \N__3885\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3896\,
            I => \N__3882\
        );

    \I__640\ : InMux
    port map (
            O => \N__3895\,
            I => \N__3879\
        );

    \I__639\ : InMux
    port map (
            O => \N__3894\,
            I => \N__3876\
        );

    \I__638\ : InMux
    port map (
            O => \N__3893\,
            I => \N__3869\
        );

    \I__637\ : InMux
    port map (
            O => \N__3892\,
            I => \N__3869\
        );

    \I__636\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3869\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3888\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3885\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__633\ : Odrv4
    port map (
            O => \N__3882\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3879\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3876\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3869\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__3856\,
            I => \N__3853\
        );

    \I__628\ : InMux
    port map (
            O => \N__3853\,
            I => \N__3847\
        );

    \I__627\ : CascadeMux
    port map (
            O => \N__3852\,
            I => \N__3843\
        );

    \I__626\ : InMux
    port map (
            O => \N__3851\,
            I => \N__3838\
        );

    \I__625\ : InMux
    port map (
            O => \N__3850\,
            I => \N__3838\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3847\,
            I => \N__3835\
        );

    \I__623\ : InMux
    port map (
            O => \N__3846\,
            I => \N__3830\
        );

    \I__622\ : InMux
    port map (
            O => \N__3843\,
            I => \N__3830\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3838\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__620\ : Odrv4
    port map (
            O => \N__3835\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3830\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__618\ : InMux
    port map (
            O => \N__3823\,
            I => \N__3820\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3820\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a3_0_1_0\
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__3817\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a3_0_1_0_cascade_\
        );

    \I__615\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3810\
        );

    \I__614\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3807\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3810\,
            I => \U409_TRANSFER_ACK.N_54_4\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3807\,
            I => \U409_TRANSFER_ACK.N_54_4\
        );

    \I__611\ : InMux
    port map (
            O => \N__3802\,
            I => \N__3799\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3799\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0Z0Z_0\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__3796\,
            I => \N__3792\
        );

    \I__608\ : InMux
    port map (
            O => \N__3795\,
            I => \N__3787\
        );

    \I__607\ : InMux
    port map (
            O => \N__3792\,
            I => \N__3781\
        );

    \I__606\ : InMux
    port map (
            O => \N__3791\,
            I => \N__3781\
        );

    \I__605\ : InMux
    port map (
            O => \N__3790\,
            I => \N__3778\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3787\,
            I => \N__3775\
        );

    \I__603\ : InMux
    port map (
            O => \N__3786\,
            I => \N__3772\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3781\,
            I => \N__3769\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3778\,
            I => \N__3766\
        );

    \I__600\ : Span4Mux_v
    port map (
            O => \N__3775\,
            I => \N__3763\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3772\,
            I => \N__3760\
        );

    \I__598\ : Span4Mux_v
    port map (
            O => \N__3769\,
            I => \N__3757\
        );

    \I__597\ : Span4Mux_v
    port map (
            O => \N__3766\,
            I => \N__3754\
        );

    \I__596\ : Sp12to4
    port map (
            O => \N__3763\,
            I => \N__3749\
        );

    \I__595\ : Span12Mux_v
    port map (
            O => \N__3760\,
            I => \N__3749\
        );

    \I__594\ : Span4Mux_h
    port map (
            O => \N__3757\,
            I => \N__3746\
        );

    \I__593\ : Span4Mux_h
    port map (
            O => \N__3754\,
            I => \N__3743\
        );

    \I__592\ : Odrv12
    port map (
            O => \N__3749\,
            I => \A_c_23\
        );

    \I__591\ : Odrv4
    port map (
            O => \N__3746\,
            I => \A_c_23\
        );

    \I__590\ : Odrv4
    port map (
            O => \N__3743\,
            I => \A_c_23\
        );

    \I__589\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3733\,
            I => \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3Z0Z_4\
        );

    \I__587\ : InMux
    port map (
            O => \N__3730\,
            I => \N__3727\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3727\,
            I => \N__3723\
        );

    \I__585\ : InMux
    port map (
            O => \N__3726\,
            I => \N__3720\
        );

    \I__584\ : Odrv4
    port map (
            O => \N__3723\,
            I => \U409_ADDRESS_DECODE.N_16_i\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3720\,
            I => \U409_ADDRESS_DECODE.N_16_i\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__3715\,
            I => \un1_RAMSPACEn_i_i_a3_cascade_\
        );

    \I__581\ : IoInMux
    port map (
            O => \N__3712\,
            I => \N__3709\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3709\,
            I => \N__3706\
        );

    \I__579\ : Span4Mux_s1_v
    port map (
            O => \N__3706\,
            I => \N__3703\
        );

    \I__578\ : Sp12to4
    port map (
            O => \N__3703\,
            I => \N__3700\
        );

    \I__577\ : Span12Mux_h
    port map (
            O => \N__3700\,
            I => \N__3697\
        );

    \I__576\ : Span12Mux_v
    port map (
            O => \N__3697\,
            I => \N__3694\
        );

    \I__575\ : Odrv12
    port map (
            O => \N__3694\,
            I => \N_11_i\
        );

    \I__574\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3687\
        );

    \I__573\ : InMux
    port map (
            O => \N__3690\,
            I => \N__3684\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__3687\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3684\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__570\ : InMux
    port map (
            O => \N__3679\,
            I => \N__3675\
        );

    \I__569\ : InMux
    port map (
            O => \N__3678\,
            I => \N__3672\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3675\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__3672\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__566\ : CascadeMux
    port map (
            O => \N__3667\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__3664\,
            I => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\
        );

    \I__564\ : IoInMux
    port map (
            O => \N__3661\,
            I => \N__3658\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3658\,
            I => \N__3655\
        );

    \I__562\ : Span4Mux_s1_v
    port map (
            O => \N__3655\,
            I => \N__3652\
        );

    \I__561\ : Span4Mux_v
    port map (
            O => \N__3652\,
            I => \N__3649\
        );

    \I__560\ : Sp12to4
    port map (
            O => \N__3649\,
            I => \N__3646\
        );

    \I__559\ : Span12Mux_s10_h
    port map (
            O => \N__3646\,
            I => \N__3643\
        );

    \I__558\ : Span12Mux_v
    port map (
            O => \N__3643\,
            I => \N__3638\
        );

    \I__557\ : InMux
    port map (
            O => \N__3642\,
            I => \N__3633\
        );

    \I__556\ : InMux
    port map (
            O => \N__3641\,
            I => \N__3633\
        );

    \I__555\ : Odrv12
    port map (
            O => \N__3638\,
            I => \TACK_OUTn\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3633\,
            I => \TACK_OUTn\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__3628\,
            I => \N__3624\
        );

    \I__552\ : InMux
    port map (
            O => \N__3627\,
            I => \N__3621\
        );

    \I__551\ : InMux
    port map (
            O => \N__3624\,
            I => \N__3618\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3621\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_6\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3618\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_6\
        );

    \I__548\ : InMux
    port map (
            O => \N__3613\,
            I => \N__3610\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3610\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3\
        );

    \I__546\ : InMux
    port map (
            O => \N__3607\,
            I => \N__3600\
        );

    \I__545\ : InMux
    port map (
            O => \N__3606\,
            I => \N__3597\
        );

    \I__544\ : InMux
    port map (
            O => \N__3605\,
            I => \N__3594\
        );

    \I__543\ : InMux
    port map (
            O => \N__3604\,
            I => \N__3591\
        );

    \I__542\ : InMux
    port map (
            O => \N__3603\,
            I => \N__3588\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3600\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__3597\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3594\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3591\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3588\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__536\ : InMux
    port map (
            O => \N__3577\,
            I => \N__3572\
        );

    \I__535\ : InMux
    port map (
            O => \N__3576\,
            I => \N__3568\
        );

    \I__534\ : InMux
    port map (
            O => \N__3575\,
            I => \N__3565\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3572\,
            I => \N__3562\
        );

    \I__532\ : InMux
    port map (
            O => \N__3571\,
            I => \N__3559\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3568\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3565\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__529\ : Odrv4
    port map (
            O => \N__3562\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3559\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__527\ : CascadeMux
    port map (
            O => \N__3550\,
            I => \N__3547\
        );

    \I__526\ : InMux
    port map (
            O => \N__3547\,
            I => \N__3544\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3544\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__3541\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__523\ : InMux
    port map (
            O => \N__3538\,
            I => \N__3534\
        );

    \I__522\ : InMux
    port map (
            O => \N__3537\,
            I => \N__3531\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3534\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3531\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__519\ : CascadeMux
    port map (
            O => \N__3526\,
            I => \N__3522\
        );

    \I__518\ : InMux
    port map (
            O => \N__3525\,
            I => \N__3519\
        );

    \I__517\ : InMux
    port map (
            O => \N__3522\,
            I => \N__3516\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3519\,
            I => \N__3511\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3516\,
            I => \N__3511\
        );

    \I__514\ : Span4Mux_v
    port map (
            O => \N__3511\,
            I => \N__3508\
        );

    \I__513\ : Odrv4
    port map (
            O => \N__3508\,
            I => \U409_CIA.N_89\
        );

    \I__512\ : InMux
    port map (
            O => \N__3505\,
            I => \N__3497\
        );

    \I__511\ : InMux
    port map (
            O => \N__3504\,
            I => \N__3497\
        );

    \I__510\ : InMux
    port map (
            O => \N__3503\,
            I => \N__3494\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__3502\,
            I => \N__3490\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3497\,
            I => \N__3487\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3494\,
            I => \N__3484\
        );

    \I__506\ : InMux
    port map (
            O => \N__3493\,
            I => \N__3479\
        );

    \I__505\ : InMux
    port map (
            O => \N__3490\,
            I => \N__3479\
        );

    \I__504\ : Span4Mux_v
    port map (
            O => \N__3487\,
            I => \N__3476\
        );

    \I__503\ : Span4Mux_h
    port map (
            O => \N__3484\,
            I => \N__3471\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3479\,
            I => \N__3468\
        );

    \I__501\ : Span4Mux_v
    port map (
            O => \N__3476\,
            I => \N__3465\
        );

    \I__500\ : InMux
    port map (
            O => \N__3475\,
            I => \N__3460\
        );

    \I__499\ : InMux
    port map (
            O => \N__3474\,
            I => \N__3460\
        );

    \I__498\ : Span4Mux_h
    port map (
            O => \N__3471\,
            I => \N__3455\
        );

    \I__497\ : Span4Mux_v
    port map (
            O => \N__3468\,
            I => \N__3455\
        );

    \I__496\ : Span4Mux_v
    port map (
            O => \N__3465\,
            I => \N__3452\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3460\,
            I => \N__3449\
        );

    \I__494\ : Span4Mux_v
    port map (
            O => \N__3455\,
            I => \N__3446\
        );

    \I__493\ : Span4Mux_h
    port map (
            O => \N__3452\,
            I => \N__3443\
        );

    \I__492\ : Sp12to4
    port map (
            O => \N__3449\,
            I => \N__3440\
        );

    \I__491\ : Span4Mux_v
    port map (
            O => \N__3446\,
            I => \N__3437\
        );

    \I__490\ : Sp12to4
    port map (
            O => \N__3443\,
            I => \N__3432\
        );

    \I__489\ : Span12Mux_v
    port map (
            O => \N__3440\,
            I => \N__3432\
        );

    \I__488\ : Span4Mux_h
    port map (
            O => \N__3437\,
            I => \N__3429\
        );

    \I__487\ : Odrv12
    port map (
            O => \N__3432\,
            I => \A_c_22\
        );

    \I__486\ : Odrv4
    port map (
            O => \N__3429\,
            I => \A_c_22\
        );

    \I__485\ : InMux
    port map (
            O => \N__3424\,
            I => \N__3421\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3421\,
            I => \N__3418\
        );

    \I__483\ : Span4Mux_v
    port map (
            O => \N__3418\,
            I => \N__3414\
        );

    \I__482\ : InMux
    port map (
            O => \N__3417\,
            I => \N__3411\
        );

    \I__481\ : Span4Mux_h
    port map (
            O => \N__3414\,
            I => \N__3408\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3411\,
            I => \N__3405\
        );

    \I__479\ : Sp12to4
    port map (
            O => \N__3408\,
            I => \N__3400\
        );

    \I__478\ : Span12Mux_v
    port map (
            O => \N__3405\,
            I => \N__3400\
        );

    \I__477\ : Span12Mux_v
    port map (
            O => \N__3400\,
            I => \N__3397\
        );

    \I__476\ : Span12Mux_h
    port map (
            O => \N__3397\,
            I => \N__3394\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__3394\,
            I => \OVL_c\
        );

    \I__474\ : CascadeMux
    port map (
            O => \N__3391\,
            I => \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3Z0Z_4_cascade_\
        );

    \I__473\ : IoInMux
    port map (
            O => \N__3388\,
            I => \N__3385\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3385\,
            I => \N__3382\
        );

    \I__471\ : Span4Mux_s2_v
    port map (
            O => \N__3382\,
            I => \N__3379\
        );

    \I__470\ : Span4Mux_h
    port map (
            O => \N__3379\,
            I => \N__3376\
        );

    \I__469\ : Sp12to4
    port map (
            O => \N__3376\,
            I => \N__3373\
        );

    \I__468\ : Span12Mux_v
    port map (
            O => \N__3373\,
            I => \N__3370\
        );

    \I__467\ : Odrv12
    port map (
            O => \N__3370\,
            I => \N_53_i\
        );

    \I__466\ : InMux
    port map (
            O => \N__3367\,
            I => \N__3364\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3364\,
            I => \N__3361\
        );

    \I__464\ : Odrv4
    port map (
            O => \N__3361\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_17\
        );

    \I__463\ : InMux
    port map (
            O => \N__3358\,
            I => \N__3355\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3355\,
            I => \N__3352\
        );

    \I__461\ : Span4Mux_v
    port map (
            O => \N__3352\,
            I => \N__3349\
        );

    \I__460\ : Odrv4
    port map (
            O => \N__3349\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_16\
        );

    \I__459\ : InMux
    port map (
            O => \N__3346\,
            I => \N__3339\
        );

    \I__458\ : InMux
    port map (
            O => \N__3345\,
            I => \N__3339\
        );

    \I__457\ : InMux
    port map (
            O => \N__3344\,
            I => \N__3336\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__3339\,
            I => \N__3331\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__3336\,
            I => \N__3331\
        );

    \I__454\ : Span12Mux_h
    port map (
            O => \N__3331\,
            I => \N__3328\
        );

    \I__453\ : Span12Mux_v
    port map (
            O => \N__3328\,
            I => \N__3325\
        );

    \I__452\ : Odrv12
    port map (
            O => \N__3325\,
            I => \TM_c_0\
        );

    \I__451\ : InMux
    port map (
            O => \N__3322\,
            I => \N__3316\
        );

    \I__450\ : InMux
    port map (
            O => \N__3321\,
            I => \N__3316\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3316\,
            I => \N__3312\
        );

    \I__448\ : InMux
    port map (
            O => \N__3315\,
            I => \N__3309\
        );

    \I__447\ : Span4Mux_h
    port map (
            O => \N__3312\,
            I => \N__3304\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__3309\,
            I => \N__3304\
        );

    \I__445\ : Span4Mux_h
    port map (
            O => \N__3304\,
            I => \N__3301\
        );

    \I__444\ : Sp12to4
    port map (
            O => \N__3301\,
            I => \N__3298\
        );

    \I__443\ : Odrv12
    port map (
            O => \N__3298\,
            I => \TM_c_1\
        );

    \I__442\ : IoInMux
    port map (
            O => \N__3295\,
            I => \N__3292\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3292\,
            I => \N__3289\
        );

    \I__440\ : IoSpan4Mux
    port map (
            O => \N__3289\,
            I => \N__3286\
        );

    \I__439\ : Span4Mux_s0_v
    port map (
            O => \N__3286\,
            I => \N__3283\
        );

    \I__438\ : Sp12to4
    port map (
            O => \N__3283\,
            I => \N__3280\
        );

    \I__437\ : Span12Mux_v
    port map (
            O => \N__3280\,
            I => \N__3277\
        );

    \I__436\ : Odrv12
    port map (
            O => \N__3277\,
            I => \PORTSIZE_i_a2\
        );

    \I__435\ : InMux
    port map (
            O => \N__3274\,
            I => \N__3271\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3271\,
            I => \N__3268\
        );

    \I__433\ : Span4Mux_v
    port map (
            O => \N__3268\,
            I => \N__3265\
        );

    \I__432\ : Span4Mux_v
    port map (
            O => \N__3265\,
            I => \N__3262\
        );

    \I__431\ : Odrv4
    port map (
            O => \N__3262\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_12\
        );

    \I__430\ : InMux
    port map (
            O => \N__3259\,
            I => \N__3256\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3256\,
            I => \N__3253\
        );

    \I__428\ : Span4Mux_h
    port map (
            O => \N__3253\,
            I => \N__3249\
        );

    \I__427\ : InMux
    port map (
            O => \N__3252\,
            I => \N__3246\
        );

    \I__426\ : Odrv4
    port map (
            O => \N__3249\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3246\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__424\ : InMux
    port map (
            O => \N__3241\,
            I => \N__3235\
        );

    \I__423\ : InMux
    port map (
            O => \N__3240\,
            I => \N__3235\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3235\,
            I => \N__3231\
        );

    \I__421\ : InMux
    port map (
            O => \N__3234\,
            I => \N__3228\
        );

    \I__420\ : Span4Mux_v
    port map (
            O => \N__3231\,
            I => \N__3225\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3228\,
            I => \N__3222\
        );

    \I__418\ : Odrv4
    port map (
            O => \N__3225\,
            I => \U409_CIA_PORTSIZE_i_a2_0_3\
        );

    \I__417\ : Odrv12
    port map (
            O => \N__3222\,
            I => \U409_CIA_PORTSIZE_i_a2_0_3\
        );

    \I__416\ : CascadeMux
    port map (
            O => \N__3217\,
            I => \N__3214\
        );

    \I__415\ : InMux
    port map (
            O => \N__3214\,
            I => \N__3209\
        );

    \I__414\ : InMux
    port map (
            O => \N__3213\,
            I => \N__3206\
        );

    \I__413\ : InMux
    port map (
            O => \N__3212\,
            I => \N__3203\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__3209\,
            I => \N__3199\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3206\,
            I => \N__3194\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__3203\,
            I => \N__3194\
        );

    \I__409\ : InMux
    port map (
            O => \N__3202\,
            I => \N__3191\
        );

    \I__408\ : Span4Mux_v
    port map (
            O => \N__3199\,
            I => \N__3186\
        );

    \I__407\ : Span4Mux_v
    port map (
            O => \N__3194\,
            I => \N__3186\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3191\,
            I => \N__3183\
        );

    \I__405\ : Sp12to4
    port map (
            O => \N__3186\,
            I => \N__3180\
        );

    \I__404\ : Span4Mux_h
    port map (
            O => \N__3183\,
            I => \N__3177\
        );

    \I__403\ : Span12Mux_h
    port map (
            O => \N__3180\,
            I => \N__3172\
        );

    \I__402\ : Sp12to4
    port map (
            O => \N__3177\,
            I => \N__3172\
        );

    \I__401\ : Span12Mux_v
    port map (
            O => \N__3172\,
            I => \N__3169\
        );

    \I__400\ : Odrv12
    port map (
            O => \N__3169\,
            I => \A_c_19\
        );

    \I__399\ : CascadeMux
    port map (
            O => \N__3166\,
            I => \N__3162\
        );

    \I__398\ : InMux
    port map (
            O => \N__3165\,
            I => \N__3158\
        );

    \I__397\ : InMux
    port map (
            O => \N__3162\,
            I => \N__3155\
        );

    \I__396\ : InMux
    port map (
            O => \N__3161\,
            I => \N__3152\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__3158\,
            I => \N__3145\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3155\,
            I => \N__3145\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3152\,
            I => \N__3145\
        );

    \I__392\ : Span4Mux_v
    port map (
            O => \N__3145\,
            I => \N__3142\
        );

    \I__391\ : Sp12to4
    port map (
            O => \N__3142\,
            I => \N__3139\
        );

    \I__390\ : Span12Mux_h
    port map (
            O => \N__3139\,
            I => \N__3136\
        );

    \I__389\ : Span12Mux_v
    port map (
            O => \N__3136\,
            I => \N__3133\
        );

    \I__388\ : Odrv12
    port map (
            O => \N__3133\,
            I => \A_c_18\
        );

    \I__387\ : CascadeMux
    port map (
            O => \N__3130\,
            I => \N__3127\
        );

    \I__386\ : InMux
    port map (
            O => \N__3127\,
            I => \N__3124\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__3124\,
            I => \N__3120\
        );

    \I__384\ : InMux
    port map (
            O => \N__3123\,
            I => \N__3117\
        );

    \I__383\ : Span4Mux_h
    port map (
            O => \N__3120\,
            I => \N__3112\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3117\,
            I => \N__3112\
        );

    \I__381\ : Span4Mux_v
    port map (
            O => \N__3112\,
            I => \N__3109\
        );

    \I__380\ : Span4Mux_h
    port map (
            O => \N__3109\,
            I => \N__3106\
        );

    \I__379\ : Sp12to4
    port map (
            O => \N__3106\,
            I => \N__3103\
        );

    \I__378\ : Odrv12
    port map (
            O => \N__3103\,
            I => \TT_c_0\
        );

    \I__377\ : InMux
    port map (
            O => \N__3100\,
            I => \N__3094\
        );

    \I__376\ : InMux
    port map (
            O => \N__3099\,
            I => \N__3094\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__3094\,
            I => \N__3090\
        );

    \I__374\ : InMux
    port map (
            O => \N__3093\,
            I => \N__3087\
        );

    \I__373\ : Span4Mux_h
    port map (
            O => \N__3090\,
            I => \N__3082\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3087\,
            I => \N__3082\
        );

    \I__371\ : Span4Mux_v
    port map (
            O => \N__3082\,
            I => \N__3079\
        );

    \I__370\ : Span4Mux_v
    port map (
            O => \N__3079\,
            I => \N__3076\
        );

    \I__369\ : Span4Mux_h
    port map (
            O => \N__3076\,
            I => \N__3073\
        );

    \I__368\ : Odrv4
    port map (
            O => \N__3073\,
            I => \A_c_26\
        );

    \I__367\ : InMux
    port map (
            O => \N__3070\,
            I => \N__3064\
        );

    \I__366\ : InMux
    port map (
            O => \N__3069\,
            I => \N__3064\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__3064\,
            I => \N__3061\
        );

    \I__364\ : Span4Mux_v
    port map (
            O => \N__3061\,
            I => \N__3058\
        );

    \I__363\ : Span4Mux_h
    port map (
            O => \N__3058\,
            I => \N__3055\
        );

    \I__362\ : Sp12to4
    port map (
            O => \N__3055\,
            I => \N__3052\
        );

    \I__361\ : Odrv12
    port map (
            O => \N__3052\,
            I => \TT_c_1\
        );

    \I__360\ : CascadeMux
    port map (
            O => \N__3049\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_11_cascade_\
        );

    \I__359\ : InMux
    port map (
            O => \N__3046\,
            I => \N__3043\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3043\,
            I => \N__3040\
        );

    \I__357\ : Odrv4
    port map (
            O => \N__3040\,
            I => \U409_TRANSFER_ACK.N_17\
        );

    \I__356\ : InMux
    port map (
            O => \N__3037\,
            I => \N__3033\
        );

    \I__355\ : InMux
    port map (
            O => \N__3036\,
            I => \N__3030\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__3033\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_4\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__3030\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_4\
        );

    \I__352\ : CascadeMux
    port map (
            O => \N__3025\,
            I => \N__3021\
        );

    \I__351\ : InMux
    port map (
            O => \N__3024\,
            I => \N__3018\
        );

    \I__350\ : InMux
    port map (
            O => \N__3021\,
            I => \N__3015\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__3018\,
            I => \N__3010\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3015\,
            I => \N__3010\
        );

    \I__347\ : Odrv12
    port map (
            O => \N__3010\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_11\
        );

    \I__346\ : InMux
    port map (
            O => \N__3007\,
            I => \N__3004\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__3004\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_14\
        );

    \I__344\ : InMux
    port map (
            O => \N__3001\,
            I => \N__2998\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2998\,
            I => \N__2994\
        );

    \I__342\ : InMux
    port map (
            O => \N__2997\,
            I => \N__2991\
        );

    \I__341\ : Span4Mux_v
    port map (
            O => \N__2994\,
            I => \N__2988\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2991\,
            I => \N__2985\
        );

    \I__339\ : Span4Mux_h
    port map (
            O => \N__2988\,
            I => \N__2982\
        );

    \I__338\ : Span4Mux_v
    port map (
            O => \N__2985\,
            I => \N__2979\
        );

    \I__337\ : Odrv4
    port map (
            O => \N__2982\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_10\
        );

    \I__336\ : Odrv4
    port map (
            O => \N__2979\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_10\
        );

    \I__335\ : InMux
    port map (
            O => \N__2974\,
            I => \N__2971\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2971\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1\
        );

    \I__333\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2965\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2965\,
            I => \N__2961\
        );

    \I__331\ : InMux
    port map (
            O => \N__2964\,
            I => \N__2958\
        );

    \I__330\ : Span4Mux_v
    port map (
            O => \N__2961\,
            I => \N__2953\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2958\,
            I => \N__2953\
        );

    \I__328\ : Span4Mux_h
    port map (
            O => \N__2953\,
            I => \N__2950\
        );

    \I__327\ : Span4Mux_v
    port map (
            O => \N__2950\,
            I => \N__2947\
        );

    \I__326\ : Odrv4
    port map (
            O => \N__2947\,
            I => \A_c_31\
        );

    \I__325\ : CascadeMux
    port map (
            O => \N__2944\,
            I => \N__2940\
        );

    \I__324\ : CascadeMux
    port map (
            O => \N__2943\,
            I => \N__2937\
        );

    \I__323\ : InMux
    port map (
            O => \N__2940\,
            I => \N__2934\
        );

    \I__322\ : InMux
    port map (
            O => \N__2937\,
            I => \N__2931\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2934\,
            I => \N__2926\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2931\,
            I => \N__2926\
        );

    \I__319\ : Span4Mux_v
    port map (
            O => \N__2926\,
            I => \N__2923\
        );

    \I__318\ : Span4Mux_v
    port map (
            O => \N__2923\,
            I => \N__2920\
        );

    \I__317\ : Span4Mux_h
    port map (
            O => \N__2920\,
            I => \N__2917\
        );

    \I__316\ : Odrv4
    port map (
            O => \N__2917\,
            I => \A_c_24\
        );

    \I__315\ : InMux
    port map (
            O => \N__2914\,
            I => \N__2910\
        );

    \I__314\ : InMux
    port map (
            O => \N__2913\,
            I => \N__2907\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2910\,
            I => \N__2902\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2907\,
            I => \N__2902\
        );

    \I__311\ : Span4Mux_v
    port map (
            O => \N__2902\,
            I => \N__2899\
        );

    \I__310\ : Span4Mux_h
    port map (
            O => \N__2899\,
            I => \N__2896\
        );

    \I__309\ : Odrv4
    port map (
            O => \N__2896\,
            I => \A_c_25\
        );

    \I__308\ : InMux
    port map (
            O => \N__2893\,
            I => \N__2890\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2890\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_3\
        );

    \I__306\ : InMux
    port map (
            O => \N__2887\,
            I => \N__2884\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2884\,
            I => \N__2880\
        );

    \I__304\ : InMux
    port map (
            O => \N__2883\,
            I => \N__2877\
        );

    \I__303\ : Span4Mux_h
    port map (
            O => \N__2880\,
            I => \N__2872\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2877\,
            I => \N__2872\
        );

    \I__301\ : Span4Mux_v
    port map (
            O => \N__2872\,
            I => \N__2869\
        );

    \I__300\ : Span4Mux_h
    port map (
            O => \N__2869\,
            I => \N__2866\
        );

    \I__299\ : Odrv4
    port map (
            O => \N__2866\,
            I => \A_c_30\
        );

    \I__298\ : CascadeMux
    port map (
            O => \N__2863\,
            I => \N__2860\
        );

    \I__297\ : InMux
    port map (
            O => \N__2860\,
            I => \N__2854\
        );

    \I__296\ : InMux
    port map (
            O => \N__2859\,
            I => \N__2854\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2854\,
            I => \N__2851\
        );

    \I__294\ : Span4Mux_h
    port map (
            O => \N__2851\,
            I => \N__2848\
        );

    \I__293\ : Span4Mux_v
    port map (
            O => \N__2848\,
            I => \N__2845\
        );

    \I__292\ : Span4Mux_v
    port map (
            O => \N__2845\,
            I => \N__2842\
        );

    \I__291\ : Odrv4
    port map (
            O => \N__2842\,
            I => \A_c_28\
        );

    \I__290\ : InMux
    port map (
            O => \N__2839\,
            I => \N__2833\
        );

    \I__289\ : InMux
    port map (
            O => \N__2838\,
            I => \N__2833\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2833\,
            I => \N__2830\
        );

    \I__287\ : Sp12to4
    port map (
            O => \N__2830\,
            I => \N__2827\
        );

    \I__286\ : Span12Mux_v
    port map (
            O => \N__2827\,
            I => \N__2824\
        );

    \I__285\ : Odrv12
    port map (
            O => \N__2824\,
            I => \A_c_29\
        );

    \I__284\ : CascadeMux
    port map (
            O => \N__2821\,
            I => \N__2817\
        );

    \I__283\ : InMux
    port map (
            O => \N__2820\,
            I => \N__2814\
        );

    \I__282\ : InMux
    port map (
            O => \N__2817\,
            I => \N__2811\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2814\,
            I => \N__2806\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2811\,
            I => \N__2806\
        );

    \I__279\ : Odrv12
    port map (
            O => \N__2806\,
            I => \A_c_27\
        );

    \I__278\ : InMux
    port map (
            O => \N__2803\,
            I => \N__2800\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2800\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4\
        );

    \I__276\ : InMux
    port map (
            O => \N__2797\,
            I => \N__2794\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2794\,
            I => \N__2790\
        );

    \I__274\ : CascadeMux
    port map (
            O => \N__2793\,
            I => \N__2787\
        );

    \I__273\ : Span4Mux_v
    port map (
            O => \N__2790\,
            I => \N__2784\
        );

    \I__272\ : InMux
    port map (
            O => \N__2787\,
            I => \N__2781\
        );

    \I__271\ : Sp12to4
    port map (
            O => \N__2784\,
            I => \N__2776\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2781\,
            I => \N__2776\
        );

    \I__269\ : Odrv12
    port map (
            O => \N__2776\,
            I => \A_c_20\
        );

    \I__268\ : CascadeMux
    port map (
            O => \N__2773\,
            I => \U409_TRANSFER_ACK.N_41_cascade_\
        );

    \I__267\ : InMux
    port map (
            O => \N__2770\,
            I => \N__2767\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2767\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3Z0Z_2\
        );

    \I__265\ : InMux
    port map (
            O => \N__2764\,
            I => \N__2761\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2761\,
            I => \N__2758\
        );

    \I__263\ : Span4Mux_v
    port map (
            O => \N__2758\,
            I => \N__2755\
        );

    \I__262\ : Sp12to4
    port map (
            O => \N__2755\,
            I => \N__2752\
        );

    \I__261\ : Span12Mux_s3_h
    port map (
            O => \N__2752\,
            I => \N__2749\
        );

    \I__260\ : Span12Mux_v
    port map (
            O => \N__2749\,
            I => \N__2746\
        );

    \I__259\ : Odrv12
    port map (
            O => \N__2746\,
            I => \A_c_16\
        );

    \I__258\ : InMux
    port map (
            O => \N__2743\,
            I => \N__2740\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2740\,
            I => \N__2737\
        );

    \I__256\ : Span4Mux_v
    port map (
            O => \N__2737\,
            I => \N__2734\
        );

    \I__255\ : Sp12to4
    port map (
            O => \N__2734\,
            I => \N__2731\
        );

    \I__254\ : Span12Mux_v
    port map (
            O => \N__2731\,
            I => \N__2728\
        );

    \I__253\ : Odrv12
    port map (
            O => \N__2728\,
            I => \A_c_17\
        );

    \I__252\ : ClkMux
    port map (
            O => \N__2725\,
            I => \N__2677\
        );

    \I__251\ : ClkMux
    port map (
            O => \N__2724\,
            I => \N__2677\
        );

    \I__250\ : ClkMux
    port map (
            O => \N__2723\,
            I => \N__2677\
        );

    \I__249\ : ClkMux
    port map (
            O => \N__2722\,
            I => \N__2677\
        );

    \I__248\ : ClkMux
    port map (
            O => \N__2721\,
            I => \N__2677\
        );

    \I__247\ : ClkMux
    port map (
            O => \N__2720\,
            I => \N__2677\
        );

    \I__246\ : ClkMux
    port map (
            O => \N__2719\,
            I => \N__2677\
        );

    \I__245\ : ClkMux
    port map (
            O => \N__2718\,
            I => \N__2677\
        );

    \I__244\ : ClkMux
    port map (
            O => \N__2717\,
            I => \N__2677\
        );

    \I__243\ : ClkMux
    port map (
            O => \N__2716\,
            I => \N__2677\
        );

    \I__242\ : ClkMux
    port map (
            O => \N__2715\,
            I => \N__2677\
        );

    \I__241\ : ClkMux
    port map (
            O => \N__2714\,
            I => \N__2677\
        );

    \I__240\ : ClkMux
    port map (
            O => \N__2713\,
            I => \N__2677\
        );

    \I__239\ : ClkMux
    port map (
            O => \N__2712\,
            I => \N__2677\
        );

    \I__238\ : ClkMux
    port map (
            O => \N__2711\,
            I => \N__2677\
        );

    \I__237\ : ClkMux
    port map (
            O => \N__2710\,
            I => \N__2677\
        );

    \I__236\ : GlobalMux
    port map (
            O => \N__2677\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            I => \N__2712\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            I => \N__2711\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            I => \N__2710\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__2713\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            I => \N__2721\
        );

    \INVU409_TRANSFER_ACK.ROMENnC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            I => \N__2717\
        );

    \INVU409_TRANSFER_ACK.TACK_EN_iC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            I => \N__2715\
        );

    \INVU409_TRANSFER_ACK.CIA_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            I => \N__2714\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            I => \N__2723\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            I => \N__2720\
        );

    \INVU409_TRANSFER_ACK.TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            I => \N__2716\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            I => \N__2724\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            I => \N__2722\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            I => \N__2719\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\,
            I => \N__2718\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            I => \N__2725\
        );

    \IN_MUX_bfv_13_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_2_0_\
        );

    \IN_MUX_bfv_13_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_13_3_0_\
        );

    \IN_MUX_bfv_15_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_1_0_\
        );

    \IN_MUX_bfv_15_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_15_2_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_12_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_CIA.PORTSIZE_i_a2_0_3_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2764\,
            in1 => \N__3790\,
            in2 => \N__2793\,
            in3 => \N__2743\,
            lcout => \U409_CIA_PORTSIZE_i_a2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_11_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2968\,
            in1 => \N__2914\,
            in2 => \N__2944\,
            in3 => \N__4308\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__2893\,
            in1 => \N__2964\,
            in2 => \N__2943\,
            in3 => \N__2803\,
            lcout => \N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_3_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2887\,
            in2 => \_gnd_net_\,
            in3 => \N__2913\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_10_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2883\,
            in1 => \N__2839\,
            in2 => \N__2863\,
            in3 => \N__2820\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2859\,
            in1 => \N__2838\,
            in2 => \N__2821\,
            in3 => \N__3093\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_0_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__3424\,
            in1 => \N__3791\,
            in2 => \N__3502\,
            in3 => \N__4336\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.N_41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__2797\,
            in1 => \N__2770\,
            in2 => \N__2773\,
            in3 => \N__3493\,
            lcout => \U409_TRANSFER_ACK.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_2_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__4337\,
            in1 => \_gnd_net_\,
            in2 => \N__3796\,
            in3 => \N__3202\,
            lcout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.PORTSIZE_i_a2_0_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3234\,
            in1 => \N__3212\,
            in2 => \_gnd_net_\,
            in3 => \N__3161\,
            lcout => \U409_CIA.N_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_0_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3241\,
            in1 => \N__3475\,
            in2 => \N__3130\,
            in3 => \N__3036\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a2_0_0_a2_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3474\,
            in1 => \N__3213\,
            in2 => \N__3166\,
            in3 => \N__3240\,
            lcout => \N_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_2_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3069\,
            in1 => \N__3099\,
            in2 => \N__3217\,
            in3 => \N__3165\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_1_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4265\,
            in1 => \N__3123\,
            in2 => \N__3025\,
            in3 => \N__3037\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3100\,
            in1 => \N__3070\,
            in2 => \N__3049\,
            in3 => \N__2997\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_3_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__3315\,
            in1 => \N__3046\,
            in2 => \_gnd_net_\,
            in3 => \N__3344\,
            lcout => \U409_TRANSFER_ACK.N_28_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_4_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5371\,
            in2 => \_gnd_net_\,
            in3 => \N__4634\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_1_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3024\,
            in1 => \N__3007\,
            in2 => \_gnd_net_\,
            in3 => \N__3001\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2974\,
            in1 => \N__3901\,
            in2 => \_gnd_net_\,
            in3 => \N__3605\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4078\,
            in1 => \N__4036\,
            in2 => \N__3856\,
            in3 => \N__3577\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3367\,
            in1 => \N__3358\,
            in2 => \N__4805\,
            in3 => \N__3252\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un2_ROMEN_0_i_0_x3_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__3346\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3322\,
            lcout => \U409_ADDRESS_DECODE.N_16_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a3_0_a2_0_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__3345\,
            in1 => \N__3321\,
            in2 => \N__4605\,
            in3 => \N__5367\,
            lcout => \N_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.PORTSIZE_i_a2_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010000000"
        )
    port map (
            in0 => \N__4372\,
            in1 => \N__3503\,
            in2 => \N__3526\,
            in3 => \N__4328\,
            lcout => \PORTSIZE_i_a2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__3274\,
            in1 => \N__3259\,
            in2 => \N__4806\,
            in3 => \N__3691\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5243\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__3900\,
            in1 => \N__3576\,
            in2 => \_gnd_net_\,
            in3 => \N__3607\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__4443\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__3627\,
            in1 => \N__3679\,
            in2 => \_gnd_net_\,
            in3 => \N__4003\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__4443\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__4077\,
            in1 => \N__3978\,
            in2 => \N__4042\,
            in3 => \N__3959\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__4443\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3927\,
            in2 => \N__3961\,
            in3 => \N__3537\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__4444\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__4774\,
            in1 => \N__3823\,
            in2 => \N__3628\,
            in3 => \N__3814\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3899\,
            in2 => \N__3541\,
            in3 => \N__3606\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__4444\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3977\,
            in1 => \N__4038\,
            in2 => \_gnd_net_\,
            in3 => \N__3954\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__4444\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__3538\,
            in1 => \N__4096\,
            in2 => \N__3931\,
            in3 => \N__3960\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__4439\
        );

    \U409_CIA.VMA_RNO_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__3525\,
            in1 => \N__3505\,
            in2 => \N__4392\,
            in3 => \N__4351\,
            lcout => \U409_CIA.VMA_3_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3_4_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__3504\,
            in1 => \N__5366\,
            in2 => \N__4354\,
            in3 => \N__3417\,
            lcout => \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3Z0Z_4\,
            ltout => \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.N_53_i_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__3786\,
            in1 => \N__3726\,
            in2 => \N__3391\,
            in3 => \N__4600\,
            lcout => \N_53_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__4211\,
            in1 => \N__5349\,
            in2 => \_gnd_net_\,
            in3 => \N__4190\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110011111"
        )
    port map (
            in0 => \N__4210\,
            in1 => \N__4189\,
            in2 => \N__5364\,
            in3 => \N__4169\,
            lcout => \U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000110000"
        )
    port map (
            in0 => \N__4212\,
            in1 => \N__4191\,
            in2 => \N__5363\,
            in3 => \N__4170\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNINULI_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3690\,
            in1 => \N__4224\,
            in2 => \N__4117\,
            in3 => \N__3678\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER6\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111011101"
        )
    port map (
            in0 => \N__4209\,
            in1 => \N__4188\,
            in2 => \N__3667\,
            in3 => \N__3641\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__3642\,
            in1 => \_gnd_net_\,
            in2 => \N__3664\,
            in3 => \N__5348\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4076\,
            in2 => \_gnd_net_\,
            in3 => \N__4037\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3895\,
            in1 => \N__3575\,
            in2 => \_gnd_net_\,
            in3 => \N__3604\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__3924\,
            in1 => \N__3891\,
            in2 => \N__3550\,
            in3 => \N__3613\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4071\,
            in1 => \N__4034\,
            in2 => \N__3852\,
            in3 => \N__4094\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3603\,
            in2 => \_gnd_net_\,
            in3 => \N__3571\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIG5942_7_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4095\,
            in1 => \N__4075\,
            in2 => \N__4045\,
            in3 => \N__4035\,
            lcout => \U409_TRANSFER_ACK.N_54_4\,
            ltout => \U409_TRANSFER_ACK.N_54_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__3925\,
            in1 => \N__3892\,
            in2 => \N__4006\,
            in3 => \N__3846\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_5\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000101"
        )
    port map (
            in0 => \N__3893\,
            in1 => \_gnd_net_\,
            in2 => \N__3997\,
            in3 => \N__3802\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__4438\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__3994\,
            in1 => \N__3851\,
            in2 => \N__3985\,
            in3 => \N__3958\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__4425\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIUGMJ1_5_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3926\,
            in1 => \N__3894\,
            in2 => \N__4651\,
            in3 => \N__3850\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a3_0_1_0\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_f0_0_a3_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_0_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__4778\,
            in1 => \_gnd_net_\,
            in2 => \N__3817\,
            in3 => \N__3813\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_i_a3_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3795\,
            in1 => \N__3736\,
            in2 => \N__4604\,
            in3 => \N__3730\,
            lcout => \un1_RAMSPACEn_i_i_a3\,
            ltout => \un1_RAMSPACEn_i_i_a3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.N_11_i_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__4387\,
            in1 => \N__4352\,
            in2 => \N__3715\,
            in3 => \N__4280\,
            lcout => \N_11_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_i_a3_0_a2_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4388\,
            in1 => \N__4353\,
            in2 => \_gnd_net_\,
            in3 => \N__4281\,
            lcout => OPEN,
            ltout => \un1_REGSPACEn_i_i_a3_0_a2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__4471\,
            in1 => \N__4465\,
            in2 => \N__4447\,
            in3 => \N__5365\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.N_52_i_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__4393\,
            in1 => \N__4329\,
            in2 => \_gnd_net_\,
            in3 => \N__4282\,
            lcout => \N_52_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__4657\,
            in1 => \N__4225\,
            in2 => \_gnd_net_\,
            in3 => \N__4858\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5237\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__4213\,
            in1 => \N__4192\,
            in2 => \N__5362\,
            in3 => \N__4171\,
            lcout => \TACK_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            ce => \N__4156\,
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110000"
        )
    port map (
            in0 => \N__4102\,
            in1 => \N__4542\,
            in2 => \N__4134\,
            in3 => \N__4558\,
            lcout => \ROMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            ce => 'H',
            sr => \N__5244\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111100100000"
        )
    port map (
            in0 => \N__4510\,
            in1 => \N__5068\,
            in2 => \N__4552\,
            in3 => \N__4116\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            ce => 'H',
            sr => \N__5244\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5061\,
            in1 => \N__4530\,
            in2 => \N__5105\,
            in3 => \N__5131\,
            lcout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI6OQO2_0_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4498\,
            in1 => \N__4650\,
            in2 => \N__4609\,
            in3 => \N__4773\,
            lcout => \U409_TRANSFER_ACK.N_28_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5130\,
            in1 => \N__5093\,
            in2 => \N__4508\,
            in3 => \N__5060\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__5132\,
            in1 => \N__5094\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_EN_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010111000000"
        )
    port map (
            in0 => \N__4504\,
            in1 => \N__4543\,
            in2 => \N__4531\,
            in3 => \N__5032\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5238\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100001111000"
        )
    port map (
            in0 => \N__5063\,
            in1 => \N__4502\,
            in2 => \N__5106\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5238\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111101110000000"
        )
    port map (
            in0 => \N__5064\,
            in1 => \N__4503\,
            in2 => \N__5107\,
            in3 => \N__5134\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5238\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111010000"
        )
    port map (
            in0 => \N__5133\,
            in1 => \N__5098\,
            in2 => \N__4509\,
            in3 => \N__5062\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__5238\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_1_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4926\,
            in1 => \N__4685\,
            in2 => \N__4912\,
            in3 => \N__4837\,
            lcout => \U409_TRANSFER_ACK.N_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_o2_0_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4908\,
            in2 => \_gnd_net_\,
            in3 => \N__4925\,
            lcout => \U409_TRANSFER_ACK.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__5391\,
            in1 => \N__4680\,
            in2 => \N__4900\,
            in3 => \N__4835\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.N_63_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__4856\,
            in1 => \N__4879\,
            in2 => \N__4873\,
            in3 => \N__4866\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.m9_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5297\,
            in2 => \N__4870\,
            in3 => \N__4813\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000010000"
        )
    port map (
            in0 => \N__4857\,
            in1 => \N__4843\,
            in2 => \N__5315\,
            in3 => \N__4867\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4681\,
            in2 => \_gnd_net_\,
            in3 => \N__4834\,
            lcout => \U409_TRANSFER_ACK.N_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m12_0_a3_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__4836\,
            in1 => \N__4898\,
            in2 => \N__4687\,
            in3 => \N__5393\,
            lcout => \U409_TRANSFER_ACK.N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNIFTON_0_0_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4679\,
            in2 => \_gnd_net_\,
            in3 => \N__4833\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.CIA_STATE_d_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_i_a3_2_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4803\,
            in1 => \N__4897\,
            in2 => \N__4816\,
            in3 => \N__5392\,
            lcout => \U409_TRANSFER_ACK.N_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__4899\,
            in1 => \N__5394\,
            in2 => \N__4807\,
            in3 => \N__4686\,
            lcout => \U409_TRANSFER_ACK.N_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5129\,
            in1 => \N__5092\,
            in2 => \_gnd_net_\,
            in3 => \N__5059\,
            lcout => \U409_TRANSFER_ACK.N_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__5011\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4972\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNI692L_0_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5280\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5158\,
            lcout => \CIA_ENABLE\,
            ltout => \CIA_ENABLE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4966\,
            in3 => \N__4963\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5157\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5281\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__5245\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4927\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__5245\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5395\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \N__5230\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5427\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__5239\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5301\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__5565\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5634\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_2_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5563\,
            in2 => \_gnd_net_\,
            in3 => \N__5733\,
            lcout => OPEN,
            ltout => \U409_CIA.N_93_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_1_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5451\,
            in1 => \N__5473\,
            in2 => \N__5176\,
            in3 => \N__5633\,
            lcout => OPEN,
            ltout => \U409_CIA.VMA_RNOZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__5150\,
            in1 => \N__5564\,
            in2 => \N__5173\,
            in3 => \N__5170\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_1_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__5751\,
            in1 => \N__5732\,
            in2 => \N__5656\,
            in3 => \N__5679\,
            lcout => \U409_CIA.un1_CIA_CLK_COUNT_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIMC921_7_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5651\,
            in1 => \N__5678\,
            in2 => \_gnd_net_\,
            in3 => \N__5750\,
            lcout => \U409_CIA.N_91\,
            ltout => \U409_CIA.N_91_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNICTDR2_0_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5566\,
            in1 => \N__5632\,
            in2 => \N__5137\,
            in3 => \N__5479\,
            lcout => \U409_CIA.CIA_CLK_COUNT11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIBFRM_2_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5769\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5697\,
            lcout => \U409_CIA.CLK_CIA6_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIH7921_2_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5696\,
            in1 => \N__5730\,
            in2 => \_gnd_net_\,
            in3 => \N__5768\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_0_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110001101"
        )
    port map (
            in0 => \N__5542\,
            in1 => \N__5472\,
            in2 => \N__5426\,
            in3 => \N__5731\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA_r_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111011001100"
        )
    port map (
            in0 => \N__5461\,
            in1 => \N__5419\,
            in2 => \N__5455\,
            in3 => \N__5452\,
            lcout => \CLK_CIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_13_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6316\,
            in2 => \_gnd_net_\,
            in3 => \N__5814\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_13_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__6229\,
            in1 => \N__6390\,
            in2 => \N__5491\,
            in3 => \N__6351\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_13_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6475\,
            in1 => \N__6517\,
            in2 => \N__6622\,
            in3 => \N__6562\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_13_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6009\,
            in1 => \N__5972\,
            in2 => \N__5401\,
            in3 => \N__6604\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_13_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__6097\,
            in1 => \N__6133\,
            in2 => \_gnd_net_\,
            in3 => \N__6169\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_13_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5848\,
            in1 => \N__6496\,
            in2 => \N__5398\,
            in3 => \N__6538\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_13_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__5520\,
            in1 => \N__6010\,
            in2 => \N__5536\,
            in3 => \N__5925\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6678\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5810\,
            in2 => \N__6312\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_2_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_13_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5826\,
            in2 => \_gnd_net_\,
            in3 => \N__5509\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__6679\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_13_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6042\,
            in2 => \_gnd_net_\,
            in3 => \N__5506\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__6679\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_13_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6021\,
            in2 => \_gnd_net_\,
            in3 => \N__5503\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_13_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6075\,
            in2 => \_gnd_net_\,
            in3 => \N__5500\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__6679\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_13_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6420\,
            in3 => \N__5497\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_13_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6252\,
            in2 => \_gnd_net_\,
            in3 => \N__5494\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__6679\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_13_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6435\,
            in2 => \_gnd_net_\,
            in3 => \N__5482\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6450\,
            in2 => \_gnd_net_\,
            in3 => \N__5590\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_13_3_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6270\,
            in2 => \_gnd_net_\,
            in3 => \N__5587\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__6681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6063\,
            in2 => \_gnd_net_\,
            in3 => \N__5584\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__6681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5838\,
            in2 => \_gnd_net_\,
            in3 => \N__5581\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__6681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6282\,
            in2 => \_gnd_net_\,
            in3 => \N__5578\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__6681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6402\,
            in2 => \_gnd_net_\,
            in3 => \N__5575\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_13_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6240\,
            in2 => \_gnd_net_\,
            in3 => \N__5572\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_13_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5794\,
            in2 => \_gnd_net_\,
            in3 => \N__5569\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6681\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_2_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__5627\,
            in1 => \N__5562\,
            in2 => \N__5635\,
            in3 => \_gnd_net_\,
            lcout => \U409_CIA.CLK_CIA6_1\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5770\,
            in2 => \_gnd_net_\,
            in3 => \N__5755\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__5604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5706\,
            in1 => \N__5752\,
            in2 => \_gnd_net_\,
            in3 => \N__5737\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \N__5604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5734\,
            in2 => \_gnd_net_\,
            in3 => \N__5710\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__5604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5707\,
            in1 => \N__5698\,
            in2 => \_gnd_net_\,
            in3 => \N__5683\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            clk => \N__5604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_6_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5680\,
            in2 => \_gnd_net_\,
            in3 => \N__5662\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\,
            clk => \N__5604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_7_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5655\,
            in2 => \_gnd_net_\,
            in3 => \N__5659\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5631\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_14_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__6003\,
            in1 => \N__5969\,
            in2 => \N__6175\,
            in3 => \N__5926\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_14_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5968\,
            in1 => \N__6006\,
            in2 => \N__5938\,
            in3 => \N__6085\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_14_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__6004\,
            in1 => \N__5970\,
            in2 => \N__6733\,
            in3 => \N__5927\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_14_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5967\,
            in1 => \N__6005\,
            in2 => \N__5937\,
            in3 => \N__6709\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6577\,
            in1 => \N__6148\,
            in2 => \N__6193\,
            in3 => \N__6696\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_14_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6592\,
            in1 => \N__6745\,
            in2 => \N__6115\,
            in3 => \N__6721\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_14_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__6547\,
            in1 => \N__5971\,
            in2 => \N__5842\,
            in3 => \N__5934\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_14_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6170\,
            in2 => \_gnd_net_\,
            in3 => \N__6192\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6680\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_14_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5839\,
            in1 => \N__5827\,
            in2 => \N__5815\,
            in3 => \N__5793\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_14_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__6388\,
            in1 => \N__6350\,
            in2 => \N__5782\,
            in3 => \N__6228\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_14_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__6007\,
            in1 => \N__6505\,
            in2 => \N__5977\,
            in3 => \N__5935\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_14_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6076\,
            in1 => \N__6022\,
            in2 => \_gnd_net_\,
            in3 => \N__6307\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_14_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6064\,
            in1 => \N__6052\,
            in2 => \N__6046\,
            in3 => \N__6043\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_14_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__6387\,
            in1 => \N__6226\,
            in2 => \N__6031\,
            in3 => \N__6028\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_14_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__6008\,
            in1 => \N__5976\,
            in2 => \N__6463\,
            in3 => \N__5936\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_14_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__6389\,
            in1 => \N__5886\,
            in2 => \N__6355\,
            in3 => \N__6227\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6682\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__6347\,
            in1 => \N__6224\,
            in2 => \N__5875\,
            in3 => \N__6385\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_14_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__6222\,
            in1 => \N__5863\,
            in2 => \N__6391\,
            in3 => \N__6349\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_14_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__6348\,
            in1 => \N__6225\,
            in2 => \N__5857\,
            in3 => \N__6386\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_14_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6451\,
            in1 => \N__6439\,
            in2 => \N__6424\,
            in3 => \N__6403\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_14_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__6346\,
            in1 => \N__6223\,
            in2 => \N__6319\,
            in3 => \N__6311\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6684\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_14_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__6283\,
            in1 => \N__6271\,
            in2 => \N__6259\,
            in3 => \N__6241\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6188\,
            in2 => \N__6174\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_1_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_15_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6147\,
            in2 => \_gnd_net_\,
            in3 => \N__6136\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__6683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_15_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6129\,
            in2 => \_gnd_net_\,
            in3 => \N__6118\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__6683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_15_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6111\,
            in2 => \_gnd_net_\,
            in3 => \N__6100\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__6683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_15_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6096\,
            in2 => \_gnd_net_\,
            in3 => \N__6079\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_15_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6621\,
            in2 => \_gnd_net_\,
            in3 => \N__6595\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_15_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6591\,
            in2 => \_gnd_net_\,
            in3 => \N__6580\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__6683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_15_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6576\,
            in2 => \_gnd_net_\,
            in3 => \N__6565\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__6683\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_15_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6558\,
            in2 => \_gnd_net_\,
            in3 => \N__6541\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_2_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_15_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6531\,
            in2 => \_gnd_net_\,
            in3 => \N__6520\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__6685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_15_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6516\,
            in2 => \_gnd_net_\,
            in3 => \N__6499\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_15_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6489\,
            in2 => \_gnd_net_\,
            in3 => \N__6478\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__6685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_15_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6474\,
            in2 => \_gnd_net_\,
            in3 => \N__6454\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_15_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6744\,
            in2 => \_gnd_net_\,
            in3 => \N__6724\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_15_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6720\,
            in2 => \_gnd_net_\,
            in3 => \N__6703\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_15_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6697\,
            in2 => \_gnd_net_\,
            in3 => \N__6700\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6685\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_iobuf_RNO_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6655\,
            lcout => \N_525_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 14 2025 00:16:40

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    TM : in std_logic_vector(1 downto 0);
    TT : in std_logic_vector(1 downto 0);
    D : inout std_logic_vector(7 downto 4);
    A : in std_logic_vector(31 downto 1);
    PIO_S0 : out std_logic;
    PORTSIZE : out std_logic;
    TICK60 : out std_logic;
    CIACS0n : out std_logic;
    CPUCONFn : in std_logic;
    CLK6 : in std_logic;
    CLK_CIA : out std_logic;
    BUFENn : out std_logic;
    AUTOBOOT : in std_logic;
    RnW : in std_logic;
    PIO_P2 : out std_logic;
    CIACS1n : out std_logic;
    BRIDGE_ENn : out std_logic;
    PIO_S1 : out std_logic;
    PIO_P0 : out std_logic;
    TICK50 : out std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : out std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    REGSPACEn : out std_logic;
    TSn : in std_logic;
    RTC_ENn : out std_logic;
    PIO_S2 : out std_logic;
    ATA_ENn : out std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    CONFIGENn : out std_logic;
    TACKn : inout std_logic;
    ROMENn : out std_logic;
    PIO_P1 : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__3990\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_14\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_a3_0Z0Z_2_cascade_\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4_cascade_\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_27\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_5\ : std_logic;
signal \U409_AUTOCONFIG.N_42\ : std_logic;
signal \U409_AUTOCONFIG.N_111_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_1_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_62\ : std_logic;
signal \U409_ADDRESS_DECODE.N_54_cascade_\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U409_AUTOCONFIG.N_92\ : std_logic;
signal \U409_AUTOCONFIG.N_86_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_57\ : std_logic;
signal \N_89_1\ : std_logic;
signal \N_89_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_3\ : std_logic;
signal \A_c_25\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_9\ : std_logic;
signal \U409_AUTOCONFIG.N_38\ : std_logic;
signal \U409_AUTOCONFIG.N_48\ : std_logic;
signal \U409_AUTOCONFIG.N_111\ : std_logic;
signal \U409_AUTOCONFIG.N_41\ : std_logic;
signal \U409_AUTOCONFIG.N_43\ : std_logic;
signal \U409_AUTOCONFIG.N_66\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_i_1_cascade_\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_OUT_3C_net\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.N_112_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.N_112\ : std_logic;
signal \U409_AUTOCONFIG.N_74_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_i_0\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U409_AUTOCONFIG.N_44\ : std_logic;
signal \U409_AUTOCONFIG.N_86\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_85_i_i_0\ : std_logic;
signal \N_121\ : std_logic;
signal \N_121_cascade_\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_7\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG_D_OUT_0_i_0\ : std_logic;
signal \U409_AUTOCONFIG.N_27\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.N_31\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\ : std_logic;
signal \U409_AUTOCONFIG.N_22\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONF_1_sqmuxa_0_a2_0Z0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.N_20\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net\ : std_logic;
signal \CPUCONFn_c\ : std_logic;
signal \U409_AUTOCONFIG.N_52\ : std_logic;
signal \U409_AUTOCONFIG.N_52_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_56\ : std_logic;
signal \U409_AUTOCONFIG.N_67\ : std_logic;
signal \U409_AUTOCONFIG.N_56_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0Z0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa\ : std_logic;
signal \U409_ADDRESS_DECODE.HIROMZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.LOWROMZ0Z_2_cascade_\ : std_logic;
signal \D_1_i\ : std_logic;
signal \U409_AUTOCONFIG.AC_STARTZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_1_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_10\ : std_logic;
signal \N_120_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_11\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn_i\ : std_logic;
signal \U409_ADDRESS_DECODE.N_102\ : std_logic;
signal \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3Z0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG_D_OUT_0_i_1\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG_D_OUT_0_i_2\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG_D_OUT_0_i_3\ : std_logic;
signal \U409_AUTOCONFIG.STATEZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.STATEZ0Z_0\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_CONFC_net\ : std_logic;
signal \TM_c_0\ : std_logic;
signal \CONFIGURED\ : std_logic;
signal \TM_c_1\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_\ : std_logic;
signal \ATA_BASE_1\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACE\ : std_logic;
signal \N_120_i\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1\ : std_logic;
signal \A_c_31\ : std_logic;
signal \N_120\ : std_logic;
signal \U409_ADDRESS_DECODE.PORTSIZEZ0Z_0_cascade_\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_29\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_0\ : std_logic;
signal \CONFIGENn_c\ : std_logic;
signal \D_in_7\ : std_logic;
signal \BRIDGE_BASE_3\ : std_logic;
signal \BRIDGE_BASE_2\ : std_logic;
signal \BRIDGE_BASE_1\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\ : std_logic;
signal \INVU409_AUTOCONFIG.CONFIGENnC_net\ : std_logic;
signal \A_c_23\ : std_logic;
signal \ATA_BASE_7\ : std_logic;
signal \A_c_22\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\ : std_logic;
signal \A_c_1\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONFZ0\ : std_logic;
signal \U409_AUTOCONFIG.N_122\ : std_logic;
signal \A_c_19\ : std_logic;
signal \ATA_BASE_3\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACE_1Z0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_ROMEN_0\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_ENZ0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_ATA_ENn_i\ : std_logic;
signal \U409_TRANSFER_ACK.CO1\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_cascade_\ : std_logic;
signal \D_in_4\ : std_logic;
signal \ATA_BASE_4\ : std_logic;
signal \D_in_5\ : std_logic;
signal \ATA_BASE_5\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_1\ : std_logic;
signal \ATA_BASE_6\ : std_logic;
signal \INVU409_AUTOCONFIG.ATA_BASE_4C_net\ : std_logic;
signal \un1_AUTOCONFIG_SPACE\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_0\ : std_logic;
signal \D_in_6\ : std_logic;
signal \ATA_BASE_2\ : std_logic;
signal \INVU409_AUTOCONFIG.ATA_BASE_2C_net\ : std_logic;
signal \U409_ADDRESS_DECODE.LOWROMZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE_ROMEN_1\ : std_logic;
signal \A_c_21\ : std_logic;
signal \OVL_c\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\ : std_logic;
signal \A_c_28\ : std_logic;
signal \BRIDGE_BASE_0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \ROMENn_c\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROMENn_nessC_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_ENC_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_OUTnC_net\ : std_logic;
signal \AC_TACK\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_OUTn_3_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_2\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn\ : std_logic;
signal \BUFENn_c\ : std_logic;
signal \U409_TRANSFER_ACK.N_119\ : std_logic;
signal \GB_BUFFER_CLK40_IN_c_g_THRU_CO\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U409_TRANSFER_ACK.N_17_mux_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_6_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_3_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_17_mux\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a3_3\ : std_logic;
signal \U409_TRANSFER_ACK.N_87_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_77\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\ : std_logic;
signal \TSn_c\ : std_logic;
signal \CLK40_IN_c_g\ : std_logic;
signal \U409_TRANSFER_ACK.N_87\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.TICK603_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_1C_net\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \U409_CIA.CLK_CIA_r_1_0_cascade_\ : std_logic;
signal \CLK_CIA_c\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \U409_CIA.CLK_CIA6_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_3_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\ : std_logic;
signal \U409_CIA.CLK_CIA6_4_cascade_\ : std_logic;
signal \U409_CIA.VMA_RNOZ0Z_0_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \bfn_16_7_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_6\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_6\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_7\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_3_2\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \AUTOCONFIG_SPACE\ : std_logic;
signal \CIA_SPACE\ : std_logic;
signal \TCIn_1_i\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \CIA_ENABLE\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \PIO_P1_wire\ : std_logic;
signal \CPUCONFn_wire\ : std_logic;
signal \RTC_ENn_wire\ : std_logic;
signal \TM_wire\ : std_logic_vector(1 downto 0);
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \PIO_P2_wire\ : std_logic;
signal \BRIDGE_ENn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CONFIGENn_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \PIO_P0_wire\ : std_logic;
signal \ATA_ENn_wire\ : std_logic;
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \CLK_CIA_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \PIO_S0_wire\ : std_logic;
signal \PIO_S2_wire\ : std_logic;
signal \PIO_S1_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    \CLK40_IN_wire\ <= CLK40_IN;
    \A_wire\ <= A;
    \TT_wire\ <= TT;
    PIO_P1 <= \PIO_P1_wire\;
    \CPUCONFn_wire\ <= CPUCONFn;
    RTC_ENn <= \RTC_ENn_wire\;
    \TM_wire\ <= TM;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    TBIn <= \TBIn_wire\;
    \TSn_wire\ <= TSn;
    PORTSIZE <= \PORTSIZE_wire\;
    PIO_P2 <= \PIO_P2_wire\;
    BRIDGE_ENn <= \BRIDGE_ENn_wire\;
    \RESETn_wire\ <= RESETn;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TCIn <= \TCIn_wire\;
    \RnW_wire\ <= RnW;
    CONFIGENn <= \CONFIGENn_wire\;
    TICK60 <= \TICK60_wire\;
    PIO_P0 <= \PIO_P0_wire\;
    ATA_ENn <= \ATA_ENn_wire\;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    CLK_CIA <= \CLK_CIA_wire\;
    BUFENn <= \BUFENn_wire\;
    PIO_S0 <= \PIO_S0_wire\;
    PIO_S2 <= \PIO_S2_wire\;
    PIO_S1 <= \PIO_S1_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__7680\,
            RESETB => \N__7665\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11322\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11324\,
            DIN => \N__11323\,
            DOUT => \N__11322\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11324\,
            PADOUT => \N__11323\,
            PADIN => \N__11322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11312\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11314\,
            DIN => \N__11313\,
            DOUT => \N__11312\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11314\,
            PADOUT => \N__11313\,
            PADIN => \N__11312\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11302\,
            GLOBALBUFFEROUTPUT => \CLK40_IN_c_g\
        );

    \CLK40_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11304\,
            DIN => \N__11303\,
            DOUT => \N__11302\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11304\,
            PADOUT => \N__11303\,
            PADIN => \N__11302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11293\,
            DIN => \N__11292\,
            DOUT => \N__11291\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11293\,
            PADOUT => \N__11292\,
            PADIN => \N__11291\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11284\,
            DIN => \N__11283\,
            DOUT => \N__11282\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11284\,
            PADOUT => \N__11283\,
            PADIN => \N__11282\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_P1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11275\,
            DIN => \N__11274\,
            DOUT => \N__11273\,
            PACKAGEPIN => \PIO_P1_wire\
        );

    \PIO_P1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11275\,
            PADOUT => \N__11274\,
            PADIN => \N__11273\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10647\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11266\,
            DIN => \N__11265\,
            DOUT => \N__11264\,
            PACKAGEPIN => D(7)
        );

    \D_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11266\,
            PADOUT => \N__11265\,
            PADIN => \N__11264\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5160\,
            DIN0 => \D_in_7\,
            DOUT0 => \N__5223\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11257\,
            DIN => \N__11256\,
            DOUT => \N__11255\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11257\,
            PADOUT => \N__11256\,
            PADIN => \N__11255\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUCONFn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11248\,
            DIN => \N__11247\,
            DOUT => \N__11246\,
            PACKAGEPIN => \CPUCONFn_wire\
        );

    \CPUCONFn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11248\,
            PADOUT => \N__11247\,
            PADIN => \N__11246\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CPUCONFn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RTC_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11239\,
            DIN => \N__11238\,
            DOUT => \N__11237\,
            PACKAGEPIN => \RTC_ENn_wire\
        );

    \RTC_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11239\,
            PADOUT => \N__11238\,
            PADIN => \N__11237\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5427\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11230\,
            DIN => \N__11229\,
            DOUT => \N__11228\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11230\,
            PADOUT => \N__11229\,
            PADIN => \N__11228\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11221\,
            DIN => \N__11220\,
            DOUT => \N__11219\,
            PACKAGEPIN => D(4)
        );

    \D_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11221\,
            PADOUT => \N__11220\,
            PADIN => \N__11219\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5135\,
            DIN0 => \D_in_4\,
            DOUT0 => \N__4530\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11212\,
            DIN => \N__11211\,
            DOUT => \N__11210\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11212\,
            PADOUT => \N__11211\,
            PADIN => \N__11210\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11203\,
            DIN => \N__11202\,
            DOUT => \N__11201\,
            PACKAGEPIN => \TM_wire\(1)
        );

    \TM_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11203\,
            PADOUT => \N__11202\,
            PADIN => \N__11201\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11194\,
            DIN => \N__11193\,
            DOUT => \N__11192\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11194\,
            PADOUT => \N__11193\,
            PADIN => \N__11192\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11185\,
            DIN => \N__11184\,
            DOUT => \N__11183\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11185\,
            PADOUT => \N__11184\,
            PADIN => \N__11183\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6840\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11176\,
            DIN => \N__11175\,
            DOUT => \N__11174\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11176\,
            PADOUT => \N__11175\,
            PADIN => \N__11174\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11167\,
            DIN => \N__11166\,
            DOUT => \N__11165\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11167\,
            PADOUT => \N__11166\,
            PADIN => \N__11165\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7578\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11158\,
            DIN => \N__11157\,
            DOUT => \N__11156\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11158\,
            PADOUT => \N__11157\,
            PADIN => \N__11156\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10359\,
            DIN0 => OPEN,
            DOUT0 => \N__7982\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11149\,
            DIN => \N__11148\,
            DOUT => \N__11147\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11149\,
            PADOUT => \N__11148\,
            PADIN => \N__11147\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11140\,
            DIN => \N__11139\,
            DOUT => \N__11138\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11140\,
            PADOUT => \N__11139\,
            PADIN => \N__11138\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5928\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_P2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11131\,
            DIN => \N__11130\,
            DOUT => \N__11129\,
            PACKAGEPIN => \PIO_P2_wire\
        );

    \PIO_P2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11131\,
            PADOUT => \N__11130\,
            PADIN => \N__11129\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4056\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11122\,
            DIN => \N__11121\,
            DOUT => \N__11120\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11122\,
            PADOUT => \N__11121\,
            PADIN => \N__11120\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BRIDGE_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11113\,
            DIN => \N__11112\,
            DOUT => \N__11111\,
            PACKAGEPIN => \BRIDGE_ENn_wire\
        );

    \BRIDGE_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11113\,
            PADOUT => \N__11112\,
            PADIN => \N__11111\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6957\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11104\,
            DIN => \N__11103\,
            DOUT => \N__11102\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11104\,
            PADOUT => \N__11103\,
            PADIN => \N__11102\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11095\,
            DIN => \N__11094\,
            DOUT => \N__11093\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11095\,
            PADOUT => \N__11094\,
            PADIN => \N__11093\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11086\,
            DIN => \N__11085\,
            DOUT => \N__11084\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11086\,
            PADOUT => \N__11085\,
            PADIN => \N__11084\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11077\,
            DIN => \N__11076\,
            DOUT => \N__11075\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11077\,
            PADOUT => \N__11076\,
            PADIN => \N__11075\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11068\,
            DIN => \N__11067\,
            DOUT => \N__11066\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11068\,
            PADOUT => \N__11067\,
            PADIN => \N__11066\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11059\,
            DIN => \N__11058\,
            DOUT => \N__11057\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11059\,
            PADOUT => \N__11058\,
            PADIN => \N__11057\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11050\,
            DIN => \N__11049\,
            DOUT => \N__11048\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11050\,
            PADOUT => \N__11049\,
            PADIN => \N__11048\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10674\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11041\,
            DIN => \N__11040\,
            DOUT => \N__11039\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11041\,
            PADOUT => \N__11040\,
            PADIN => \N__11039\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9459\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11032\,
            DIN => \N__11031\,
            DOUT => \N__11030\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11032\,
            PADOUT => \N__11031\,
            PADIN => \N__11030\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11023\,
            DIN => \N__11022\,
            DOUT => \N__11021\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11023\,
            PADOUT => \N__11022\,
            PADIN => \N__11021\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11014\,
            DIN => \N__11013\,
            DOUT => \N__11012\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11014\,
            PADOUT => \N__11013\,
            PADIN => \N__11012\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11005\,
            DIN => \N__11004\,
            DOUT => \N__11003\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11005\,
            PADOUT => \N__11004\,
            PADIN => \N__11003\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10996\,
            DIN => \N__10995\,
            DOUT => \N__10994\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__10996\,
            PADOUT => \N__10995\,
            PADIN => \N__10994\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10212\,
            DIN0 => OPEN,
            DOUT0 => \N__7983\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10987\,
            DIN => \N__10986\,
            DOUT => \N__10985\,
            PACKAGEPIN => D(5)
        );

    \D_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__10987\,
            PADOUT => \N__10986\,
            PADIN => \N__10985\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5155\,
            DIN0 => \D_in_5\,
            DOUT0 => \N__5316\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10978\,
            DIN => \N__10977\,
            DOUT => \N__10976\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10978\,
            PADOUT => \N__10977\,
            PADIN => \N__10976\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10969\,
            DIN => \N__10968\,
            DOUT => \N__10967\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10969\,
            PADOUT => \N__10968\,
            PADIN => \N__10967\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10960\,
            DIN => \N__10959\,
            DOUT => \N__10958\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10960\,
            PADOUT => \N__10959\,
            PADIN => \N__10958\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CONFIGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10951\,
            DIN => \N__10950\,
            DOUT => \N__10949\,
            PACKAGEPIN => \CONFIGENn_wire\
        );

    \CONFIGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10951\,
            PADOUT => \N__10950\,
            PADIN => \N__10949\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5814\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10942\,
            DIN => \N__10941\,
            DOUT => \N__10940\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10942\,
            PADOUT => \N__10941\,
            PADIN => \N__10940\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9291\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10933\,
            DIN => \N__10932\,
            DOUT => \N__10931\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10933\,
            PADOUT => \N__10932\,
            PADIN => \N__10931\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_P0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10924\,
            DIN => \N__10923\,
            DOUT => \N__10922\,
            PACKAGEPIN => \PIO_P0_wire\
        );

    \PIO_P0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10924\,
            PADOUT => \N__10923\,
            PADIN => \N__10922\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10716\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10915\,
            DIN => \N__10914\,
            DOUT => \N__10913\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10915\,
            PADOUT => \N__10914\,
            PADIN => \N__10913\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10906\,
            DIN => \N__10905\,
            DOUT => \N__10904\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10906\,
            PADOUT => \N__10905\,
            PADIN => \N__10904\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ATA_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10897\,
            DIN => \N__10896\,
            DOUT => \N__10895\,
            PACKAGEPIN => \ATA_ENn_wire\
        );

    \ATA_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10897\,
            PADOUT => \N__10896\,
            PADIN => \N__10895\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6789\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10888\,
            DIN => \N__10887\,
            DOUT => \N__10886\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10888\,
            PADOUT => \N__10887\,
            PADIN => \N__10886\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10879\,
            DIN => \N__10878\,
            DOUT => \N__10877\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10879\,
            PADOUT => \N__10878\,
            PADIN => \N__10877\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10611\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10870\,
            DIN => \N__10869\,
            DOUT => \N__10868\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10870\,
            PADOUT => \N__10869\,
            PADIN => \N__10868\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5400\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10861\,
            DIN => \N__10860\,
            DOUT => \N__10859\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10861\,
            PADOUT => \N__10860\,
            PADIN => \N__10859\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_CIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10852\,
            DIN => \N__10851\,
            DOUT => \N__10850\,
            PACKAGEPIN => \CLK_CIA_wire\
        );

    \CLK_CIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10852\,
            PADOUT => \N__10851\,
            PADIN => \N__10850\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9213\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10843\,
            DIN => \N__10842\,
            DOUT => \N__10841\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10843\,
            PADOUT => \N__10842\,
            PADIN => \N__10841\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10834\,
            DIN => \N__10833\,
            DOUT => \N__10832\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__10834\,
            PADOUT => \N__10833\,
            PADIN => \N__10832\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10355\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__7975\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10825\,
            DIN => \N__10824\,
            DOUT => \N__10823\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10825\,
            PADOUT => \N__10824\,
            PADIN => \N__10823\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10816\,
            DIN => \N__10815\,
            DOUT => \N__10814\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10816\,
            PADOUT => \N__10815\,
            PADIN => \N__10814\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7704\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_S0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10807\,
            DIN => \N__10806\,
            DOUT => \N__10805\,
            PACKAGEPIN => \PIO_S0_wire\
        );

    \PIO_S0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10807\,
            PADOUT => \N__10806\,
            PADIN => \N__10805\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4080\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10798\,
            DIN => \N__10797\,
            DOUT => \N__10796\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10798\,
            PADOUT => \N__10797\,
            PADIN => \N__10796\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_S2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10789\,
            DIN => \N__10788\,
            DOUT => \N__10787\,
            PACKAGEPIN => \PIO_S2_wire\
        );

    \PIO_S2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10789\,
            PADOUT => \N__10788\,
            PADIN => \N__10787\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7664\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10780\,
            DIN => \N__10779\,
            DOUT => \N__10778\,
            PACKAGEPIN => D(6)
        );

    \D_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__10780\,
            PADOUT => \N__10779\,
            PADIN => \N__10778\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5156\,
            DIN0 => \D_in_6\,
            DOUT0 => \N__5268\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10771\,
            DIN => \N__10770\,
            DOUT => \N__10769\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10771\,
            PADOUT => \N__10770\,
            PADIN => \N__10769\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10762\,
            DIN => \N__10761\,
            DOUT => \N__10760\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10762\,
            PADOUT => \N__10761\,
            PADIN => \N__10760\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_S1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10753\,
            DIN => \N__10752\,
            DOUT => \N__10751\,
            PACKAGEPIN => \PIO_S1_wire\
        );

    \PIO_S1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10753\,
            PADOUT => \N__10752\,
            PADIN => \N__10751\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4638\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10744\,
            DIN => \N__10743\,
            DOUT => \N__10742\,
            PACKAGEPIN => \TM_wire\(0)
        );

    \TM_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10744\,
            PADOUT => \N__10743\,
            PADIN => \N__10742\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10735\,
            DIN => \N__10734\,
            DOUT => \N__10733\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10735\,
            PADOUT => \N__10734\,
            PADIN => \N__10733\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2593\ : IoInMux
    port map (
            O => \N__10716\,
            I => \N__10713\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__10713\,
            I => \N__10710\
        );

    \I__2591\ : Span4Mux_s0_h
    port map (
            O => \N__10710\,
            I => \N__10706\
        );

    \I__2590\ : InMux
    port map (
            O => \N__10709\,
            I => \N__10703\
        );

    \I__2589\ : Sp12to4
    port map (
            O => \N__10706\,
            I => \N__10700\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__10703\,
            I => \N__10697\
        );

    \I__2587\ : Span12Mux_s10_v
    port map (
            O => \N__10700\,
            I => \N__10694\
        );

    \I__2586\ : Span12Mux_s10_v
    port map (
            O => \N__10697\,
            I => \N__10691\
        );

    \I__2585\ : Span12Mux_h
    port map (
            O => \N__10694\,
            I => \N__10688\
        );

    \I__2584\ : Span12Mux_h
    port map (
            O => \N__10691\,
            I => \N__10685\
        );

    \I__2583\ : Span12Mux_h
    port map (
            O => \N__10688\,
            I => \N__10682\
        );

    \I__2582\ : Span12Mux_h
    port map (
            O => \N__10685\,
            I => \N__10679\
        );

    \I__2581\ : Odrv12
    port map (
            O => \N__10682\,
            I => \A_c_12\
        );

    \I__2580\ : Odrv12
    port map (
            O => \N__10679\,
            I => \A_c_12\
        );

    \I__2579\ : IoInMux
    port map (
            O => \N__10674\,
            I => \N__10671\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__10671\,
            I => \N__10668\
        );

    \I__2577\ : Span4Mux_s3_h
    port map (
            O => \N__10668\,
            I => \N__10665\
        );

    \I__2576\ : Span4Mux_v
    port map (
            O => \N__10665\,
            I => \N__10662\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__10662\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__2574\ : InMux
    port map (
            O => \N__10659\,
            I => \N__10653\
        );

    \I__2573\ : InMux
    port map (
            O => \N__10658\,
            I => \N__10653\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__10653\,
            I => \N__10650\
        );

    \I__2571\ : Odrv12
    port map (
            O => \N__10650\,
            I => \CIA_ENABLE\
        );

    \I__2570\ : IoInMux
    port map (
            O => \N__10647\,
            I => \N__10644\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__10644\,
            I => \N__10641\
        );

    \I__2568\ : IoSpan4Mux
    port map (
            O => \N__10641\,
            I => \N__10637\
        );

    \I__2567\ : InMux
    port map (
            O => \N__10640\,
            I => \N__10634\
        );

    \I__2566\ : IoSpan4Mux
    port map (
            O => \N__10637\,
            I => \N__10631\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__10634\,
            I => \N__10628\
        );

    \I__2564\ : Span4Mux_s3_h
    port map (
            O => \N__10631\,
            I => \N__10623\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__10628\,
            I => \N__10623\
        );

    \I__2562\ : Sp12to4
    port map (
            O => \N__10623\,
            I => \N__10620\
        );

    \I__2561\ : Span12Mux_h
    port map (
            O => \N__10620\,
            I => \N__10617\
        );

    \I__2560\ : Span12Mux_h
    port map (
            O => \N__10617\,
            I => \N__10614\
        );

    \I__2559\ : Odrv12
    port map (
            O => \N__10614\,
            I => \A_c_13\
        );

    \I__2558\ : IoInMux
    port map (
            O => \N__10611\,
            I => \N__10608\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__10608\,
            I => \N__10605\
        );

    \I__2556\ : Span4Mux_s3_h
    port map (
            O => \N__10605\,
            I => \N__10602\
        );

    \I__2555\ : Span4Mux_v
    port map (
            O => \N__10602\,
            I => \N__10599\
        );

    \I__2554\ : Odrv4
    port map (
            O => \N__10599\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__2553\ : InMux
    port map (
            O => \N__10596\,
            I => \N__10593\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10593\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\
        );

    \I__2551\ : InMux
    port map (
            O => \N__10590\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__2550\ : InMux
    port map (
            O => \N__10587\,
            I => \N__10584\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__10584\,
            I => \N__10578\
        );

    \I__2548\ : InMux
    port map (
            O => \N__10583\,
            I => \N__10575\
        );

    \I__2547\ : InMux
    port map (
            O => \N__10582\,
            I => \N__10572\
        );

    \I__2546\ : InMux
    port map (
            O => \N__10581\,
            I => \N__10569\
        );

    \I__2545\ : Odrv4
    port map (
            O => \N__10578\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__10575\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__10572\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__10569\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2541\ : InMux
    port map (
            O => \N__10560\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__2540\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10554\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__10554\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO\
        );

    \I__2538\ : InMux
    port map (
            O => \N__10551\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__2537\ : InMux
    port map (
            O => \N__10548\,
            I => \N__10542\
        );

    \I__2536\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10539\
        );

    \I__2535\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10536\
        );

    \I__2534\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10533\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10542\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__10539\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__10536\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__10533\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__2529\ : InMux
    port map (
            O => \N__10524\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\
        );

    \I__2528\ : InMux
    port map (
            O => \N__10521\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__10518\,
            I => \N__10512\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__10517\,
            I => \N__10509\
        );

    \I__2525\ : InMux
    port map (
            O => \N__10516\,
            I => \N__10506\
        );

    \I__2524\ : InMux
    port map (
            O => \N__10515\,
            I => \N__10503\
        );

    \I__2523\ : InMux
    port map (
            O => \N__10512\,
            I => \N__10498\
        );

    \I__2522\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10498\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__10506\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__10503\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__10498\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__2518\ : ClkMux
    port map (
            O => \N__10491\,
            I => \N__10479\
        );

    \I__2517\ : ClkMux
    port map (
            O => \N__10490\,
            I => \N__10479\
        );

    \I__2516\ : ClkMux
    port map (
            O => \N__10489\,
            I => \N__10479\
        );

    \I__2515\ : ClkMux
    port map (
            O => \N__10488\,
            I => \N__10479\
        );

    \I__2514\ : GlobalMux
    port map (
            O => \N__10479\,
            I => \N__10476\
        );

    \I__2513\ : gio2CtrlBuf
    port map (
            O => \N__10476\,
            I => \CLK28_IN_c_g\
        );

    \I__2512\ : InMux
    port map (
            O => \N__10473\,
            I => \N__10466\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10461\
        );

    \I__2510\ : InMux
    port map (
            O => \N__10471\,
            I => \N__10461\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10470\,
            I => \N__10456\
        );

    \I__2508\ : InMux
    port map (
            O => \N__10469\,
            I => \N__10456\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__10466\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__10461\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__10456\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__2504\ : InMux
    port map (
            O => \N__10449\,
            I => \N__10446\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10446\,
            I => \N__10440\
        );

    \I__2502\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10437\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10444\,
            I => \N__10432\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10432\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__10440\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__10437\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__10432\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__2496\ : CascadeMux
    port map (
            O => \N__10425\,
            I => \N__10419\
        );

    \I__2495\ : CascadeMux
    port map (
            O => \N__10424\,
            I => \N__10415\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10423\,
            I => \N__10412\
        );

    \I__2493\ : InMux
    port map (
            O => \N__10422\,
            I => \N__10407\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10407\
        );

    \I__2491\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10402\
        );

    \I__2490\ : InMux
    port map (
            O => \N__10415\,
            I => \N__10402\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__10412\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__10407\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__10402\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__10395\,
            I => \N__10387\
        );

    \I__2485\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10384\
        );

    \I__2484\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10377\
        );

    \I__2483\ : InMux
    port map (
            O => \N__10392\,
            I => \N__10377\
        );

    \I__2482\ : InMux
    port map (
            O => \N__10391\,
            I => \N__10377\
        );

    \I__2481\ : InMux
    port map (
            O => \N__10390\,
            I => \N__10372\
        );

    \I__2480\ : InMux
    port map (
            O => \N__10387\,
            I => \N__10372\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__10384\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__10377\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__10372\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2476\ : InMux
    port map (
            O => \N__10365\,
            I => \N__10362\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__10362\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_3_2\
        );

    \I__2474\ : IoInMux
    port map (
            O => \N__10359\,
            I => \N__10356\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__10356\,
            I => \N__10352\
        );

    \I__2472\ : IoInMux
    port map (
            O => \N__10355\,
            I => \N__10349\
        );

    \I__2471\ : IoSpan4Mux
    port map (
            O => \N__10352\,
            I => \N__10346\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__10349\,
            I => \N__10343\
        );

    \I__2469\ : Span4Mux_s0_v
    port map (
            O => \N__10346\,
            I => \N__10338\
        );

    \I__2468\ : Span4Mux_s0_v
    port map (
            O => \N__10343\,
            I => \N__10338\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__10338\,
            I => \N__10334\
        );

    \I__2466\ : InMux
    port map (
            O => \N__10337\,
            I => \N__10331\
        );

    \I__2465\ : Sp12to4
    port map (
            O => \N__10334\,
            I => \N__10328\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__10331\,
            I => \N__10325\
        );

    \I__2463\ : Span12Mux_s9_h
    port map (
            O => \N__10328\,
            I => \N__10321\
        );

    \I__2462\ : Span4Mux_v
    port map (
            O => \N__10325\,
            I => \N__10318\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__10324\,
            I => \N__10315\
        );

    \I__2460\ : Span12Mux_v
    port map (
            O => \N__10321\,
            I => \N__10312\
        );

    \I__2459\ : Span4Mux_h
    port map (
            O => \N__10318\,
            I => \N__10309\
        );

    \I__2458\ : InMux
    port map (
            O => \N__10315\,
            I => \N__10306\
        );

    \I__2457\ : Odrv12
    port map (
            O => \N__10312\,
            I => \TACK_EN\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__10309\,
            I => \TACK_EN\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__10306\,
            I => \TACK_EN\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10299\,
            I => \N__10296\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__10296\,
            I => \N__10292\
        );

    \I__2452\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10289\
        );

    \I__2451\ : Span4Mux_h
    port map (
            O => \N__10292\,
            I => \N__10283\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10289\,
            I => \N__10283\
        );

    \I__2449\ : InMux
    port map (
            O => \N__10288\,
            I => \N__10280\
        );

    \I__2448\ : Span4Mux_h
    port map (
            O => \N__10283\,
            I => \N__10276\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__10280\,
            I => \N__10273\
        );

    \I__2446\ : InMux
    port map (
            O => \N__10279\,
            I => \N__10270\
        );

    \I__2445\ : Span4Mux_h
    port map (
            O => \N__10276\,
            I => \N__10265\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__10273\,
            I => \N__10260\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__10270\,
            I => \N__10260\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10269\,
            I => \N__10255\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10255\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__10265\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__2439\ : Odrv4
    port map (
            O => \N__10260\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__10255\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10248\,
            I => \N__10245\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__10245\,
            I => \N__10242\
        );

    \I__2435\ : Span4Mux_v
    port map (
            O => \N__10242\,
            I => \N__10239\
        );

    \I__2434\ : Span4Mux_v
    port map (
            O => \N__10239\,
            I => \N__10235\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10238\,
            I => \N__10232\
        );

    \I__2432\ : Sp12to4
    port map (
            O => \N__10235\,
            I => \N__10226\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__10232\,
            I => \N__10226\
        );

    \I__2430\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10223\
        );

    \I__2429\ : Span12Mux_h
    port map (
            O => \N__10226\,
            I => \N__10220\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__10223\,
            I => \N__10217\
        );

    \I__2427\ : Odrv12
    port map (
            O => \N__10220\,
            I => \CIA_SPACE\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__10217\,
            I => \CIA_SPACE\
        );

    \I__2425\ : IoInMux
    port map (
            O => \N__10212\,
            I => \N__10209\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__10209\,
            I => \N__10206\
        );

    \I__2423\ : Span4Mux_s1_v
    port map (
            O => \N__10206\,
            I => \N__10203\
        );

    \I__2422\ : Sp12to4
    port map (
            O => \N__10203\,
            I => \N__10200\
        );

    \I__2421\ : Span12Mux_h
    port map (
            O => \N__10200\,
            I => \N__10197\
        );

    \I__2420\ : Span12Mux_v
    port map (
            O => \N__10197\,
            I => \N__10194\
        );

    \I__2419\ : Odrv12
    port map (
            O => \N__10194\,
            I => \TCIn_1_i\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10191\,
            I => \N__10188\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__10188\,
            I => \N__10184\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10187\,
            I => \N__10181\
        );

    \I__2415\ : Span4Mux_v
    port map (
            O => \N__10184\,
            I => \N__10171\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__10181\,
            I => \N__10171\
        );

    \I__2413\ : CascadeMux
    port map (
            O => \N__10180\,
            I => \N__10164\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__10179\,
            I => \N__10161\
        );

    \I__2411\ : InMux
    port map (
            O => \N__10178\,
            I => \N__10157\
        );

    \I__2410\ : CascadeMux
    port map (
            O => \N__10177\,
            I => \N__10154\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10176\,
            I => \N__10150\
        );

    \I__2408\ : Span4Mux_v
    port map (
            O => \N__10171\,
            I => \N__10141\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10170\,
            I => \N__10138\
        );

    \I__2406\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10135\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10124\
        );

    \I__2404\ : InMux
    port map (
            O => \N__10167\,
            I => \N__10124\
        );

    \I__2403\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10124\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10124\
        );

    \I__2401\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10124\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__10157\,
            I => \N__10121\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10116\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10153\,
            I => \N__10116\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__10150\,
            I => \N__10113\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10149\,
            I => \N__10110\
        );

    \I__2395\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10107\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10104\
        );

    \I__2393\ : CascadeMux
    port map (
            O => \N__10146\,
            I => \N__10101\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__10145\,
            I => \N__10098\
        );

    \I__2391\ : CascadeMux
    port map (
            O => \N__10144\,
            I => \N__10095\
        );

    \I__2390\ : Span4Mux_h
    port map (
            O => \N__10141\,
            I => \N__10081\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__10138\,
            I => \N__10081\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__10135\,
            I => \N__10081\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10124\,
            I => \N__10081\
        );

    \I__2386\ : Span4Mux_h
    port map (
            O => \N__10121\,
            I => \N__10081\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__10116\,
            I => \N__10081\
        );

    \I__2384\ : Span4Mux_v
    port map (
            O => \N__10113\,
            I => \N__10073\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__10110\,
            I => \N__10073\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__10107\,
            I => \N__10073\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10104\,
            I => \N__10070\
        );

    \I__2380\ : InMux
    port map (
            O => \N__10101\,
            I => \N__10063\
        );

    \I__2379\ : InMux
    port map (
            O => \N__10098\,
            I => \N__10063\
        );

    \I__2378\ : InMux
    port map (
            O => \N__10095\,
            I => \N__10063\
        );

    \I__2377\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10057\
        );

    \I__2376\ : Span4Mux_v
    port map (
            O => \N__10081\,
            I => \N__10054\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10080\,
            I => \N__10051\
        );

    \I__2374\ : Span4Mux_v
    port map (
            O => \N__10073\,
            I => \N__10048\
        );

    \I__2373\ : Span4Mux_h
    port map (
            O => \N__10070\,
            I => \N__10043\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10063\,
            I => \N__10043\
        );

    \I__2371\ : InMux
    port map (
            O => \N__10062\,
            I => \N__10038\
        );

    \I__2370\ : InMux
    port map (
            O => \N__10061\,
            I => \N__10038\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10060\,
            I => \N__10035\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__10057\,
            I => \N__10028\
        );

    \I__2367\ : Span4Mux_h
    port map (
            O => \N__10054\,
            I => \N__10028\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__10051\,
            I => \N__10028\
        );

    \I__2365\ : Span4Mux_h
    port map (
            O => \N__10048\,
            I => \N__10024\
        );

    \I__2364\ : Span4Mux_h
    port map (
            O => \N__10043\,
            I => \N__10017\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10038\,
            I => \N__10017\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10035\,
            I => \N__10017\
        );

    \I__2361\ : Span4Mux_v
    port map (
            O => \N__10028\,
            I => \N__10014\
        );

    \I__2360\ : InMux
    port map (
            O => \N__10027\,
            I => \N__10011\
        );

    \I__2359\ : Span4Mux_h
    port map (
            O => \N__10024\,
            I => \N__10006\
        );

    \I__2358\ : Span4Mux_v
    port map (
            O => \N__10017\,
            I => \N__10006\
        );

    \I__2357\ : Sp12to4
    port map (
            O => \N__10014\,
            I => \N__10002\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10011\,
            I => \N__9999\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__10006\,
            I => \N__9996\
        );

    \I__2354\ : InMux
    port map (
            O => \N__10005\,
            I => \N__9993\
        );

    \I__2353\ : Span12Mux_h
    port map (
            O => \N__10002\,
            I => \N__9990\
        );

    \I__2352\ : Span12Mux_v
    port map (
            O => \N__9999\,
            I => \N__9983\
        );

    \I__2351\ : Sp12to4
    port map (
            O => \N__9996\,
            I => \N__9983\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__9993\,
            I => \N__9983\
        );

    \I__2349\ : Span12Mux_v
    port map (
            O => \N__9990\,
            I => \N__9978\
        );

    \I__2348\ : Span12Mux_h
    port map (
            O => \N__9983\,
            I => \N__9978\
        );

    \I__2347\ : Odrv12
    port map (
            O => \N__9978\,
            I => \RESETn_c\
        );

    \I__2346\ : InMux
    port map (
            O => \N__9975\,
            I => \N__9971\
        );

    \I__2345\ : InMux
    port map (
            O => \N__9974\,
            I => \N__9968\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__9971\,
            I => \N__9965\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__9968\,
            I => \N__9962\
        );

    \I__2342\ : Span12Mux_s11_v
    port map (
            O => \N__9965\,
            I => \N__9958\
        );

    \I__2341\ : Span4Mux_h
    port map (
            O => \N__9962\,
            I => \N__9955\
        );

    \I__2340\ : InMux
    port map (
            O => \N__9961\,
            I => \N__9952\
        );

    \I__2339\ : Odrv12
    port map (
            O => \N__9958\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__9955\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__9952\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__9945\,
            I => \U409_CIA.CIA_CLK_COUNT11_3_cascade_\
        );

    \I__2335\ : InMux
    port map (
            O => \N__9942\,
            I => \N__9939\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__9939\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0\
        );

    \I__2333\ : InMux
    port map (
            O => \N__9936\,
            I => \N__9933\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__9933\,
            I => \U409_CIA.CIA_CLK_COUNT11_3\
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__9930\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__9927\,
            I => \U409_CIA.CLK_CIA6_4_cascade_\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__9924\,
            I => \U409_CIA.VMA_RNOZ0Z_0_cascade_\
        );

    \I__2328\ : InMux
    port map (
            O => \N__9921\,
            I => \N__9911\
        );

    \I__2327\ : InMux
    port map (
            O => \N__9920\,
            I => \N__9911\
        );

    \I__2326\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9904\
        );

    \I__2325\ : InMux
    port map (
            O => \N__9918\,
            I => \N__9904\
        );

    \I__2324\ : InMux
    port map (
            O => \N__9917\,
            I => \N__9904\
        );

    \I__2323\ : InMux
    port map (
            O => \N__9916\,
            I => \N__9901\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__9911\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__9904\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__9901\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2319\ : InMux
    port map (
            O => \N__9894\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__2318\ : CascadeMux
    port map (
            O => \N__9891\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__2317\ : InMux
    port map (
            O => \N__9888\,
            I => \N__9885\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__9885\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__9882\,
            I => \N__9879\
        );

    \I__2314\ : InMux
    port map (
            O => \N__9879\,
            I => \N__9875\
        );

    \I__2313\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9872\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__9875\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__9872\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2310\ : InMux
    port map (
            O => \N__9867\,
            I => \N__9863\
        );

    \I__2309\ : InMux
    port map (
            O => \N__9866\,
            I => \N__9860\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__9863\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__9860\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2306\ : CascadeMux
    port map (
            O => \N__9855\,
            I => \N__9852\
        );

    \I__2305\ : InMux
    port map (
            O => \N__9852\,
            I => \N__9848\
        );

    \I__2304\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9845\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__9848\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__9845\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2301\ : InMux
    port map (
            O => \N__9840\,
            I => \N__9837\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__9837\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__2299\ : InMux
    port map (
            O => \N__9834\,
            I => \N__9830\
        );

    \I__2298\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9827\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__9830\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__9827\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2295\ : InMux
    port map (
            O => \N__9822\,
            I => \N__9819\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__9819\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__2293\ : InMux
    port map (
            O => \N__9816\,
            I => \N__9812\
        );

    \I__2292\ : InMux
    port map (
            O => \N__9815\,
            I => \N__9809\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__9812\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__9809\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__2289\ : InMux
    port map (
            O => \N__9804\,
            I => \N__9801\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__9801\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__2287\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9794\
        );

    \I__2286\ : InMux
    port map (
            O => \N__9797\,
            I => \N__9791\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__9794\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__9791\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__2283\ : InMux
    port map (
            O => \N__9786\,
            I => \N__9773\
        );

    \I__2282\ : InMux
    port map (
            O => \N__9785\,
            I => \N__9773\
        );

    \I__2281\ : InMux
    port map (
            O => \N__9784\,
            I => \N__9768\
        );

    \I__2280\ : InMux
    port map (
            O => \N__9783\,
            I => \N__9768\
        );

    \I__2279\ : InMux
    port map (
            O => \N__9782\,
            I => \N__9759\
        );

    \I__2278\ : InMux
    port map (
            O => \N__9781\,
            I => \N__9759\
        );

    \I__2277\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9759\
        );

    \I__2276\ : InMux
    port map (
            O => \N__9779\,
            I => \N__9759\
        );

    \I__2275\ : InMux
    port map (
            O => \N__9778\,
            I => \N__9756\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__9773\,
            I => \N__9753\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__9768\,
            I => \N__9750\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__9759\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__9756\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2270\ : Odrv4
    port map (
            O => \N__9753\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__9750\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__9741\,
            I => \N__9737\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9727\
        );

    \I__2266\ : InMux
    port map (
            O => \N__9737\,
            I => \N__9724\
        );

    \I__2265\ : InMux
    port map (
            O => \N__9736\,
            I => \N__9719\
        );

    \I__2264\ : InMux
    port map (
            O => \N__9735\,
            I => \N__9719\
        );

    \I__2263\ : InMux
    port map (
            O => \N__9734\,
            I => \N__9716\
        );

    \I__2262\ : InMux
    port map (
            O => \N__9733\,
            I => \N__9707\
        );

    \I__2261\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9707\
        );

    \I__2260\ : InMux
    port map (
            O => \N__9731\,
            I => \N__9707\
        );

    \I__2259\ : InMux
    port map (
            O => \N__9730\,
            I => \N__9707\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__9727\,
            I => \N__9704\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__9724\,
            I => \N__9699\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__9719\,
            I => \N__9699\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__9716\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__9707\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2253\ : Odrv4
    port map (
            O => \N__9704\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__9699\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__9690\,
            I => \N__9687\
        );

    \I__2250\ : InMux
    port map (
            O => \N__9687\,
            I => \N__9677\
        );

    \I__2249\ : InMux
    port map (
            O => \N__9686\,
            I => \N__9674\
        );

    \I__2248\ : InMux
    port map (
            O => \N__9685\,
            I => \N__9669\
        );

    \I__2247\ : InMux
    port map (
            O => \N__9684\,
            I => \N__9669\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__9683\,
            I => \N__9666\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__9682\,
            I => \N__9663\
        );

    \I__2244\ : CascadeMux
    port map (
            O => \N__9681\,
            I => \N__9660\
        );

    \I__2243\ : CascadeMux
    port map (
            O => \N__9680\,
            I => \N__9657\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__9677\,
            I => \N__9652\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__9674\,
            I => \N__9652\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__9669\,
            I => \N__9649\
        );

    \I__2239\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9644\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9663\,
            I => \N__9644\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9639\
        );

    \I__2236\ : InMux
    port map (
            O => \N__9657\,
            I => \N__9639\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__9652\,
            I => \N__9634\
        );

    \I__2234\ : Span4Mux_v
    port map (
            O => \N__9649\,
            I => \N__9634\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__9644\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__9639\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__9634\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2230\ : InMux
    port map (
            O => \N__9627\,
            I => \N__9624\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__9624\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9617\
        );

    \I__2227\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9614\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9617\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__9614\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__2224\ : ClkMux
    port map (
            O => \N__9609\,
            I => \N__9573\
        );

    \I__2223\ : ClkMux
    port map (
            O => \N__9608\,
            I => \N__9573\
        );

    \I__2222\ : ClkMux
    port map (
            O => \N__9607\,
            I => \N__9573\
        );

    \I__2221\ : ClkMux
    port map (
            O => \N__9606\,
            I => \N__9573\
        );

    \I__2220\ : ClkMux
    port map (
            O => \N__9605\,
            I => \N__9573\
        );

    \I__2219\ : ClkMux
    port map (
            O => \N__9604\,
            I => \N__9573\
        );

    \I__2218\ : ClkMux
    port map (
            O => \N__9603\,
            I => \N__9573\
        );

    \I__2217\ : ClkMux
    port map (
            O => \N__9602\,
            I => \N__9573\
        );

    \I__2216\ : ClkMux
    port map (
            O => \N__9601\,
            I => \N__9573\
        );

    \I__2215\ : ClkMux
    port map (
            O => \N__9600\,
            I => \N__9573\
        );

    \I__2214\ : ClkMux
    port map (
            O => \N__9599\,
            I => \N__9573\
        );

    \I__2213\ : ClkMux
    port map (
            O => \N__9598\,
            I => \N__9573\
        );

    \I__2212\ : GlobalMux
    port map (
            O => \N__9573\,
            I => \N__9570\
        );

    \I__2211\ : gio2CtrlBuf
    port map (
            O => \N__9570\,
            I => \CLK6_c_g\
        );

    \I__2210\ : InMux
    port map (
            O => \N__9567\,
            I => \N__9564\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__9564\,
            I => \U409_CIA.CLK_CIA6_3\
        );

    \I__2208\ : InMux
    port map (
            O => \N__9561\,
            I => \N__9557\
        );

    \I__2207\ : InMux
    port map (
            O => \N__9560\,
            I => \N__9554\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__9557\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9554\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9549\,
            I => \N__9546\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__9546\,
            I => \N__9543\
        );

    \I__2202\ : Span4Mux_h
    port map (
            O => \N__9543\,
            I => \N__9540\
        );

    \I__2201\ : Odrv4
    port map (
            O => \N__9540\,
            I => \U409_TICK.TICK503_11\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__9537\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__2199\ : InMux
    port map (
            O => \N__9534\,
            I => \N__9530\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9533\,
            I => \N__9527\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__9530\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__9527\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9519\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__9519\,
            I => \N__9515\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9518\,
            I => \N__9512\
        );

    \I__2192\ : Odrv4
    port map (
            O => \N__9515\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__9512\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2190\ : InMux
    port map (
            O => \N__9507\,
            I => \N__9503\
        );

    \I__2189\ : InMux
    port map (
            O => \N__9506\,
            I => \N__9500\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__9503\,
            I => \N__9497\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__9500\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2186\ : Odrv4
    port map (
            O => \N__9497\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__9492\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9489\,
            I => \N__9486\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__9486\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9479\
        );

    \I__2181\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9476\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__9479\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9476\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__9471\,
            I => \N__9468\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9468\,
            I => \N__9465\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9465\,
            I => \N__9462\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__9462\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__2174\ : IoInMux
    port map (
            O => \N__9459\,
            I => \N__9456\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__9456\,
            I => \N__9453\
        );

    \I__2172\ : Span4Mux_s2_v
    port map (
            O => \N__9453\,
            I => \N__9450\
        );

    \I__2171\ : Span4Mux_v
    port map (
            O => \N__9450\,
            I => \N__9447\
        );

    \I__2170\ : Sp12to4
    port map (
            O => \N__9447\,
            I => \N__9444\
        );

    \I__2169\ : Span12Mux_h
    port map (
            O => \N__9444\,
            I => \N__9440\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9443\,
            I => \N__9437\
        );

    \I__2167\ : Odrv12
    port map (
            O => \N__9440\,
            I => \TICK50_c\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__9437\,
            I => \TICK50_c\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__9432\,
            I => \N__9429\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9429\,
            I => \N__9426\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__9426\,
            I => \N__9423\
        );

    \I__2162\ : Span4Mux_h
    port map (
            O => \N__9423\,
            I => \N__9420\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__9420\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__9417\,
            I => \N__9413\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9410\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9407\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9410\,
            I => \N__9404\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__9407\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__9404\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9390\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9383\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9383\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9383\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9395\,
            I => \N__9376\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9394\,
            I => \N__9376\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9376\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__9390\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__9383\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__9376\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9369\,
            I => \N__9359\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9368\,
            I => \N__9352\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9367\,
            I => \N__9352\
        );

    \I__2141\ : InMux
    port map (
            O => \N__9366\,
            I => \N__9352\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9365\,
            I => \N__9343\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9343\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9343\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9343\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9359\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__9352\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9343\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__9336\,
            I => \N__9330\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__9335\,
            I => \N__9326\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__9334\,
            I => \N__9322\
        );

    \I__2130\ : CascadeMux
    port map (
            O => \N__9333\,
            I => \N__9319\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9330\,
            I => \N__9315\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9310\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9326\,
            I => \N__9310\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9301\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9322\,
            I => \N__9301\
        );

    \I__2124\ : InMux
    port map (
            O => \N__9319\,
            I => \N__9301\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9301\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9315\,
            I => \N__9298\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__9310\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9301\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__9298\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2118\ : IoInMux
    port map (
            O => \N__9291\,
            I => \N__9288\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9288\,
            I => \N__9285\
        );

    \I__2116\ : Span4Mux_s3_v
    port map (
            O => \N__9285\,
            I => \N__9282\
        );

    \I__2115\ : Span4Mux_v
    port map (
            O => \N__9282\,
            I => \N__9279\
        );

    \I__2114\ : Span4Mux_v
    port map (
            O => \N__9279\,
            I => \N__9276\
        );

    \I__2113\ : Span4Mux_h
    port map (
            O => \N__9276\,
            I => \N__9272\
        );

    \I__2112\ : InMux
    port map (
            O => \N__9275\,
            I => \N__9269\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__9272\,
            I => \TICK60_c\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9269\,
            I => \TICK60_c\
        );

    \I__2109\ : InMux
    port map (
            O => \N__9264\,
            I => \N__9260\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9257\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__9260\,
            I => \N__9254\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__9257\,
            I => \N__9251\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__9254\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__9251\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2103\ : InMux
    port map (
            O => \N__9246\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9243\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9240\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9237\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9234\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9231\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__2097\ : InMux
    port map (
            O => \N__9228\,
            I => \N__9224\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9227\,
            I => \N__9221\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__9224\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__9221\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__9216\,
            I => \U409_CIA.CLK_CIA_r_1_0_cascade_\
        );

    \I__2092\ : IoInMux
    port map (
            O => \N__9213\,
            I => \N__9210\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__9210\,
            I => \N__9207\
        );

    \I__2090\ : IoSpan4Mux
    port map (
            O => \N__9207\,
            I => \N__9204\
        );

    \I__2089\ : Span4Mux_s3_v
    port map (
            O => \N__9204\,
            I => \N__9201\
        );

    \I__2088\ : Sp12to4
    port map (
            O => \N__9201\,
            I => \N__9196\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9200\,
            I => \N__9193\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__9199\,
            I => \N__9189\
        );

    \I__2085\ : Span12Mux_s10_v
    port map (
            O => \N__9196\,
            I => \N__9186\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__9193\,
            I => \N__9183\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9180\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9189\,
            I => \N__9177\
        );

    \I__2081\ : Odrv12
    port map (
            O => \N__9186\,
            I => \CLK_CIA_c\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__9183\,
            I => \CLK_CIA_c\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9180\,
            I => \CLK_CIA_c\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__9177\,
            I => \CLK_CIA_c\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9168\,
            I => \N__9165\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9165\,
            I => \N__9161\
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__9164\,
            I => \N__9158\
        );

    \I__2074\ : Span4Mux_h
    port map (
            O => \N__9161\,
            I => \N__9155\
        );

    \I__2073\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9152\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__9155\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__9152\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__9147\,
            I => \N__9144\
        );

    \I__2069\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9141\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9141\,
            I => \N__9137\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9140\,
            I => \N__9134\
        );

    \I__2066\ : Odrv12
    port map (
            O => \N__9137\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9134\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2064\ : InMux
    port map (
            O => \N__9129\,
            I => \N__9125\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__9128\,
            I => \N__9121\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9125\,
            I => \N__9117\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__9124\,
            I => \N__9114\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9121\,
            I => \N__9111\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9120\,
            I => \N__9108\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__9117\,
            I => \N__9105\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9114\,
            I => \N__9102\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__9111\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__9108\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__9105\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9102\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__9093\,
            I => \N__9090\
        );

    \I__2051\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9086\
        );

    \I__2050\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9083\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9086\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9083\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9078\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9075\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9072\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9069\,
            I => \N__9066\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__9066\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9063\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9060\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9057\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9054\,
            I => \N__9050\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9053\,
            I => \N__9047\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__9050\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9047\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9042\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9039\,
            I => \bfn_14_6_0_\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9036\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9033\,
            I => \N__9030\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9030\,
            I => \N__9020\
        );

    \I__2030\ : SRMux
    port map (
            O => \N__9029\,
            I => \N__8991\
        );

    \I__2029\ : SRMux
    port map (
            O => \N__9028\,
            I => \N__8991\
        );

    \I__2028\ : SRMux
    port map (
            O => \N__9027\,
            I => \N__8991\
        );

    \I__2027\ : SRMux
    port map (
            O => \N__9026\,
            I => \N__8991\
        );

    \I__2026\ : SRMux
    port map (
            O => \N__9025\,
            I => \N__8991\
        );

    \I__2025\ : SRMux
    port map (
            O => \N__9024\,
            I => \N__8991\
        );

    \I__2024\ : SRMux
    port map (
            O => \N__9023\,
            I => \N__8991\
        );

    \I__2023\ : Glb2LocalMux
    port map (
            O => \N__9020\,
            I => \N__8991\
        );

    \I__2022\ : SRMux
    port map (
            O => \N__9019\,
            I => \N__8991\
        );

    \I__2021\ : SRMux
    port map (
            O => \N__9018\,
            I => \N__8991\
        );

    \I__2020\ : SRMux
    port map (
            O => \N__9017\,
            I => \N__8991\
        );

    \I__2019\ : SRMux
    port map (
            O => \N__9016\,
            I => \N__8991\
        );

    \I__2018\ : GlobalMux
    port map (
            O => \N__8991\,
            I => \N__8988\
        );

    \I__2017\ : gio2CtrlBuf
    port map (
            O => \N__8988\,
            I => \RESETn_c_i_g\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__8985\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_\
        );

    \I__2015\ : InMux
    port map (
            O => \N__8982\,
            I => \N__8978\
        );

    \I__2014\ : InMux
    port map (
            O => \N__8981\,
            I => \N__8975\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__8978\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__8975\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__8970\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out_cascade_\
        );

    \I__2010\ : InMux
    port map (
            O => \N__8967\,
            I => \N__8959\
        );

    \I__2009\ : InMux
    port map (
            O => \N__8966\,
            I => \N__8959\
        );

    \I__2008\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8954\
        );

    \I__2007\ : InMux
    port map (
            O => \N__8964\,
            I => \N__8954\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__8959\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__8954\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__2004\ : InMux
    port map (
            O => \N__8949\,
            I => \N__8938\
        );

    \I__2003\ : InMux
    port map (
            O => \N__8948\,
            I => \N__8938\
        );

    \I__2002\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8938\
        );

    \I__2001\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8933\
        );

    \I__2000\ : InMux
    port map (
            O => \N__8945\,
            I => \N__8933\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__8938\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__8933\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1997\ : InMux
    port map (
            O => \N__8928\,
            I => \N__8919\
        );

    \I__1996\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8919\
        );

    \I__1995\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8914\
        );

    \I__1994\ : InMux
    port map (
            O => \N__8925\,
            I => \N__8914\
        );

    \I__1993\ : InMux
    port map (
            O => \N__8924\,
            I => \N__8911\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__8919\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__8914\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__8911\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1989\ : CascadeMux
    port map (
            O => \N__8904\,
            I => \N__8900\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__8903\,
            I => \N__8895\
        );

    \I__1987\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8885\
        );

    \I__1986\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8885\
        );

    \I__1985\ : InMux
    port map (
            O => \N__8898\,
            I => \N__8885\
        );

    \I__1984\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8880\
        );

    \I__1983\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8880\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8875\
        );

    \I__1981\ : InMux
    port map (
            O => \N__8892\,
            I => \N__8875\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__8885\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__8880\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__8875\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1977\ : InMux
    port map (
            O => \N__8868\,
            I => \N__8862\
        );

    \I__1976\ : InMux
    port map (
            O => \N__8867\,
            I => \N__8857\
        );

    \I__1975\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8857\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8865\,
            I => \N__8854\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__8862\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__8857\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__8854\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__8847\,
            I => \N__8843\
        );

    \I__1969\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8838\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8838\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__8838\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__1966\ : InMux
    port map (
            O => \N__8835\,
            I => \N__8826\
        );

    \I__1965\ : InMux
    port map (
            O => \N__8834\,
            I => \N__8826\
        );

    \I__1964\ : InMux
    port map (
            O => \N__8833\,
            I => \N__8823\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8818\
        );

    \I__1962\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8818\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8826\,
            I => \N__8815\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8823\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__8818\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__8815\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__8808\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__8805\,
            I => \N__8799\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8804\,
            I => \N__8788\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8803\,
            I => \N__8788\
        );

    \I__1953\ : InMux
    port map (
            O => \N__8802\,
            I => \N__8788\
        );

    \I__1952\ : InMux
    port map (
            O => \N__8799\,
            I => \N__8788\
        );

    \I__1951\ : InMux
    port map (
            O => \N__8798\,
            I => \N__8783\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8797\,
            I => \N__8783\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__8788\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__8783\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1947\ : SRMux
    port map (
            O => \N__8778\,
            I => \N__8774\
        );

    \I__1946\ : SRMux
    port map (
            O => \N__8777\,
            I => \N__8770\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__8774\,
            I => \N__8767\
        );

    \I__1944\ : SRMux
    port map (
            O => \N__8773\,
            I => \N__8763\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__8770\,
            I => \N__8760\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__8767\,
            I => \N__8757\
        );

    \I__1941\ : SRMux
    port map (
            O => \N__8766\,
            I => \N__8754\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__8763\,
            I => \N__8751\
        );

    \I__1939\ : Span4Mux_v
    port map (
            O => \N__8760\,
            I => \N__8748\
        );

    \I__1938\ : Span4Mux_v
    port map (
            O => \N__8757\,
            I => \N__8743\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__8754\,
            I => \N__8743\
        );

    \I__1936\ : Span4Mux_v
    port map (
            O => \N__8751\,
            I => \N__8740\
        );

    \I__1935\ : Sp12to4
    port map (
            O => \N__8748\,
            I => \N__8735\
        );

    \I__1934\ : Sp12to4
    port map (
            O => \N__8743\,
            I => \N__8735\
        );

    \I__1933\ : Odrv4
    port map (
            O => \N__8740\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1932\ : Odrv12
    port map (
            O => \N__8735\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8730\,
            I => \N__8725\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8729\,
            I => \N__8722\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8728\,
            I => \N__8719\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__8725\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__8722\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__8719\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8712\,
            I => \N__8709\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8709\,
            I => \N__8705\
        );

    \I__1923\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8702\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__8705\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__8702\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8693\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8696\,
            I => \N__8690\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8693\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__8690\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__8685\,
            I => \N__8682\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8682\,
            I => \N__8678\
        );

    \I__1914\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8675\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8678\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__8675\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1911\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8666\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8663\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__8666\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8663\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__1907\ : InMux
    port map (
            O => \N__8658\,
            I => \N__8655\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__8655\,
            I => \N__8651\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8648\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__8651\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__8648\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8643\,
            I => \N__8639\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8636\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__8639\,
            I => \N__8633\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__8636\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__8633\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8628\,
            I => \N__8625\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__8625\,
            I => \U409_TICK.TICK603_11\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8622\,
            I => \N__8618\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8615\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__8618\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__8615\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__1891\ : CascadeMux
    port map (
            O => \N__8610\,
            I => \U409_TICK.TICK603_8_cascade_\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8607\,
            I => \N__8604\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8604\,
            I => \N__8600\
        );

    \I__1888\ : InMux
    port map (
            O => \N__8603\,
            I => \N__8597\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__8600\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__8597\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__8592\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__8589\,
            I => \N__8586\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8586\,
            I => \N__8580\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8577\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8584\,
            I => \N__8572\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8572\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__8580\,
            I => \N__8569\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8577\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8572\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__8569\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__1875\ : CascadeMux
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8559\,
            I => \N__8553\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8553\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8553\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8541\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8541\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8541\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8541\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__1867\ : InMux
    port map (
            O => \N__8538\,
            I => \N__8532\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8537\,
            I => \N__8525\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8536\,
            I => \N__8525\
        );

    \I__1864\ : InMux
    port map (
            O => \N__8535\,
            I => \N__8525\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8532\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8525\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1861\ : InMux
    port map (
            O => \N__8520\,
            I => \N__8515\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8510\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8518\,
            I => \N__8510\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8515\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__8510\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8505\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8502\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__1854\ : InMux
    port map (
            O => \N__8499\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8496\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8493\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__1851\ : InMux
    port map (
            O => \N__8490\,
            I => \N__8487\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8487\,
            I => \N__8484\
        );

    \I__1849\ : Odrv12
    port map (
            O => \N__8484\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__8481\,
            I => \N__8478\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8478\,
            I => \N__8475\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__8475\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8472\,
            I => \N__8469\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8469\,
            I => \N__8466\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__8466\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__1842\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8459\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8456\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8459\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8456\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8451\,
            I => \N__8448\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8448\,
            I => \N__8444\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8441\
        );

    \I__1835\ : Odrv4
    port map (
            O => \N__8444\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__8441\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__8436\,
            I => \N__8432\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8429\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8426\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8429\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__8426\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8416\
        );

    \I__1827\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8413\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8419\,
            I => \N__8410\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__8416\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8413\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8410\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8403\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8400\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8397\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8394\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8391\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8388\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8385\,
            I => \N__8382\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8382\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8379\,
            I => \bfn_13_7_0_\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8376\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8373\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8364\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8369\,
            I => \N__8361\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8368\,
            I => \N__8358\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8367\,
            I => \N__8355\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8364\,
            I => \N__8350\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8361\,
            I => \N__8350\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__8358\,
            I => \N__8345\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8355\,
            I => \N__8340\
        );

    \I__1803\ : Span4Mux_v
    port map (
            O => \N__8350\,
            I => \N__8340\
        );

    \I__1802\ : InMux
    port map (
            O => \N__8349\,
            I => \N__8337\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8334\
        );

    \I__1800\ : Span4Mux_v
    port map (
            O => \N__8345\,
            I => \N__8331\
        );

    \I__1799\ : Span4Mux_h
    port map (
            O => \N__8340\,
            I => \N__8326\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8337\,
            I => \N__8326\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8334\,
            I => \N__8321\
        );

    \I__1796\ : Sp12to4
    port map (
            O => \N__8331\,
            I => \N__8321\
        );

    \I__1795\ : Span4Mux_h
    port map (
            O => \N__8326\,
            I => \N__8318\
        );

    \I__1794\ : Span12Mux_h
    port map (
            O => \N__8321\,
            I => \N__8313\
        );

    \I__1793\ : Sp12to4
    port map (
            O => \N__8318\,
            I => \N__8313\
        );

    \I__1792\ : Span12Mux_v
    port map (
            O => \N__8313\,
            I => \N__8310\
        );

    \I__1791\ : Odrv12
    port map (
            O => \N__8310\,
            I => \TSn_c\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__8307\,
            I => \N__8298\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__8306\,
            I => \N__8295\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8305\,
            I => \N__8292\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8304\,
            I => \N__8289\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8286\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8283\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8280\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8298\,
            I => \N__8277\
        );

    \I__1782\ : InMux
    port map (
            O => \N__8295\,
            I => \N__8274\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__8292\,
            I => \N__8271\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8289\,
            I => \N__8259\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8286\,
            I => \N__8256\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__8283\,
            I => \N__8253\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__8280\,
            I => \N__8250\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8277\,
            I => \N__8247\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8274\,
            I => \N__8244\
        );

    \I__1774\ : Glb2LocalMux
    port map (
            O => \N__8271\,
            I => \N__8211\
        );

    \I__1773\ : ClkMux
    port map (
            O => \N__8270\,
            I => \N__8211\
        );

    \I__1772\ : ClkMux
    port map (
            O => \N__8269\,
            I => \N__8211\
        );

    \I__1771\ : ClkMux
    port map (
            O => \N__8268\,
            I => \N__8211\
        );

    \I__1770\ : ClkMux
    port map (
            O => \N__8267\,
            I => \N__8211\
        );

    \I__1769\ : ClkMux
    port map (
            O => \N__8266\,
            I => \N__8211\
        );

    \I__1768\ : ClkMux
    port map (
            O => \N__8265\,
            I => \N__8211\
        );

    \I__1767\ : ClkMux
    port map (
            O => \N__8264\,
            I => \N__8211\
        );

    \I__1766\ : ClkMux
    port map (
            O => \N__8263\,
            I => \N__8211\
        );

    \I__1765\ : ClkMux
    port map (
            O => \N__8262\,
            I => \N__8211\
        );

    \I__1764\ : Glb2LocalMux
    port map (
            O => \N__8259\,
            I => \N__8211\
        );

    \I__1763\ : Glb2LocalMux
    port map (
            O => \N__8256\,
            I => \N__8211\
        );

    \I__1762\ : Glb2LocalMux
    port map (
            O => \N__8253\,
            I => \N__8211\
        );

    \I__1761\ : Glb2LocalMux
    port map (
            O => \N__8250\,
            I => \N__8211\
        );

    \I__1760\ : Glb2LocalMux
    port map (
            O => \N__8247\,
            I => \N__8211\
        );

    \I__1759\ : Glb2LocalMux
    port map (
            O => \N__8244\,
            I => \N__8211\
        );

    \I__1758\ : GlobalMux
    port map (
            O => \N__8211\,
            I => \N__8208\
        );

    \I__1757\ : gio2CtrlBuf
    port map (
            O => \N__8208\,
            I => \CLK40_IN_c_g\
        );

    \I__1756\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8201\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8204\,
            I => \N__8198\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8201\,
            I => \U409_TRANSFER_ACK.N_87\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__8198\,
            I => \U409_TRANSFER_ACK.N_87\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__8193\,
            I => \N__8187\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__8192\,
            I => \N__8184\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8181\
        );

    \I__1749\ : InMux
    port map (
            O => \N__8190\,
            I => \N__8174\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8187\,
            I => \N__8174\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8184\,
            I => \N__8174\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__8181\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8174\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1744\ : IoInMux
    port map (
            O => \N__8169\,
            I => \N__8166\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8166\,
            I => \N__8163\
        );

    \I__1742\ : Span12Mux_s1_v
    port map (
            O => \N__8163\,
            I => \N__8160\
        );

    \I__1741\ : Odrv12
    port map (
            O => \N__8160\,
            I => \RESETn_c_i\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8157\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__1739\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8150\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8147\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__8150\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__8147\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__8142\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3_cascade_\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__8139\,
            I => \N__8136\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8136\,
            I => \N__8130\
        );

    \I__1732\ : InMux
    port map (
            O => \N__8135\,
            I => \N__8130\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__8130\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8127\,
            I => \N__8124\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__8124\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a3_3\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__8121\,
            I => \U409_TRANSFER_ACK.N_87_cascade_\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8114\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8117\,
            I => \N__8111\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8114\,
            I => \U409_TRANSFER_ACK.N_77\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8111\,
            I => \U409_TRANSFER_ACK.N_77\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__8106\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8094\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8102\,
            I => \N__8094\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8101\,
            I => \N__8094\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8094\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__8091\,
            I => \U409_TRANSFER_ACK.N_17_mux_cascade_\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__8088\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__8085\,
            I => \U409_TRANSFER_ACK.N_6_0_cascade_\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8082\,
            I => \N__8079\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8079\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8076\,
            I => \N__8070\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8075\,
            I => \N__8070\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8070\,
            I => \U409_TRANSFER_ACK.N_3_0\
        );

    \I__1710\ : CascadeMux
    port map (
            O => \N__8067\,
            I => \N__8061\
        );

    \I__1709\ : CascadeMux
    port map (
            O => \N__8066\,
            I => \N__8058\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8054\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8045\
        );

    \I__1706\ : InMux
    port map (
            O => \N__8061\,
            I => \N__8045\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8058\,
            I => \N__8045\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8057\,
            I => \N__8045\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__8054\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8045\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8040\,
            I => \N__8037\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8037\,
            I => \U409_TRANSFER_ACK.N_17_mux\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__8034\,
            I => \N__8029\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8033\,
            I => \N__8024\
        );

    \I__1697\ : InMux
    port map (
            O => \N__8032\,
            I => \N__8024\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8029\,
            I => \N__8021\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8024\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__8021\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8016\,
            I => \N__8012\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8015\,
            I => \N__8009\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__8012\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__8009\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8004\,
            I => \N__7998\
        );

    \I__1688\ : InMux
    port map (
            O => \N__8003\,
            I => \N__7991\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8002\,
            I => \N__7991\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8001\,
            I => \N__7991\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__7998\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__7991\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__7986\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\
        );

    \I__1682\ : IoInMux
    port map (
            O => \N__7983\,
            I => \N__7979\
        );

    \I__1681\ : IoInMux
    port map (
            O => \N__7982\,
            I => \N__7976\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__7979\,
            I => \N__7970\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__7976\,
            I => \N__7970\
        );

    \I__1678\ : IoInMux
    port map (
            O => \N__7975\,
            I => \N__7967\
        );

    \I__1677\ : IoSpan4Mux
    port map (
            O => \N__7970\,
            I => \N__7964\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__7967\,
            I => \N__7961\
        );

    \I__1675\ : Span4Mux_s3_v
    port map (
            O => \N__7964\,
            I => \N__7958\
        );

    \I__1674\ : Span4Mux_s3_v
    port map (
            O => \N__7961\,
            I => \N__7955\
        );

    \I__1673\ : Sp12to4
    port map (
            O => \N__7958\,
            I => \N__7950\
        );

    \I__1672\ : Sp12to4
    port map (
            O => \N__7955\,
            I => \N__7950\
        );

    \I__1671\ : Span12Mux_s9_h
    port map (
            O => \N__7950\,
            I => \N__7947\
        );

    \I__1670\ : Span12Mux_v
    port map (
            O => \N__7947\,
            I => \N__7942\
        );

    \I__1669\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7937\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7945\,
            I => \N__7937\
        );

    \I__1667\ : Odrv12
    port map (
            O => \N__7942\,
            I => \TACK_OUTn\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__7937\,
            I => \TACK_OUTn\
        );

    \I__1665\ : InMux
    port map (
            O => \N__7932\,
            I => \N__7929\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__7929\,
            I => \U409_TRANSFER_ACK.TACK_OUTn_3_0\
        );

    \I__1663\ : InMux
    port map (
            O => \N__7926\,
            I => \N__7922\
        );

    \I__1662\ : InMux
    port map (
            O => \N__7925\,
            I => \N__7918\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__7922\,
            I => \N__7915\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__7921\,
            I => \N__7910\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__7918\,
            I => \N__7904\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__7915\,
            I => \N__7904\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7914\,
            I => \N__7901\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7913\,
            I => \N__7894\
        );

    \I__1655\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7894\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7894\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__7904\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__7901\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__7894\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__7887\,
            I => \N__7884\
        );

    \I__1649\ : InMux
    port map (
            O => \N__7884\,
            I => \N__7881\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__7881\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_2\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7873\
        );

    \I__1646\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7870\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__7876\,
            I => \N__7866\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7873\,
            I => \N__7862\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7870\,
            I => \N__7859\
        );

    \I__1642\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7856\
        );

    \I__1641\ : InMux
    port map (
            O => \N__7866\,
            I => \N__7851\
        );

    \I__1640\ : InMux
    port map (
            O => \N__7865\,
            I => \N__7851\
        );

    \I__1639\ : Odrv4
    port map (
            O => \N__7862\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__7859\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__7856\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__7851\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1635\ : InMux
    port map (
            O => \N__7842\,
            I => \N__7838\
        );

    \I__1634\ : InMux
    port map (
            O => \N__7841\,
            I => \N__7835\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7838\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__7835\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7830\,
            I => \N__7826\
        );

    \I__1630\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7823\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__7826\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__7823\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__7818\,
            I => \N__7814\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__7817\,
            I => \N__7811\
        );

    \I__1625\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7808\
        );

    \I__1624\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7805\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7808\,
            I => \N__7800\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__7805\,
            I => \N__7800\
        );

    \I__1621\ : Span4Mux_h
    port map (
            O => \N__7800\,
            I => \N__7797\
        );

    \I__1620\ : Odrv4
    port map (
            O => \N__7797\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\
        );

    \I__1619\ : InMux
    port map (
            O => \N__7794\,
            I => \N__7790\
        );

    \I__1618\ : InMux
    port map (
            O => \N__7793\,
            I => \N__7787\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__7790\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__7787\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1615\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7779\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7779\,
            I => \N__7776\
        );

    \I__1613\ : Sp12to4
    port map (
            O => \N__7776\,
            I => \N__7773\
        );

    \I__1612\ : Span12Mux_h
    port map (
            O => \N__7773\,
            I => \N__7770\
        );

    \I__1611\ : Span12Mux_v
    port map (
            O => \N__7770\,
            I => \N__7767\
        );

    \I__1610\ : Odrv12
    port map (
            O => \N__7767\,
            I => \TACKn_in\
        );

    \I__1609\ : InMux
    port map (
            O => \N__7764\,
            I => \N__7761\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__7761\,
            I => \N__7757\
        );

    \I__1607\ : InMux
    port map (
            O => \N__7760\,
            I => \N__7754\
        );

    \I__1606\ : Span4Mux_v
    port map (
            O => \N__7757\,
            I => \N__7750\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__7754\,
            I => \N__7747\
        );

    \I__1604\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7744\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__7750\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0\
        );

    \I__1602\ : Odrv4
    port map (
            O => \N__7747\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__7744\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0\
        );

    \I__1600\ : CascadeMux
    port map (
            O => \N__7737\,
            I => \N__7733\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__7736\,
            I => \N__7730\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7725\
        );

    \I__1597\ : InMux
    port map (
            O => \N__7730\,
            I => \N__7725\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__7725\,
            I => \N__7721\
        );

    \I__1595\ : InMux
    port map (
            O => \N__7724\,
            I => \N__7718\
        );

    \I__1594\ : Odrv12
    port map (
            O => \N__7721\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__7718\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__1592\ : InMux
    port map (
            O => \N__7713\,
            I => \N__7707\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7712\,
            I => \N__7707\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__7707\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn\
        );

    \I__1589\ : IoInMux
    port map (
            O => \N__7704\,
            I => \N__7701\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__7701\,
            I => \N__7698\
        );

    \I__1587\ : Span12Mux_s1_v
    port map (
            O => \N__7698\,
            I => \N__7695\
        );

    \I__1586\ : Span12Mux_v
    port map (
            O => \N__7695\,
            I => \N__7692\
        );

    \I__1585\ : Odrv12
    port map (
            O => \N__7692\,
            I => \BUFENn_c\
        );

    \I__1584\ : InMux
    port map (
            O => \N__7689\,
            I => \N__7686\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__7686\,
            I => \N__7683\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__7683\,
            I => \U409_TRANSFER_ACK.N_119\
        );

    \I__1581\ : IoInMux
    port map (
            O => \N__7680\,
            I => \N__7677\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__7677\,
            I => \N__7674\
        );

    \I__1579\ : Span4Mux_s3_v
    port map (
            O => \N__7674\,
            I => \N__7671\
        );

    \I__1578\ : Span4Mux_h
    port map (
            O => \N__7671\,
            I => \N__7668\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__7668\,
            I => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\
        );

    \I__1576\ : IoInMux
    port map (
            O => \N__7665\,
            I => \N__7661\
        );

    \I__1575\ : IoInMux
    port map (
            O => \N__7664\,
            I => \N__7658\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__7661\,
            I => \N__7655\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7658\,
            I => \N__7652\
        );

    \I__1572\ : Span4Mux_s0_v
    port map (
            O => \N__7655\,
            I => \N__7649\
        );

    \I__1571\ : IoSpan4Mux
    port map (
            O => \N__7652\,
            I => \N__7646\
        );

    \I__1570\ : Span4Mux_v
    port map (
            O => \N__7649\,
            I => \N__7643\
        );

    \I__1569\ : Span4Mux_s3_h
    port map (
            O => \N__7646\,
            I => \N__7640\
        );

    \I__1568\ : Span4Mux_v
    port map (
            O => \N__7643\,
            I => \N__7637\
        );

    \I__1567\ : Sp12to4
    port map (
            O => \N__7640\,
            I => \N__7634\
        );

    \I__1566\ : Span4Mux_v
    port map (
            O => \N__7637\,
            I => \N__7631\
        );

    \I__1565\ : Odrv12
    port map (
            O => \N__7634\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__7631\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7626\,
            I => \N__7619\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7625\,
            I => \N__7616\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7624\,
            I => \N__7609\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7623\,
            I => \N__7609\
        );

    \I__1559\ : InMux
    port map (
            O => \N__7622\,
            I => \N__7609\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7619\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7616\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7609\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1555\ : InMux
    port map (
            O => \N__7602\,
            I => \N__7593\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7601\,
            I => \N__7593\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7600\,
            I => \N__7590\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7599\,
            I => \N__7585\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7598\,
            I => \N__7585\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7593\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7590\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7585\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1547\ : IoInMux
    port map (
            O => \N__7578\,
            I => \N__7575\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__7575\,
            I => \N__7572\
        );

    \I__1545\ : Span4Mux_s3_v
    port map (
            O => \N__7572\,
            I => \N__7569\
        );

    \I__1544\ : Sp12to4
    port map (
            O => \N__7569\,
            I => \N__7566\
        );

    \I__1543\ : Span12Mux_h
    port map (
            O => \N__7566\,
            I => \N__7563\
        );

    \I__1542\ : Odrv12
    port map (
            O => \N__7563\,
            I => \ROMENn_c\
        );

    \I__1541\ : CEMux
    port map (
            O => \N__7560\,
            I => \N__7557\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7557\,
            I => \N__7554\
        );

    \I__1539\ : Span4Mux_h
    port map (
            O => \N__7554\,
            I => \N__7551\
        );

    \I__1538\ : Odrv4
    port map (
            O => \N__7551\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_0\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7548\,
            I => \N__7545\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7545\,
            I => \N__7541\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7544\,
            I => \N__7538\
        );

    \I__1534\ : Span4Mux_h
    port map (
            O => \N__7541\,
            I => \N__7535\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7538\,
            I => \AC_TACK\
        );

    \I__1532\ : Odrv4
    port map (
            O => \N__7535\,
            I => \AC_TACK\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__7530\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\
        );

    \I__1530\ : InMux
    port map (
            O => \N__7527\,
            I => \N__7523\
        );

    \I__1529\ : InMux
    port map (
            O => \N__7526\,
            I => \N__7520\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7523\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7520\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7515\,
            I => \N__7509\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7514\,
            I => \N__7502\
        );

    \I__1524\ : InMux
    port map (
            O => \N__7513\,
            I => \N__7502\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7502\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7509\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7502\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__7497\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_cascade_\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__7494\,
            I => \N__7491\
        );

    \I__1518\ : InMux
    port map (
            O => \N__7491\,
            I => \N__7488\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__7488\,
            I => \N__7485\
        );

    \I__1516\ : Span4Mux_v
    port map (
            O => \N__7485\,
            I => \N__7481\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7484\,
            I => \N__7478\
        );

    \I__1514\ : Span4Mux_h
    port map (
            O => \N__7481\,
            I => \N__7475\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7478\,
            I => \N__7472\
        );

    \I__1512\ : Sp12to4
    port map (
            O => \N__7475\,
            I => \N__7467\
        );

    \I__1511\ : Span12Mux_h
    port map (
            O => \N__7472\,
            I => \N__7467\
        );

    \I__1510\ : Span12Mux_v
    port map (
            O => \N__7467\,
            I => \N__7464\
        );

    \I__1509\ : Odrv12
    port map (
            O => \N__7464\,
            I => \D_in_4\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7461\,
            I => \N__7457\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7460\,
            I => \N__7454\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7457\,
            I => \ATA_BASE_4\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7454\,
            I => \ATA_BASE_4\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__7449\,
            I => \N__7446\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7446\,
            I => \N__7443\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7443\,
            I => \N__7440\
        );

    \I__1501\ : Span4Mux_v
    port map (
            O => \N__7440\,
            I => \N__7436\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7439\,
            I => \N__7433\
        );

    \I__1499\ : Span4Mux_v
    port map (
            O => \N__7436\,
            I => \N__7429\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7433\,
            I => \N__7426\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__7432\,
            I => \N__7423\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__7429\,
            I => \N__7420\
        );

    \I__1495\ : Span4Mux_h
    port map (
            O => \N__7426\,
            I => \N__7417\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7423\,
            I => \N__7414\
        );

    \I__1493\ : Sp12to4
    port map (
            O => \N__7420\,
            I => \N__7411\
        );

    \I__1492\ : Sp12to4
    port map (
            O => \N__7417\,
            I => \N__7406\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7414\,
            I => \N__7406\
        );

    \I__1490\ : Span12Mux_h
    port map (
            O => \N__7411\,
            I => \N__7401\
        );

    \I__1489\ : Span12Mux_v
    port map (
            O => \N__7406\,
            I => \N__7401\
        );

    \I__1488\ : Odrv12
    port map (
            O => \N__7401\,
            I => \D_in_5\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7398\,
            I => \N__7394\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7397\,
            I => \N__7391\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7394\,
            I => \ATA_BASE_5\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7391\,
            I => \ATA_BASE_5\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7380\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7373\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7384\,
            I => \N__7373\
        );

    \I__1480\ : InMux
    port map (
            O => \N__7383\,
            I => \N__7373\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7380\,
            I => \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_1\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7373\,
            I => \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_1\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7368\,
            I => \N__7364\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7361\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__7364\,
            I => \ATA_BASE_6\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7361\,
            I => \ATA_BASE_6\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__7356\,
            I => \N__7348\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7355\,
            I => \N__7339\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7354\,
            I => \N__7339\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7353\,
            I => \N__7339\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7352\,
            I => \N__7327\
        );

    \I__1468\ : InMux
    port map (
            O => \N__7351\,
            I => \N__7327\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7348\,
            I => \N__7327\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7347\,
            I => \N__7327\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7346\,
            I => \N__7327\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7339\,
            I => \N__7322\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7338\,
            I => \N__7319\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7327\,
            I => \N__7316\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7326\,
            I => \N__7311\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7311\
        );

    \I__1459\ : Span4Mux_h
    port map (
            O => \N__7322\,
            I => \N__7308\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7319\,
            I => \N__7305\
        );

    \I__1457\ : Span4Mux_h
    port map (
            O => \N__7316\,
            I => \N__7300\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7311\,
            I => \N__7300\
        );

    \I__1455\ : Odrv4
    port map (
            O => \N__7308\,
            I => \un1_AUTOCONFIG_SPACE\
        );

    \I__1454\ : Odrv4
    port map (
            O => \N__7305\,
            I => \un1_AUTOCONFIG_SPACE\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__7300\,
            I => \un1_AUTOCONFIG_SPACE\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7288\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7283\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7291\,
            I => \N__7283\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7288\,
            I => \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_0\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7283\,
            I => \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_0\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__7278\,
            I => \N__7274\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__7277\,
            I => \N__7271\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7274\,
            I => \N__7268\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7265\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7268\,
            I => \N__7259\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__7265\,
            I => \N__7259\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7264\,
            I => \N__7256\
        );

    \I__1440\ : Span4Mux_v
    port map (
            O => \N__7259\,
            I => \N__7253\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__7256\,
            I => \N__7250\
        );

    \I__1438\ : Sp12to4
    port map (
            O => \N__7253\,
            I => \N__7247\
        );

    \I__1437\ : Span4Mux_h
    port map (
            O => \N__7250\,
            I => \N__7244\
        );

    \I__1436\ : Span12Mux_h
    port map (
            O => \N__7247\,
            I => \N__7239\
        );

    \I__1435\ : Sp12to4
    port map (
            O => \N__7244\,
            I => \N__7239\
        );

    \I__1434\ : Span12Mux_v
    port map (
            O => \N__7239\,
            I => \N__7236\
        );

    \I__1433\ : Odrv12
    port map (
            O => \N__7236\,
            I => \D_in_6\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7233\,
            I => \N__7229\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7232\,
            I => \N__7226\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__7229\,
            I => \ATA_BASE_2\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7226\,
            I => \ATA_BASE_2\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__7221\,
            I => \N__7217\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7220\,
            I => \N__7214\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7217\,
            I => \N__7211\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7214\,
            I => \N__7208\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7211\,
            I => \U409_ADDRESS_DECODE.LOWROMZ0Z_3\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__7208\,
            I => \U409_ADDRESS_DECODE.LOWROMZ0Z_3\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7203\,
            I => \N__7197\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7202\,
            I => \N__7197\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7197\,
            I => \N__7193\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7196\,
            I => \N__7190\
        );

    \I__1418\ : Span4Mux_v
    port map (
            O => \N__7193\,
            I => \N__7186\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__7190\,
            I => \N__7183\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7180\
        );

    \I__1415\ : Odrv4
    port map (
            O => \N__7186\,
            I => \U409_ADDRESS_DECODE_ROMEN_1\
        );

    \I__1414\ : Odrv12
    port map (
            O => \N__7183\,
            I => \U409_ADDRESS_DECODE_ROMEN_1\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7180\,
            I => \U409_ADDRESS_DECODE_ROMEN_1\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__7173\,
            I => \N__7170\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7170\,
            I => \N__7163\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7169\,
            I => \N__7154\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7168\,
            I => \N__7154\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7151\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__7166\,
            I => \N__7147\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7163\,
            I => \N__7143\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7162\,
            I => \N__7140\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7161\,
            I => \N__7137\
        );

    \I__1403\ : InMux
    port map (
            O => \N__7160\,
            I => \N__7134\
        );

    \I__1402\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7131\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7154\,
            I => \N__7126\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7151\,
            I => \N__7126\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7150\,
            I => \N__7123\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7147\,
            I => \N__7120\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7146\,
            I => \N__7117\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__7143\,
            I => \N__7114\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7140\,
            I => \N__7105\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7137\,
            I => \N__7105\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7134\,
            I => \N__7105\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7131\,
            I => \N__7105\
        );

    \I__1391\ : Span4Mux_v
    port map (
            O => \N__7126\,
            I => \N__7102\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7123\,
            I => \N__7095\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7120\,
            I => \N__7095\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__7117\,
            I => \N__7095\
        );

    \I__1387\ : Span4Mux_h
    port map (
            O => \N__7114\,
            I => \N__7090\
        );

    \I__1386\ : Span4Mux_v
    port map (
            O => \N__7105\,
            I => \N__7090\
        );

    \I__1385\ : Span4Mux_h
    port map (
            O => \N__7102\,
            I => \N__7085\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__7095\,
            I => \N__7085\
        );

    \I__1383\ : Sp12to4
    port map (
            O => \N__7090\,
            I => \N__7080\
        );

    \I__1382\ : Sp12to4
    port map (
            O => \N__7085\,
            I => \N__7080\
        );

    \I__1381\ : Odrv12
    port map (
            O => \N__7080\,
            I => \A_c_21\
        );

    \I__1380\ : InMux
    port map (
            O => \N__7077\,
            I => \N__7074\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__7074\,
            I => \N__7070\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7073\,
            I => \N__7067\
        );

    \I__1377\ : Span4Mux_h
    port map (
            O => \N__7070\,
            I => \N__7061\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__7067\,
            I => \N__7061\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7066\,
            I => \N__7058\
        );

    \I__1374\ : Span4Mux_v
    port map (
            O => \N__7061\,
            I => \N__7055\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7058\,
            I => \N__7052\
        );

    \I__1372\ : Sp12to4
    port map (
            O => \N__7055\,
            I => \N__7049\
        );

    \I__1371\ : Span12Mux_h
    port map (
            O => \N__7052\,
            I => \N__7046\
        );

    \I__1370\ : Span12Mux_h
    port map (
            O => \N__7049\,
            I => \N__7043\
        );

    \I__1369\ : Span12Mux_v
    port map (
            O => \N__7046\,
            I => \N__7040\
        );

    \I__1368\ : Span12Mux_v
    port map (
            O => \N__7043\,
            I => \N__7037\
        );

    \I__1367\ : Odrv12
    port map (
            O => \N__7040\,
            I => \OVL_c\
        );

    \I__1366\ : Odrv12
    port map (
            O => \N__7037\,
            I => \OVL_c\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7032\,
            I => \N__7028\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7024\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__7028\,
            I => \N__7021\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7027\,
            I => \N__7018\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7024\,
            I => \N__7015\
        );

    \I__1360\ : Span4Mux_h
    port map (
            O => \N__7021\,
            I => \N__7012\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7018\,
            I => \N__7009\
        );

    \I__1358\ : Span12Mux_h
    port map (
            O => \N__7015\,
            I => \N__7006\
        );

    \I__1357\ : Sp12to4
    port map (
            O => \N__7012\,
            I => \N__7001\
        );

    \I__1356\ : Sp12to4
    port map (
            O => \N__7009\,
            I => \N__7001\
        );

    \I__1355\ : Span12Mux_v
    port map (
            O => \N__7006\,
            I => \N__6998\
        );

    \I__1354\ : Span12Mux_v
    port map (
            O => \N__7001\,
            I => \N__6995\
        );

    \I__1353\ : Odrv12
    port map (
            O => \N__6998\,
            I => \A_c_28\
        );

    \I__1352\ : Odrv12
    port map (
            O => \N__6995\,
            I => \A_c_28\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__6990\,
            I => \N__6987\
        );

    \I__1350\ : InMux
    port map (
            O => \N__6987\,
            I => \N__6983\
        );

    \I__1349\ : CascadeMux
    port map (
            O => \N__6986\,
            I => \N__6980\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__6983\,
            I => \N__6977\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6980\,
            I => \N__6974\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__6977\,
            I => \BRIDGE_BASE_0\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__6974\,
            I => \BRIDGE_BASE_0\
        );

    \I__1344\ : InMux
    port map (
            O => \N__6969\,
            I => \N__6966\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__6966\,
            I => \N__6963\
        );

    \I__1342\ : Span4Mux_v
    port map (
            O => \N__6963\,
            I => \N__6960\
        );

    \I__1341\ : Odrv4
    port map (
            O => \N__6960\,
            I => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_3\
        );

    \I__1340\ : IoInMux
    port map (
            O => \N__6957\,
            I => \N__6954\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__6954\,
            I => \N__6951\
        );

    \I__1338\ : IoSpan4Mux
    port map (
            O => \N__6951\,
            I => \N__6948\
        );

    \I__1337\ : Span4Mux_s3_h
    port map (
            O => \N__6948\,
            I => \N__6945\
        );

    \I__1336\ : Sp12to4
    port map (
            O => \N__6945\,
            I => \N__6942\
        );

    \I__1335\ : Span12Mux_h
    port map (
            O => \N__6942\,
            I => \N__6939\
        );

    \I__1334\ : Odrv12
    port map (
            O => \N__6939\,
            I => \U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__6936\,
            I => \N__6933\
        );

    \I__1332\ : InMux
    port map (
            O => \N__6933\,
            I => \N__6929\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6926\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__6929\,
            I => \N__6920\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6926\,
            I => \N__6917\
        );

    \I__1328\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6914\
        );

    \I__1327\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6911\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6908\
        );

    \I__1325\ : Span4Mux_v
    port map (
            O => \N__6920\,
            I => \N__6903\
        );

    \I__1324\ : Span4Mux_v
    port map (
            O => \N__6917\,
            I => \N__6900\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__6914\,
            I => \N__6897\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6911\,
            I => \N__6894\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6908\,
            I => \N__6890\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6907\,
            I => \N__6887\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6906\,
            I => \N__6884\
        );

    \I__1318\ : Span4Mux_h
    port map (
            O => \N__6903\,
            I => \N__6875\
        );

    \I__1317\ : Span4Mux_h
    port map (
            O => \N__6900\,
            I => \N__6875\
        );

    \I__1316\ : Span4Mux_v
    port map (
            O => \N__6897\,
            I => \N__6875\
        );

    \I__1315\ : Span4Mux_v
    port map (
            O => \N__6894\,
            I => \N__6875\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6872\
        );

    \I__1313\ : Span4Mux_v
    port map (
            O => \N__6890\,
            I => \N__6869\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6887\,
            I => \N__6866\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6884\,
            I => \N__6859\
        );

    \I__1310\ : Sp12to4
    port map (
            O => \N__6875\,
            I => \N__6859\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6872\,
            I => \N__6859\
        );

    \I__1308\ : Sp12to4
    port map (
            O => \N__6869\,
            I => \N__6854\
        );

    \I__1307\ : Span12Mux_v
    port map (
            O => \N__6866\,
            I => \N__6854\
        );

    \I__1306\ : Span12Mux_h
    port map (
            O => \N__6859\,
            I => \N__6851\
        );

    \I__1305\ : Odrv12
    port map (
            O => \N__6854\,
            I => \A_c_20\
        );

    \I__1304\ : Odrv12
    port map (
            O => \N__6851\,
            I => \A_c_20\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6843\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__6843\,
            I => \U409_ADDRESS_DECODE.ATA_SPACE_1Z0Z_0\
        );

    \I__1301\ : IoInMux
    port map (
            O => \N__6840\,
            I => \N__6837\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6837\,
            I => \N__6834\
        );

    \I__1299\ : IoSpan4Mux
    port map (
            O => \N__6834\,
            I => \N__6831\
        );

    \I__1298\ : Span4Mux_s2_v
    port map (
            O => \N__6831\,
            I => \N__6828\
        );

    \I__1297\ : Sp12to4
    port map (
            O => \N__6828\,
            I => \N__6825\
        );

    \I__1296\ : Span12Mux_v
    port map (
            O => \N__6825\,
            I => \N__6822\
        );

    \I__1295\ : Odrv12
    port map (
            O => \N__6822\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6816\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6816\,
            I => \N__6813\
        );

    \I__1292\ : Odrv12
    port map (
            O => \N__6813\,
            I => \U409_ADDRESS_DECODE_un1_ROMEN_0\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6810\,
            I => \N__6807\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__6807\,
            I => \N__6802\
        );

    \I__1289\ : InMux
    port map (
            O => \N__6806\,
            I => \N__6799\
        );

    \I__1288\ : InMux
    port map (
            O => \N__6805\,
            I => \N__6796\
        );

    \I__1287\ : Odrv12
    port map (
            O => \N__6802\,
            I => \U409_ADDRESS_DECODE.ATA_ENZ0\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__6799\,
            I => \U409_ADDRESS_DECODE.ATA_ENZ0\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__6796\,
            I => \U409_ADDRESS_DECODE.ATA_ENZ0\
        );

    \I__1284\ : IoInMux
    port map (
            O => \N__6789\,
            I => \N__6786\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6786\,
            I => \N__6783\
        );

    \I__1282\ : IoSpan4Mux
    port map (
            O => \N__6783\,
            I => \N__6780\
        );

    \I__1281\ : Sp12to4
    port map (
            O => \N__6780\,
            I => \N__6777\
        );

    \I__1280\ : Span12Mux_s7_h
    port map (
            O => \N__6777\,
            I => \N__6774\
        );

    \I__1279\ : Span12Mux_h
    port map (
            O => \N__6774\,
            I => \N__6771\
        );

    \I__1278\ : Odrv12
    port map (
            O => \N__6771\,
            I => \U409_ADDRESS_DECODE_un1_ATA_ENn_i\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6762\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6767\,
            I => \N__6762\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6762\,
            I => \U409_TRANSFER_ACK.CO1\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6759\,
            I => \N__6755\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6758\,
            I => \N__6752\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6755\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__6752\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6741\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6746\,
            I => \N__6741\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6741\,
            I => \N__6738\
        );

    \I__1267\ : Odrv4
    port map (
            O => \N__6738\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__6735\,
            I => \N__6732\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6732\,
            I => \N__6728\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6725\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__6728\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__6725\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__6720\,
            I => \N__6717\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6717\,
            I => \N__6711\
        );

    \I__1259\ : InMux
    port map (
            O => \N__6716\,
            I => \N__6711\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__6711\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__6708\,
            I => \N__6705\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6705\,
            I => \N__6702\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6702\,
            I => \N__6699\
        );

    \I__1254\ : Span4Mux_v
    port map (
            O => \N__6699\,
            I => \N__6694\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__6698\,
            I => \N__6691\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__6697\,
            I => \N__6688\
        );

    \I__1251\ : Span4Mux_h
    port map (
            O => \N__6694\,
            I => \N__6685\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6680\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6688\,
            I => \N__6680\
        );

    \I__1248\ : Sp12to4
    port map (
            O => \N__6685\,
            I => \N__6677\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6680\,
            I => \N__6674\
        );

    \I__1246\ : Span12Mux_h
    port map (
            O => \N__6677\,
            I => \N__6669\
        );

    \I__1245\ : Span12Mux_h
    port map (
            O => \N__6674\,
            I => \N__6669\
        );

    \I__1244\ : Span12Mux_v
    port map (
            O => \N__6669\,
            I => \N__6666\
        );

    \I__1243\ : Odrv12
    port map (
            O => \N__6666\,
            I => \D_in_7\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6663\,
            I => \N__6660\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6660\,
            I => \N__6656\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6659\,
            I => \N__6653\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__6656\,
            I => \BRIDGE_BASE_3\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6653\,
            I => \BRIDGE_BASE_3\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6648\,
            I => \N__6645\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6645\,
            I => \N__6641\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__6644\,
            I => \N__6638\
        );

    \I__1234\ : Span4Mux_v
    port map (
            O => \N__6641\,
            I => \N__6635\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6638\,
            I => \N__6632\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__6635\,
            I => \BRIDGE_BASE_2\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__6632\,
            I => \BRIDGE_BASE_2\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6627\,
            I => \N__6624\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__6624\,
            I => \N__6621\
        );

    \I__1228\ : Span12Mux_v
    port map (
            O => \N__6621\,
            I => \N__6617\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6620\,
            I => \N__6614\
        );

    \I__1226\ : Odrv12
    port map (
            O => \N__6617\,
            I => \BRIDGE_BASE_1\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6614\,
            I => \BRIDGE_BASE_1\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6609\,
            I => \N__6603\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6608\,
            I => \N__6596\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6596\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6606\,
            I => \N__6596\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6603\,
            I => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6596\,
            I => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6591\,
            I => \N__6585\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__6590\,
            I => \N__6581\
        );

    \I__1216\ : CascadeMux
    port map (
            O => \N__6589\,
            I => \N__6577\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6588\,
            I => \N__6570\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6585\,
            I => \N__6567\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6584\,
            I => \N__6564\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6561\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6558\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6553\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6553\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6575\,
            I => \N__6550\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6574\,
            I => \N__6547\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6573\,
            I => \N__6544\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6570\,
            I => \N__6541\
        );

    \I__1204\ : Span4Mux_h
    port map (
            O => \N__6567\,
            I => \N__6528\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6564\,
            I => \N__6528\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6561\,
            I => \N__6528\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6558\,
            I => \N__6528\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6553\,
            I => \N__6528\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6550\,
            I => \N__6528\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6547\,
            I => \N__6523\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6544\,
            I => \N__6523\
        );

    \I__1196\ : Span4Mux_v
    port map (
            O => \N__6541\,
            I => \N__6520\
        );

    \I__1195\ : Span4Mux_v
    port map (
            O => \N__6528\,
            I => \N__6517\
        );

    \I__1194\ : Span4Mux_v
    port map (
            O => \N__6523\,
            I => \N__6514\
        );

    \I__1193\ : Sp12to4
    port map (
            O => \N__6520\,
            I => \N__6507\
        );

    \I__1192\ : Sp12to4
    port map (
            O => \N__6517\,
            I => \N__6507\
        );

    \I__1191\ : Sp12to4
    port map (
            O => \N__6514\,
            I => \N__6507\
        );

    \I__1190\ : Odrv12
    port map (
            O => \N__6507\,
            I => \A_c_23\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6504\,
            I => \N__6500\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6497\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__6500\,
            I => \ATA_BASE_7\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6497\,
            I => \ATA_BASE_7\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__6492\,
            I => \N__6488\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6482\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6488\,
            I => \N__6475\
        );

    \I__1182\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6472\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6469\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6466\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6482\,
            I => \N__6463\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6460\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6457\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6454\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__6478\,
            I => \N__6451\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6475\,
            I => \N__6442\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__6472\,
            I => \N__6442\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6469\,
            I => \N__6442\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6466\,
            I => \N__6442\
        );

    \I__1170\ : Span4Mux_v
    port map (
            O => \N__6463\,
            I => \N__6439\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6460\,
            I => \N__6432\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6457\,
            I => \N__6432\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__6454\,
            I => \N__6432\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6451\,
            I => \N__6429\
        );

    \I__1165\ : Span4Mux_v
    port map (
            O => \N__6442\,
            I => \N__6426\
        );

    \I__1164\ : Span4Mux_h
    port map (
            O => \N__6439\,
            I => \N__6421\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__6432\,
            I => \N__6421\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6429\,
            I => \N__6418\
        );

    \I__1161\ : Span4Mux_v
    port map (
            O => \N__6426\,
            I => \N__6415\
        );

    \I__1160\ : Span4Mux_v
    port map (
            O => \N__6421\,
            I => \N__6412\
        );

    \I__1159\ : Span12Mux_h
    port map (
            O => \N__6418\,
            I => \N__6409\
        );

    \I__1158\ : Span4Mux_v
    port map (
            O => \N__6415\,
            I => \N__6406\
        );

    \I__1157\ : Span4Mux_v
    port map (
            O => \N__6412\,
            I => \N__6403\
        );

    \I__1156\ : Span12Mux_v
    port map (
            O => \N__6409\,
            I => \N__6400\
        );

    \I__1155\ : Sp12to4
    port map (
            O => \N__6406\,
            I => \N__6395\
        );

    \I__1154\ : Sp12to4
    port map (
            O => \N__6403\,
            I => \N__6395\
        );

    \I__1153\ : Odrv12
    port map (
            O => \N__6400\,
            I => \A_c_22\
        );

    \I__1152\ : Odrv12
    port map (
            O => \N__6395\,
            I => \A_c_22\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6387\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6387\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6384\,
            I => \N__6376\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6383\,
            I => \N__6373\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__6382\,
            I => \N__6368\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6381\,
            I => \N__6363\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6380\,
            I => \N__6363\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__6379\,
            I => \N__6354\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__6376\,
            I => \N__6346\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__6373\,
            I => \N__6346\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6343\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6336\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6336\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6363\,
            I => \N__6333\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6326\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6326\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6360\,
            I => \N__6326\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6321\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6321\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6314\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6354\,
            I => \N__6314\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6353\,
            I => \N__6314\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6311\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6351\,
            I => \N__6308\
        );

    \I__1127\ : Span4Mux_h
    port map (
            O => \N__6346\,
            I => \N__6303\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6343\,
            I => \N__6303\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6342\,
            I => \N__6300\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6341\,
            I => \N__6297\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6336\,
            I => \N__6294\
        );

    \I__1122\ : Span4Mux_v
    port map (
            O => \N__6333\,
            I => \N__6291\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6326\,
            I => \N__6286\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__6321\,
            I => \N__6286\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6314\,
            I => \N__6279\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6311\,
            I => \N__6279\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__6308\,
            I => \N__6279\
        );

    \I__1116\ : Span4Mux_h
    port map (
            O => \N__6303\,
            I => \N__6272\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__6300\,
            I => \N__6272\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6297\,
            I => \N__6272\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__6294\,
            I => \N__6269\
        );

    \I__1112\ : Span4Mux_h
    port map (
            O => \N__6291\,
            I => \N__6262\
        );

    \I__1111\ : Span4Mux_v
    port map (
            O => \N__6286\,
            I => \N__6262\
        );

    \I__1110\ : Span4Mux_v
    port map (
            O => \N__6279\,
            I => \N__6262\
        );

    \I__1109\ : Span4Mux_v
    port map (
            O => \N__6272\,
            I => \N__6259\
        );

    \I__1108\ : Span4Mux_v
    port map (
            O => \N__6269\,
            I => \N__6256\
        );

    \I__1107\ : Span4Mux_v
    port map (
            O => \N__6262\,
            I => \N__6253\
        );

    \I__1106\ : Span4Mux_h
    port map (
            O => \N__6259\,
            I => \N__6250\
        );

    \I__1105\ : Sp12to4
    port map (
            O => \N__6256\,
            I => \N__6245\
        );

    \I__1104\ : Sp12to4
    port map (
            O => \N__6253\,
            I => \N__6245\
        );

    \I__1103\ : Sp12to4
    port map (
            O => \N__6250\,
            I => \N__6242\
        );

    \I__1102\ : Span12Mux_h
    port map (
            O => \N__6245\,
            I => \N__6239\
        );

    \I__1101\ : Span12Mux_v
    port map (
            O => \N__6242\,
            I => \N__6236\
        );

    \I__1100\ : Odrv12
    port map (
            O => \N__6239\,
            I => \A_c_1\
        );

    \I__1099\ : Odrv12
    port map (
            O => \N__6236\,
            I => \A_c_1\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__6231\,
            I => \N__6227\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__6230\,
            I => \N__6223\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6227\,
            I => \N__6220\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__6226\,
            I => \N__6217\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6223\,
            I => \N__6207\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6220\,
            I => \N__6204\
        );

    \I__1092\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6201\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6216\,
            I => \N__6196\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6196\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6191\
        );

    \I__1088\ : InMux
    port map (
            O => \N__6213\,
            I => \N__6191\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6212\,
            I => \N__6184\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6211\,
            I => \N__6184\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6210\,
            I => \N__6184\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6207\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1083\ : Odrv4
    port map (
            O => \N__6204\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__6201\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__6196\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__6191\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6184\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1078\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6168\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6168\,
            I => \N__6160\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6155\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6155\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6165\,
            I => \N__6150\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6164\,
            I => \N__6150\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6163\,
            I => \N__6147\
        );

    \I__1071\ : Span4Mux_v
    port map (
            O => \N__6160\,
            I => \N__6140\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__6155\,
            I => \N__6140\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6150\,
            I => \N__6140\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6147\,
            I => \U409_AUTOCONFIG.N_122\
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__6140\,
            I => \U409_AUTOCONFIG.N_122\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6135\,
            I => \N__6128\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6134\,
            I => \N__6125\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6122\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6132\,
            I => \N__6119\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6131\,
            I => \N__6116\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__6128\,
            I => \N__6111\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6125\,
            I => \N__6106\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6122\,
            I => \N__6106\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6119\,
            I => \N__6101\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6116\,
            I => \N__6101\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6115\,
            I => \N__6098\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6114\,
            I => \N__6095\
        );

    \I__1054\ : Span4Mux_h
    port map (
            O => \N__6111\,
            I => \N__6090\
        );

    \I__1053\ : Span4Mux_v
    port map (
            O => \N__6106\,
            I => \N__6090\
        );

    \I__1052\ : Span4Mux_h
    port map (
            O => \N__6101\,
            I => \N__6083\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6098\,
            I => \N__6083\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6095\,
            I => \N__6083\
        );

    \I__1049\ : Span4Mux_v
    port map (
            O => \N__6090\,
            I => \N__6080\
        );

    \I__1048\ : Span4Mux_v
    port map (
            O => \N__6083\,
            I => \N__6077\
        );

    \I__1047\ : Sp12to4
    port map (
            O => \N__6080\,
            I => \N__6072\
        );

    \I__1046\ : Sp12to4
    port map (
            O => \N__6077\,
            I => \N__6072\
        );

    \I__1045\ : Span12Mux_h
    port map (
            O => \N__6072\,
            I => \N__6069\
        );

    \I__1044\ : Span12Mux_v
    port map (
            O => \N__6069\,
            I => \N__6066\
        );

    \I__1043\ : Odrv12
    port map (
            O => \N__6066\,
            I => \A_c_19\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6063\,
            I => \N__6059\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6062\,
            I => \N__6056\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6059\,
            I => \ATA_BASE_3\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__6056\,
            I => \ATA_BASE_3\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__6051\,
            I => \N__6048\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6048\,
            I => \N__6042\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6047\,
            I => \N__6039\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6046\,
            I => \N__6036\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6033\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6042\,
            I => \N__6029\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6039\,
            I => \N__6022\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6036\,
            I => \N__6022\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6033\,
            I => \N__6022\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__6032\,
            I => \N__6019\
        );

    \I__1028\ : Span4Mux_v
    port map (
            O => \N__6029\,
            I => \N__6016\
        );

    \I__1027\ : Span4Mux_v
    port map (
            O => \N__6022\,
            I => \N__6013\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6019\,
            I => \N__6010\
        );

    \I__1025\ : Sp12to4
    port map (
            O => \N__6016\,
            I => \N__6003\
        );

    \I__1024\ : Sp12to4
    port map (
            O => \N__6013\,
            I => \N__6003\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6010\,
            I => \N__6003\
        );

    \I__1022\ : Span12Mux_h
    port map (
            O => \N__6003\,
            I => \N__6000\
        );

    \I__1021\ : Span12Mux_v
    port map (
            O => \N__6000\,
            I => \N__5997\
        );

    \I__1020\ : Odrv12
    port map (
            O => \N__5997\,
            I => \A_c_18\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5994\,
            I => \N__5991\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5991\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2\
        );

    \I__1017\ : InMux
    port map (
            O => \N__5988\,
            I => \N__5985\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5985\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__5982\,
            I => \N__5977\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5974\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5971\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5977\,
            I => \N__5968\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5974\,
            I => \N__5965\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__5971\,
            I => \N__5962\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5968\,
            I => \N__5959\
        );

    \I__1008\ : Span4Mux_v
    port map (
            O => \N__5965\,
            I => \N__5956\
        );

    \I__1007\ : Span4Mux_h
    port map (
            O => \N__5962\,
            I => \N__5953\
        );

    \I__1006\ : Span12Mux_v
    port map (
            O => \N__5959\,
            I => \N__5950\
        );

    \I__1005\ : Sp12to4
    port map (
            O => \N__5956\,
            I => \N__5947\
        );

    \I__1004\ : Span4Mux_v
    port map (
            O => \N__5953\,
            I => \N__5944\
        );

    \I__1003\ : Odrv12
    port map (
            O => \N__5950\,
            I => \A_c_31\
        );

    \I__1002\ : Odrv12
    port map (
            O => \N__5947\,
            I => \A_c_31\
        );

    \I__1001\ : Odrv4
    port map (
            O => \N__5944\,
            I => \A_c_31\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5937\,
            I => \N__5934\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5934\,
            I => \N_120\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__5931\,
            I => \U409_ADDRESS_DECODE.PORTSIZEZ0Z_0_cascade_\
        );

    \I__997\ : IoInMux
    port map (
            O => \N__5928\,
            I => \N__5925\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5925\,
            I => \N__5922\
        );

    \I__995\ : Span4Mux_s2_v
    port map (
            O => \N__5922\,
            I => \N__5919\
        );

    \I__994\ : Span4Mux_h
    port map (
            O => \N__5919\,
            I => \N__5916\
        );

    \I__993\ : Span4Mux_v
    port map (
            O => \N__5916\,
            I => \N__5913\
        );

    \I__992\ : Span4Mux_v
    port map (
            O => \N__5913\,
            I => \N__5910\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__5910\,
            I => \PORTSIZE_0_i\
        );

    \I__990\ : InMux
    port map (
            O => \N__5907\,
            I => \N__5904\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__5904\,
            I => \N__5899\
        );

    \I__988\ : CascadeMux
    port map (
            O => \N__5903\,
            I => \N__5896\
        );

    \I__987\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5893\
        );

    \I__986\ : Span4Mux_v
    port map (
            O => \N__5899\,
            I => \N__5890\
        );

    \I__985\ : InMux
    port map (
            O => \N__5896\,
            I => \N__5887\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5893\,
            I => \N__5884\
        );

    \I__983\ : Span4Mux_h
    port map (
            O => \N__5890\,
            I => \N__5879\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5887\,
            I => \N__5879\
        );

    \I__981\ : Span4Mux_v
    port map (
            O => \N__5884\,
            I => \N__5876\
        );

    \I__980\ : Span4Mux_h
    port map (
            O => \N__5879\,
            I => \N__5873\
        );

    \I__979\ : Sp12to4
    port map (
            O => \N__5876\,
            I => \N__5870\
        );

    \I__978\ : Span4Mux_v
    port map (
            O => \N__5873\,
            I => \N__5867\
        );

    \I__977\ : Odrv12
    port map (
            O => \N__5870\,
            I => \A_c_30\
        );

    \I__976\ : Odrv4
    port map (
            O => \N__5867\,
            I => \A_c_30\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__5862\,
            I => \N__5859\
        );

    \I__974\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5856\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__5856\,
            I => \N__5853\
        );

    \I__972\ : Span4Mux_h
    port map (
            O => \N__5853\,
            I => \N__5849\
        );

    \I__971\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5846\
        );

    \I__970\ : Span4Mux_h
    port map (
            O => \N__5849\,
            I => \N__5840\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5846\,
            I => \N__5840\
        );

    \I__968\ : InMux
    port map (
            O => \N__5845\,
            I => \N__5837\
        );

    \I__967\ : Span4Mux_v
    port map (
            O => \N__5840\,
            I => \N__5834\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5837\,
            I => \N__5831\
        );

    \I__965\ : Span4Mux_v
    port map (
            O => \N__5834\,
            I => \N__5828\
        );

    \I__964\ : Span12Mux_v
    port map (
            O => \N__5831\,
            I => \N__5823\
        );

    \I__963\ : Sp12to4
    port map (
            O => \N__5828\,
            I => \N__5823\
        );

    \I__962\ : Odrv12
    port map (
            O => \N__5823\,
            I => \A_c_29\
        );

    \I__961\ : InMux
    port map (
            O => \N__5820\,
            I => \N__5817\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5817\,
            I => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_0\
        );

    \I__959\ : IoInMux
    port map (
            O => \N__5814\,
            I => \N__5811\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5811\,
            I => \N__5808\
        );

    \I__957\ : Span12Mux_s10_v
    port map (
            O => \N__5808\,
            I => \N__5805\
        );

    \I__956\ : Span12Mux_h
    port map (
            O => \N__5805\,
            I => \N__5801\
        );

    \I__955\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5798\
        );

    \I__954\ : Odrv12
    port map (
            O => \N__5801\,
            I => \CONFIGENn_c\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5798\,
            I => \CONFIGENn_c\
        );

    \I__952\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5786\
        );

    \I__951\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5777\
        );

    \I__950\ : InMux
    port map (
            O => \N__5791\,
            I => \N__5777\
        );

    \I__949\ : InMux
    port map (
            O => \N__5790\,
            I => \N__5777\
        );

    \I__948\ : InMux
    port map (
            O => \N__5789\,
            I => \N__5777\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__5786\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5777\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__945\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5765\
        );

    \I__944\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5756\
        );

    \I__943\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5756\
        );

    \I__942\ : InMux
    port map (
            O => \N__5769\,
            I => \N__5756\
        );

    \I__941\ : InMux
    port map (
            O => \N__5768\,
            I => \N__5756\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5765\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5756\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__938\ : InMux
    port map (
            O => \N__5751\,
            I => \N__5746\
        );

    \I__937\ : InMux
    port map (
            O => \N__5750\,
            I => \N__5741\
        );

    \I__936\ : InMux
    port map (
            O => \N__5749\,
            I => \N__5741\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5746\,
            I => \N__5738\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5741\,
            I => \N__5735\
        );

    \I__933\ : Span4Mux_v
    port map (
            O => \N__5738\,
            I => \N__5729\
        );

    \I__932\ : Span4Mux_v
    port map (
            O => \N__5735\,
            I => \N__5729\
        );

    \I__931\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5726\
        );

    \I__930\ : Sp12to4
    port map (
            O => \N__5729\,
            I => \N__5721\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5726\,
            I => \N__5721\
        );

    \I__928\ : Span12Mux_h
    port map (
            O => \N__5721\,
            I => \N__5718\
        );

    \I__927\ : Span12Mux_v
    port map (
            O => \N__5718\,
            I => \N__5715\
        );

    \I__926\ : Odrv12
    port map (
            O => \N__5715\,
            I => \TM_c_0\
        );

    \I__925\ : InMux
    port map (
            O => \N__5712\,
            I => \N__5707\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__5711\,
            I => \N__5700\
        );

    \I__923\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5697\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__5707\,
            I => \N__5694\
        );

    \I__921\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5689\
        );

    \I__920\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5689\
        );

    \I__919\ : InMux
    port map (
            O => \N__5704\,
            I => \N__5686\
        );

    \I__918\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5683\
        );

    \I__917\ : InMux
    port map (
            O => \N__5700\,
            I => \N__5680\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5697\,
            I => \CONFIGURED\
        );

    \I__915\ : Odrv4
    port map (
            O => \N__5694\,
            I => \CONFIGURED\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5689\,
            I => \CONFIGURED\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5686\,
            I => \CONFIGURED\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__5683\,
            I => \CONFIGURED\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5680\,
            I => \CONFIGURED\
        );

    \I__910\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5660\
        );

    \I__909\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5660\
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__5665\,
            I => \N__5657\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5660\,
            I => \N__5653\
        );

    \I__906\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5650\
        );

    \I__905\ : InMux
    port map (
            O => \N__5656\,
            I => \N__5647\
        );

    \I__904\ : Span4Mux_v
    port map (
            O => \N__5653\,
            I => \N__5642\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5650\,
            I => \N__5642\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5647\,
            I => \N__5639\
        );

    \I__901\ : Span4Mux_h
    port map (
            O => \N__5642\,
            I => \N__5636\
        );

    \I__900\ : Span12Mux_h
    port map (
            O => \N__5639\,
            I => \N__5631\
        );

    \I__899\ : Sp12to4
    port map (
            O => \N__5636\,
            I => \N__5631\
        );

    \I__898\ : Span12Mux_v
    port map (
            O => \N__5631\,
            I => \N__5628\
        );

    \I__897\ : Odrv12
    port map (
            O => \N__5628\,
            I => \TM_c_1\
        );

    \I__896\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5621\
        );

    \I__895\ : InMux
    port map (
            O => \N__5624\,
            I => \N__5618\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__5621\,
            I => \N__5614\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5618\,
            I => \N__5611\
        );

    \I__892\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5607\
        );

    \I__891\ : Span4Mux_v
    port map (
            O => \N__5614\,
            I => \N__5604\
        );

    \I__890\ : Span4Mux_v
    port map (
            O => \N__5611\,
            I => \N__5601\
        );

    \I__889\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5598\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5607\,
            I => \N__5595\
        );

    \I__887\ : Sp12to4
    port map (
            O => \N__5604\,
            I => \N__5588\
        );

    \I__886\ : Sp12to4
    port map (
            O => \N__5601\,
            I => \N__5588\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5598\,
            I => \N__5588\
        );

    \I__884\ : Span12Mux_v
    port map (
            O => \N__5595\,
            I => \N__5585\
        );

    \I__883\ : Span12Mux_h
    port map (
            O => \N__5588\,
            I => \N__5582\
        );

    \I__882\ : Span12Mux_v
    port map (
            O => \N__5585\,
            I => \N__5579\
        );

    \I__881\ : Span12Mux_v
    port map (
            O => \N__5582\,
            I => \N__5576\
        );

    \I__880\ : Odrv12
    port map (
            O => \N__5579\,
            I => \A_c_17\
        );

    \I__879\ : Odrv12
    port map (
            O => \N__5576\,
            I => \A_c_17\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__5571\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_\
        );

    \I__877\ : InMux
    port map (
            O => \N__5568\,
            I => \N__5564\
        );

    \I__876\ : InMux
    port map (
            O => \N__5567\,
            I => \N__5561\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5564\,
            I => \ATA_BASE_1\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5561\,
            I => \ATA_BASE_1\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__5556\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4_cascade_\
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__5553\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__5550\,
            I => \N__5546\
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__5549\,
            I => \N__5540\
        );

    \I__869\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5536\
        );

    \I__868\ : InMux
    port map (
            O => \N__5545\,
            I => \N__5531\
        );

    \I__867\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5531\
        );

    \I__866\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5526\
        );

    \I__865\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5526\
        );

    \I__864\ : InMux
    port map (
            O => \N__5539\,
            I => \N__5523\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5536\,
            I => \N__5520\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5531\,
            I => \N__5517\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5526\,
            I => \N__5512\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__5523\,
            I => \N__5512\
        );

    \I__859\ : Span4Mux_v
    port map (
            O => \N__5520\,
            I => \N__5507\
        );

    \I__858\ : Span4Mux_v
    port map (
            O => \N__5517\,
            I => \N__5507\
        );

    \I__857\ : Span4Mux_v
    port map (
            O => \N__5512\,
            I => \N__5504\
        );

    \I__856\ : Sp12to4
    port map (
            O => \N__5507\,
            I => \N__5499\
        );

    \I__855\ : Sp12to4
    port map (
            O => \N__5504\,
            I => \N__5499\
        );

    \I__854\ : Span12Mux_h
    port map (
            O => \N__5499\,
            I => \N__5496\
        );

    \I__853\ : Span12Mux_v
    port map (
            O => \N__5496\,
            I => \N__5493\
        );

    \I__852\ : Odrv12
    port map (
            O => \N__5493\,
            I => \RnW_c\
        );

    \I__851\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5487\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5487\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_4\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__5484\,
            I => \N__5481\
        );

    \I__848\ : InMux
    port map (
            O => \N__5481\,
            I => \N__5473\
        );

    \I__847\ : InMux
    port map (
            O => \N__5480\,
            I => \N__5473\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__5479\,
            I => \N__5467\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__5478\,
            I => \N__5464\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5473\,
            I => \N__5461\
        );

    \I__843\ : InMux
    port map (
            O => \N__5472\,
            I => \N__5456\
        );

    \I__842\ : InMux
    port map (
            O => \N__5471\,
            I => \N__5456\
        );

    \I__841\ : InMux
    port map (
            O => \N__5470\,
            I => \N__5451\
        );

    \I__840\ : InMux
    port map (
            O => \N__5467\,
            I => \N__5451\
        );

    \I__839\ : InMux
    port map (
            O => \N__5464\,
            I => \N__5448\
        );

    \I__838\ : Span4Mux_v
    port map (
            O => \N__5461\,
            I => \N__5445\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5456\,
            I => \N__5438\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5451\,
            I => \N__5438\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__5448\,
            I => \N__5438\
        );

    \I__834\ : Span4Mux_h
    port map (
            O => \N__5445\,
            I => \N__5435\
        );

    \I__833\ : Span4Mux_v
    port map (
            O => \N__5438\,
            I => \N__5432\
        );

    \I__832\ : Odrv4
    port map (
            O => \N__5435\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE\
        );

    \I__831\ : Odrv4
    port map (
            O => \N__5432\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE\
        );

    \I__830\ : IoInMux
    port map (
            O => \N__5427\,
            I => \N__5424\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__5424\,
            I => \N__5421\
        );

    \I__828\ : IoSpan4Mux
    port map (
            O => \N__5421\,
            I => \N__5418\
        );

    \I__827\ : Span4Mux_s1_h
    port map (
            O => \N__5418\,
            I => \N__5415\
        );

    \I__826\ : Sp12to4
    port map (
            O => \N__5415\,
            I => \N__5412\
        );

    \I__825\ : Span12Mux_s6_h
    port map (
            O => \N__5412\,
            I => \N__5409\
        );

    \I__824\ : Span12Mux_h
    port map (
            O => \N__5409\,
            I => \N__5406\
        );

    \I__823\ : Span12Mux_v
    port map (
            O => \N__5406\,
            I => \N__5403\
        );

    \I__822\ : Odrv12
    port map (
            O => \N__5403\,
            I => \N_120_i\
        );

    \I__821\ : IoInMux
    port map (
            O => \N__5400\,
            I => \N__5397\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5397\,
            I => \N__5394\
        );

    \I__819\ : IoSpan4Mux
    port map (
            O => \N__5394\,
            I => \N__5391\
        );

    \I__818\ : Span4Mux_s3_v
    port map (
            O => \N__5391\,
            I => \N__5388\
        );

    \I__817\ : Span4Mux_h
    port map (
            O => \N__5388\,
            I => \N__5385\
        );

    \I__816\ : Sp12to4
    port map (
            O => \N__5385\,
            I => \N__5382\
        );

    \I__815\ : Span12Mux_v
    port map (
            O => \N__5382\,
            I => \N__5379\
        );

    \I__814\ : Odrv12
    port map (
            O => \N__5379\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\
        );

    \I__813\ : InMux
    port map (
            O => \N__5376\,
            I => \N__5370\
        );

    \I__812\ : InMux
    port map (
            O => \N__5375\,
            I => \N__5370\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5370\,
            I => \N__5367\
        );

    \I__810\ : Odrv4
    port map (
            O => \N__5367\,
            I => \U409_ADDRESS_DECODE.N_102\
        );

    \I__809\ : InMux
    port map (
            O => \N__5364\,
            I => \N__5358\
        );

    \I__808\ : InMux
    port map (
            O => \N__5363\,
            I => \N__5358\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__5358\,
            I => \N__5355\
        );

    \I__806\ : Odrv4
    port map (
            O => \N__5355\,
            I => \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3Z0Z_0\
        );

    \I__805\ : InMux
    port map (
            O => \N__5352\,
            I => \N__5349\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5349\,
            I => \N__5346\
        );

    \I__803\ : Span4Mux_v
    port map (
            O => \N__5346\,
            I => \N__5342\
        );

    \I__802\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5339\
        );

    \I__801\ : Odrv4
    port map (
            O => \N__5342\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__5339\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\
        );

    \I__799\ : InMux
    port map (
            O => \N__5334\,
            I => \N__5330\
        );

    \I__798\ : CascadeMux
    port map (
            O => \N__5333\,
            I => \N__5327\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5330\,
            I => \N__5324\
        );

    \I__796\ : InMux
    port map (
            O => \N__5327\,
            I => \N__5321\
        );

    \I__795\ : Odrv4
    port map (
            O => \N__5324\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5321\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\
        );

    \I__793\ : IoInMux
    port map (
            O => \N__5316\,
            I => \N__5313\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5313\,
            I => \N__5310\
        );

    \I__791\ : Span12Mux_s5_v
    port map (
            O => \N__5310\,
            I => \N__5307\
        );

    \I__790\ : Odrv12
    port map (
            O => \N__5307\,
            I => \U409_AUTOCONFIG_D_OUT_0_i_1\
        );

    \I__789\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5300\
        );

    \I__788\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5297\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5300\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5297\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__5292\,
            I => \N__5289\
        );

    \I__784\ : InMux
    port map (
            O => \N__5289\,
            I => \N__5286\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5286\,
            I => \N__5282\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__5285\,
            I => \N__5279\
        );

    \I__781\ : Span4Mux_v
    port map (
            O => \N__5282\,
            I => \N__5276\
        );

    \I__780\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5273\
        );

    \I__779\ : Odrv4
    port map (
            O => \N__5276\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5273\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\
        );

    \I__777\ : IoInMux
    port map (
            O => \N__5268\,
            I => \N__5265\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5265\,
            I => \N__5262\
        );

    \I__775\ : Span12Mux_s10_v
    port map (
            O => \N__5262\,
            I => \N__5259\
        );

    \I__774\ : Odrv12
    port map (
            O => \N__5259\,
            I => \U409_AUTOCONFIG_D_OUT_0_i_2\
        );

    \I__773\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5252\
        );

    \I__772\ : InMux
    port map (
            O => \N__5255\,
            I => \N__5249\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5252\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5249\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__5244\,
            I => \N__5241\
        );

    \I__768\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__5238\,
            I => \N__5235\
        );

    \I__766\ : Span4Mux_v
    port map (
            O => \N__5235\,
            I => \N__5231\
        );

    \I__765\ : InMux
    port map (
            O => \N__5234\,
            I => \N__5228\
        );

    \I__764\ : Odrv4
    port map (
            O => \N__5231\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5228\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\
        );

    \I__762\ : IoInMux
    port map (
            O => \N__5223\,
            I => \N__5220\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__5220\,
            I => \N__5217\
        );

    \I__760\ : Span4Mux_s2_v
    port map (
            O => \N__5217\,
            I => \N__5214\
        );

    \I__759\ : Sp12to4
    port map (
            O => \N__5214\,
            I => \N__5211\
        );

    \I__758\ : Span12Mux_h
    port map (
            O => \N__5211\,
            I => \N__5208\
        );

    \I__757\ : Span12Mux_v
    port map (
            O => \N__5208\,
            I => \N__5205\
        );

    \I__756\ : Odrv12
    port map (
            O => \N__5205\,
            I => \U409_AUTOCONFIG_D_OUT_0_i_3\
        );

    \I__755\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5199\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5199\,
            I => \N__5196\
        );

    \I__753\ : Odrv12
    port map (
            O => \N__5196\,
            I => \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0Z0Z_0\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__5193\,
            I => \N__5189\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__5192\,
            I => \N__5185\
        );

    \I__750\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5175\
        );

    \I__749\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5175\
        );

    \I__748\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5175\
        );

    \I__747\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5175\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__5175\,
            I => \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa\
        );

    \I__745\ : InMux
    port map (
            O => \N__5172\,
            I => \N__5169\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5169\,
            I => \N__5166\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__5166\,
            I => \U409_ADDRESS_DECODE.HIROMZ0\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__5163\,
            I => \U409_ADDRESS_DECODE.LOWROMZ0Z_2_cascade_\
        );

    \I__741\ : IoInMux
    port map (
            O => \N__5160\,
            I => \N__5157\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5157\,
            I => \N__5152\
        );

    \I__739\ : IoInMux
    port map (
            O => \N__5156\,
            I => \N__5149\
        );

    \I__738\ : IoInMux
    port map (
            O => \N__5155\,
            I => \N__5146\
        );

    \I__737\ : IoSpan4Mux
    port map (
            O => \N__5152\,
            I => \N__5139\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__5149\,
            I => \N__5139\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__5146\,
            I => \N__5139\
        );

    \I__734\ : IoSpan4Mux
    port map (
            O => \N__5139\,
            I => \N__5136\
        );

    \I__733\ : Span4Mux_s2_v
    port map (
            O => \N__5136\,
            I => \N__5132\
        );

    \I__732\ : IoInMux
    port map (
            O => \N__5135\,
            I => \N__5129\
        );

    \I__731\ : Sp12to4
    port map (
            O => \N__5132\,
            I => \N__5124\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__5129\,
            I => \N__5124\
        );

    \I__729\ : Span12Mux_s10_v
    port map (
            O => \N__5124\,
            I => \N__5121\
        );

    \I__728\ : Odrv12
    port map (
            O => \N__5121\,
            I => \D_1_i\
        );

    \I__727\ : InMux
    port map (
            O => \N__5118\,
            I => \N__5115\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5115\,
            I => \U409_AUTOCONFIG.AC_STARTZ0\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__5112\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_1_cascade_\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__5109\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_4_cascade_\
        );

    \I__723\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5103\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__5103\,
            I => \N__5100\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__5100\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_10\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__5097\,
            I => \N_120_cascade_\
        );

    \I__719\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5091\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5091\,
            I => \N__5088\
        );

    \I__717\ : Span12Mux_h
    port map (
            O => \N__5088\,
            I => \N__5085\
        );

    \I__716\ : Odrv12
    port map (
            O => \N__5085\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_11\
        );

    \I__715\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__5079\,
            I => \N__5076\
        );

    \I__713\ : Span4Mux_h
    port map (
            O => \N__5076\,
            I => \N__5073\
        );

    \I__712\ : Odrv4
    port map (
            O => \N__5073\,
            I => \U409_AUTOCONFIG.N_31\
        );

    \I__711\ : InMux
    port map (
            O => \N__5070\,
            I => \N__5067\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5067\,
            I => \N__5064\
        );

    \I__709\ : Span4Mux_h
    port map (
            O => \N__5064\,
            I => \N__5061\
        );

    \I__708\ : Odrv4
    port map (
            O => \N__5061\,
            I => \U409_AUTOCONFIG.N_22\
        );

    \I__707\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5055\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5055\,
            I => \N__5052\
        );

    \I__705\ : Odrv12
    port map (
            O => \N__5052\,
            I => \U409_AUTOCONFIG.LIDE_CONF_1_sqmuxa_0_a2_0Z0Z_2\
        );

    \I__704\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5046\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5046\,
            I => \N__5043\
        );

    \I__702\ : Odrv4
    port map (
            O => \N__5043\,
            I => \U409_AUTOCONFIG.N_20\
        );

    \I__701\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5037\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5037\,
            I => \N__5034\
        );

    \I__699\ : Span12Mux_v
    port map (
            O => \N__5034\,
            I => \N__5031\
        );

    \I__698\ : Odrv12
    port map (
            O => \N__5031\,
            I => \CPUCONFn_c\
        );

    \I__697\ : InMux
    port map (
            O => \N__5028\,
            I => \N__5025\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5025\,
            I => \U409_AUTOCONFIG.N_52\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__5022\,
            I => \U409_AUTOCONFIG.N_52_cascade_\
        );

    \I__694\ : InMux
    port map (
            O => \N__5019\,
            I => \N__5011\
        );

    \I__693\ : InMux
    port map (
            O => \N__5018\,
            I => \N__5011\
        );

    \I__692\ : InMux
    port map (
            O => \N__5017\,
            I => \N__5006\
        );

    \I__691\ : InMux
    port map (
            O => \N__5016\,
            I => \N__5006\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5011\,
            I => \U409_AUTOCONFIG.N_56\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5006\,
            I => \U409_AUTOCONFIG.N_56\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__5001\,
            I => \N__4997\
        );

    \I__687\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4994\
        );

    \I__686\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4991\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4994\,
            I => \N__4988\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__4991\,
            I => \N__4985\
        );

    \I__683\ : Odrv12
    port map (
            O => \N__4988\,
            I => \U409_AUTOCONFIG.N_67\
        );

    \I__682\ : Odrv4
    port map (
            O => \N__4985\,
            I => \U409_AUTOCONFIG.N_67\
        );

    \I__681\ : CascadeMux
    port map (
            O => \N__4980\,
            I => \U409_AUTOCONFIG.N_56_cascade_\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__4977\,
            I => \N__4971\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__4976\,
            I => \N__4968\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__4975\,
            I => \N__4965\
        );

    \I__677\ : CascadeMux
    port map (
            O => \N__4974\,
            I => \N__4961\
        );

    \I__676\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4955\
        );

    \I__675\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4950\
        );

    \I__674\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4950\
        );

    \I__673\ : InMux
    port map (
            O => \N__4964\,
            I => \N__4942\
        );

    \I__672\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4942\
        );

    \I__671\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4939\
        );

    \I__670\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4934\
        );

    \I__669\ : InMux
    port map (
            O => \N__4958\,
            I => \N__4934\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4955\,
            I => \N__4929\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4950\,
            I => \N__4929\
        );

    \I__666\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4926\
        );

    \I__665\ : InMux
    port map (
            O => \N__4948\,
            I => \N__4921\
        );

    \I__664\ : InMux
    port map (
            O => \N__4947\,
            I => \N__4921\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4942\,
            I => \N__4918\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__4939\,
            I => \N__4913\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4934\,
            I => \N__4913\
        );

    \I__660\ : Span4Mux_v
    port map (
            O => \N__4929\,
            I => \N__4910\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4926\,
            I => \N__4905\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4921\,
            I => \N__4905\
        );

    \I__657\ : Span4Mux_v
    port map (
            O => \N__4918\,
            I => \N__4901\
        );

    \I__656\ : Span4Mux_v
    port map (
            O => \N__4913\,
            I => \N__4898\
        );

    \I__655\ : Span4Mux_h
    port map (
            O => \N__4910\,
            I => \N__4893\
        );

    \I__654\ : Span4Mux_v
    port map (
            O => \N__4905\,
            I => \N__4893\
        );

    \I__653\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4890\
        );

    \I__652\ : Sp12to4
    port map (
            O => \N__4901\,
            I => \N__4881\
        );

    \I__651\ : Sp12to4
    port map (
            O => \N__4898\,
            I => \N__4881\
        );

    \I__650\ : Sp12to4
    port map (
            O => \N__4893\,
            I => \N__4881\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4890\,
            I => \N__4881\
        );

    \I__648\ : Odrv12
    port map (
            O => \N__4881\,
            I => \A_c_4\
        );

    \I__647\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4875\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4875\,
            I => \N__4868\
        );

    \I__645\ : InMux
    port map (
            O => \N__4874\,
            I => \N__4863\
        );

    \I__644\ : InMux
    port map (
            O => \N__4873\,
            I => \N__4863\
        );

    \I__643\ : CascadeMux
    port map (
            O => \N__4872\,
            I => \N__4859\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__4871\,
            I => \N__4856\
        );

    \I__641\ : Span4Mux_v
    port map (
            O => \N__4868\,
            I => \N__4853\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4863\,
            I => \N__4848\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__4862\,
            I => \N__4845\
        );

    \I__638\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4838\
        );

    \I__637\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4838\
        );

    \I__636\ : Span4Mux_h
    port map (
            O => \N__4853\,
            I => \N__4835\
        );

    \I__635\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4830\
        );

    \I__634\ : InMux
    port map (
            O => \N__4851\,
            I => \N__4830\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__4848\,
            I => \N__4827\
        );

    \I__632\ : InMux
    port map (
            O => \N__4845\,
            I => \N__4820\
        );

    \I__631\ : InMux
    port map (
            O => \N__4844\,
            I => \N__4820\
        );

    \I__630\ : InMux
    port map (
            O => \N__4843\,
            I => \N__4820\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__4838\,
            I => \N__4817\
        );

    \I__628\ : Sp12to4
    port map (
            O => \N__4835\,
            I => \N__4808\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__4830\,
            I => \N__4808\
        );

    \I__626\ : Sp12to4
    port map (
            O => \N__4827\,
            I => \N__4808\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4820\,
            I => \N__4808\
        );

    \I__624\ : Span4Mux_v
    port map (
            O => \N__4817\,
            I => \N__4805\
        );

    \I__623\ : Span12Mux_h
    port map (
            O => \N__4808\,
            I => \N__4802\
        );

    \I__622\ : Span4Mux_h
    port map (
            O => \N__4805\,
            I => \N__4799\
        );

    \I__621\ : Span12Mux_v
    port map (
            O => \N__4802\,
            I => \N__4796\
        );

    \I__620\ : Sp12to4
    port map (
            O => \N__4799\,
            I => \N__4793\
        );

    \I__619\ : Odrv12
    port map (
            O => \N__4796\,
            I => \A_c_2\
        );

    \I__618\ : Odrv12
    port map (
            O => \N__4793\,
            I => \A_c_2\
        );

    \I__617\ : InMux
    port map (
            O => \N__4788\,
            I => \N__4785\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4785\,
            I => \U409_AUTOCONFIG.N_44\
        );

    \I__615\ : InMux
    port map (
            O => \N__4782\,
            I => \N__4779\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4779\,
            I => \N__4775\
        );

    \I__613\ : InMux
    port map (
            O => \N__4778\,
            I => \N__4772\
        );

    \I__612\ : Span4Mux_v
    port map (
            O => \N__4775\,
            I => \N__4765\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__4772\,
            I => \N__4762\
        );

    \I__610\ : InMux
    port map (
            O => \N__4771\,
            I => \N__4757\
        );

    \I__609\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4757\
        );

    \I__608\ : InMux
    port map (
            O => \N__4769\,
            I => \N__4752\
        );

    \I__607\ : InMux
    port map (
            O => \N__4768\,
            I => \N__4752\
        );

    \I__606\ : Odrv4
    port map (
            O => \N__4765\,
            I => \U409_AUTOCONFIG.N_86\
        );

    \I__605\ : Odrv4
    port map (
            O => \N__4762\,
            I => \U409_AUTOCONFIG.N_86\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4757\,
            I => \U409_AUTOCONFIG.N_86\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4752\,
            I => \U409_AUTOCONFIG.N_86\
        );

    \I__602\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4730\
        );

    \I__601\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4730\
        );

    \I__600\ : InMux
    port map (
            O => \N__4741\,
            I => \N__4730\
        );

    \I__599\ : InMux
    port map (
            O => \N__4740\,
            I => \N__4730\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__4739\,
            I => \N__4727\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4730\,
            I => \N__4720\
        );

    \I__596\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4717\
        );

    \I__595\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4712\
        );

    \I__594\ : InMux
    port map (
            O => \N__4725\,
            I => \N__4712\
        );

    \I__593\ : InMux
    port map (
            O => \N__4724\,
            I => \N__4709\
        );

    \I__592\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4706\
        );

    \I__591\ : Span4Mux_v
    port map (
            O => \N__4720\,
            I => \N__4702\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__4717\,
            I => \N__4695\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4712\,
            I => \N__4695\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4709\,
            I => \N__4695\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4706\,
            I => \N__4692\
        );

    \I__586\ : InMux
    port map (
            O => \N__4705\,
            I => \N__4689\
        );

    \I__585\ : Span4Mux_h
    port map (
            O => \N__4702\,
            I => \N__4684\
        );

    \I__584\ : Span4Mux_v
    port map (
            O => \N__4695\,
            I => \N__4684\
        );

    \I__583\ : Span4Mux_h
    port map (
            O => \N__4692\,
            I => \N__4679\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__4689\,
            I => \N__4679\
        );

    \I__581\ : Sp12to4
    port map (
            O => \N__4684\,
            I => \N__4676\
        );

    \I__580\ : Sp12to4
    port map (
            O => \N__4679\,
            I => \N__4673\
        );

    \I__579\ : Span12Mux_s5_h
    port map (
            O => \N__4676\,
            I => \N__4670\
        );

    \I__578\ : Span12Mux_v
    port map (
            O => \N__4673\,
            I => \N__4667\
        );

    \I__577\ : Span12Mux_v
    port map (
            O => \N__4670\,
            I => \N__4664\
        );

    \I__576\ : Odrv12
    port map (
            O => \N__4667\,
            I => \A_c_3\
        );

    \I__575\ : Odrv12
    port map (
            O => \N__4664\,
            I => \A_c_3\
        );

    \I__574\ : InMux
    port map (
            O => \N__4659\,
            I => \N__4656\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4656\,
            I => \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_85_i_i_0\
        );

    \I__572\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4649\
        );

    \I__571\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4646\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4649\,
            I => \N_121\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__4646\,
            I => \N_121\
        );

    \I__568\ : CascadeMux
    port map (
            O => \N__4641\,
            I => \N_121_cascade_\
        );

    \I__567\ : IoInMux
    port map (
            O => \N__4638\,
            I => \N__4635\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4635\,
            I => \N__4631\
        );

    \I__565\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4627\
        );

    \I__564\ : IoSpan4Mux
    port map (
            O => \N__4631\,
            I => \N__4623\
        );

    \I__563\ : InMux
    port map (
            O => \N__4630\,
            I => \N__4620\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4627\,
            I => \N__4617\
        );

    \I__561\ : InMux
    port map (
            O => \N__4626\,
            I => \N__4614\
        );

    \I__560\ : Span4Mux_s0_h
    port map (
            O => \N__4623\,
            I => \N__4611\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4620\,
            I => \N__4608\
        );

    \I__558\ : Span4Mux_v
    port map (
            O => \N__4617\,
            I => \N__4603\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__4614\,
            I => \N__4603\
        );

    \I__556\ : Sp12to4
    port map (
            O => \N__4611\,
            I => \N__4600\
        );

    \I__555\ : Span4Mux_v
    port map (
            O => \N__4608\,
            I => \N__4597\
        );

    \I__554\ : Span4Mux_v
    port map (
            O => \N__4603\,
            I => \N__4594\
        );

    \I__553\ : Span12Mux_v
    port map (
            O => \N__4600\,
            I => \N__4591\
        );

    \I__552\ : Sp12to4
    port map (
            O => \N__4597\,
            I => \N__4588\
        );

    \I__551\ : Span4Mux_v
    port map (
            O => \N__4594\,
            I => \N__4585\
        );

    \I__550\ : Span12Mux_h
    port map (
            O => \N__4591\,
            I => \N__4582\
        );

    \I__549\ : Span12Mux_h
    port map (
            O => \N__4588\,
            I => \N__4579\
        );

    \I__548\ : Span4Mux_v
    port map (
            O => \N__4585\,
            I => \N__4576\
        );

    \I__547\ : Span12Mux_h
    port map (
            O => \N__4582\,
            I => \N__4569\
        );

    \I__546\ : Span12Mux_v
    port map (
            O => \N__4579\,
            I => \N__4569\
        );

    \I__545\ : Sp12to4
    port map (
            O => \N__4576\,
            I => \N__4569\
        );

    \I__544\ : Odrv12
    port map (
            O => \N__4569\,
            I => \A_c_16\
        );

    \I__543\ : InMux
    port map (
            O => \N__4566\,
            I => \N__4563\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4563\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1\
        );

    \I__541\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4557\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4557\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2\
        );

    \I__539\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4551\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4551\,
            I => \N__4548\
        );

    \I__537\ : Span4Mux_v
    port map (
            O => \N__4548\,
            I => \N__4545\
        );

    \I__536\ : Odrv4
    port map (
            O => \N__4545\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_7\
        );

    \I__535\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4538\
        );

    \I__534\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4535\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__4538\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__4535\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\
        );

    \I__531\ : IoInMux
    port map (
            O => \N__4530\,
            I => \N__4527\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4527\,
            I => \N__4524\
        );

    \I__529\ : Span12Mux_s4_v
    port map (
            O => \N__4524\,
            I => \N__4521\
        );

    \I__528\ : Odrv12
    port map (
            O => \N__4521\,
            I => \U409_AUTOCONFIG_D_OUT_0_i_0\
        );

    \I__527\ : InMux
    port map (
            O => \N__4518\,
            I => \N__4515\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4515\,
            I => \N__4512\
        );

    \I__525\ : Span4Mux_v
    port map (
            O => \N__4512\,
            I => \N__4509\
        );

    \I__524\ : Odrv4
    port map (
            O => \N__4509\,
            I => \U409_AUTOCONFIG.N_27\
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__4506\,
            I => \N__4502\
        );

    \I__522\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4497\
        );

    \I__521\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4497\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__4497\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\
        );

    \I__519\ : InMux
    port map (
            O => \N__4494\,
            I => \N__4491\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4491\,
            I => \N__4487\
        );

    \I__517\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4484\
        );

    \I__516\ : Odrv4
    port map (
            O => \N__4487\,
            I => \U409_AUTOCONFIG.N_111\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4484\,
            I => \U409_AUTOCONFIG.N_111\
        );

    \I__514\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4474\
        );

    \I__513\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4471\
        );

    \I__512\ : InMux
    port map (
            O => \N__4477\,
            I => \N__4468\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4474\,
            I => \U409_AUTOCONFIG.N_41\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__4471\,
            I => \U409_AUTOCONFIG.N_41\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4468\,
            I => \U409_AUTOCONFIG.N_41\
        );

    \I__508\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4458\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4458\,
            I => \U409_AUTOCONFIG.N_43\
        );

    \I__506\ : InMux
    port map (
            O => \N__4455\,
            I => \N__4452\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4452\,
            I => \U409_AUTOCONFIG.N_66\
        );

    \I__504\ : CascadeMux
    port map (
            O => \N__4449\,
            I => \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_i_1_cascade_\
        );

    \I__503\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4443\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4443\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_4\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__4440\,
            I => \U409_ADDRESS_DECODE.N_112_cascade_\
        );

    \I__500\ : InMux
    port map (
            O => \N__4437\,
            I => \N__4434\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4434\,
            I => \U409_ADDRESS_DECODE.N_112\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__4431\,
            I => \U409_AUTOCONFIG.N_74_cascade_\
        );

    \I__497\ : InMux
    port map (
            O => \N__4428\,
            I => \N__4425\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__4425\,
            I => \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_i_0\
        );

    \I__495\ : InMux
    port map (
            O => \N__4422\,
            I => \N__4419\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4419\,
            I => \N__4416\
        );

    \I__493\ : Span4Mux_h
    port map (
            O => \N__4416\,
            I => \N__4413\
        );

    \I__492\ : Odrv4
    port map (
            O => \N__4413\,
            I => \N_89_1\
        );

    \I__491\ : CascadeMux
    port map (
            O => \N__4410\,
            I => \N_89_1_cascade_\
        );

    \I__490\ : InMux
    port map (
            O => \N__4407\,
            I => \N__4404\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4404\,
            I => \N__4401\
        );

    \I__488\ : Odrv4
    port map (
            O => \N__4401\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_3\
        );

    \I__487\ : InMux
    port map (
            O => \N__4398\,
            I => \N__4394\
        );

    \I__486\ : InMux
    port map (
            O => \N__4397\,
            I => \N__4391\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4394\,
            I => \N__4388\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4391\,
            I => \N__4385\
        );

    \I__483\ : Span4Mux_v
    port map (
            O => \N__4388\,
            I => \N__4382\
        );

    \I__482\ : Span4Mux_v
    port map (
            O => \N__4385\,
            I => \N__4379\
        );

    \I__481\ : Sp12to4
    port map (
            O => \N__4382\,
            I => \N__4374\
        );

    \I__480\ : Sp12to4
    port map (
            O => \N__4379\,
            I => \N__4374\
        );

    \I__479\ : Odrv12
    port map (
            O => \N__4374\,
            I => \A_c_25\
        );

    \I__478\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4368\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4368\,
            I => \N__4365\
        );

    \I__476\ : Span12Mux_h
    port map (
            O => \N__4365\,
            I => \N__4362\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__4362\,
            I => \TT_c_0\
        );

    \I__474\ : CascadeMux
    port map (
            O => \N__4359\,
            I => \N__4356\
        );

    \I__473\ : InMux
    port map (
            O => \N__4356\,
            I => \N__4353\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4353\,
            I => \N__4350\
        );

    \I__471\ : Span4Mux_h
    port map (
            O => \N__4350\,
            I => \N__4347\
        );

    \I__470\ : Sp12to4
    port map (
            O => \N__4347\,
            I => \N__4344\
        );

    \I__469\ : Odrv12
    port map (
            O => \N__4344\,
            I => \TT_c_1\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__4341\,
            I => \N__4338\
        );

    \I__467\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__465\ : Odrv4
    port map (
            O => \N__4332\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_9\
        );

    \I__464\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4323\
        );

    \I__463\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4323\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4323\,
            I => \U409_AUTOCONFIG.N_38\
        );

    \I__461\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4317\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4317\,
            I => \U409_AUTOCONFIG.N_48\
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__4314\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_1_0_cascade_\
        );

    \I__458\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4305\
        );

    \I__457\ : InMux
    port map (
            O => \N__4310\,
            I => \N__4305\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4305\,
            I => \N__4302\
        );

    \I__455\ : Odrv4
    port map (
            O => \N__4302\,
            I => \U409_AUTOCONFIG.N_62\
        );

    \I__454\ : CascadeMux
    port map (
            O => \N__4299\,
            I => \U409_ADDRESS_DECODE.N_54_cascade_\
        );

    \I__453\ : InMux
    port map (
            O => \N__4296\,
            I => \N__4288\
        );

    \I__452\ : InMux
    port map (
            O => \N__4295\,
            I => \N__4288\
        );

    \I__451\ : InMux
    port map (
            O => \N__4294\,
            I => \N__4283\
        );

    \I__450\ : InMux
    port map (
            O => \N__4293\,
            I => \N__4283\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__4288\,
            I => \N__4280\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4283\,
            I => \N__4275\
        );

    \I__447\ : Span4Mux_v
    port map (
            O => \N__4280\,
            I => \N__4272\
        );

    \I__446\ : InMux
    port map (
            O => \N__4279\,
            I => \N__4269\
        );

    \I__445\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4266\
        );

    \I__444\ : Span4Mux_v
    port map (
            O => \N__4275\,
            I => \N__4263\
        );

    \I__443\ : Sp12to4
    port map (
            O => \N__4272\,
            I => \N__4254\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4269\,
            I => \N__4254\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__4266\,
            I => \N__4254\
        );

    \I__440\ : Sp12to4
    port map (
            O => \N__4263\,
            I => \N__4254\
        );

    \I__439\ : Odrv12
    port map (
            O => \N__4254\,
            I => \A_c_5\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__4251\,
            I => \N__4247\
        );

    \I__437\ : InMux
    port map (
            O => \N__4250\,
            I => \N__4242\
        );

    \I__436\ : InMux
    port map (
            O => \N__4247\,
            I => \N__4242\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4242\,
            I => \N__4238\
        );

    \I__434\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4235\
        );

    \I__433\ : Odrv4
    port map (
            O => \N__4238\,
            I => \U409_AUTOCONFIG.N_92\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4235\,
            I => \U409_AUTOCONFIG.N_92\
        );

    \I__431\ : CascadeMux
    port map (
            O => \N__4230\,
            I => \U409_AUTOCONFIG.N_86_cascade_\
        );

    \I__430\ : InMux
    port map (
            O => \N__4227\,
            I => \N__4224\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4224\,
            I => \U409_AUTOCONFIG.N_57\
        );

    \I__428\ : InMux
    port map (
            O => \N__4221\,
            I => \N__4218\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__4218\,
            I => \N__4215\
        );

    \I__426\ : Span4Mux_v
    port map (
            O => \N__4215\,
            I => \N__4209\
        );

    \I__425\ : InMux
    port map (
            O => \N__4214\,
            I => \N__4202\
        );

    \I__424\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4202\
        );

    \I__423\ : InMux
    port map (
            O => \N__4212\,
            I => \N__4202\
        );

    \I__422\ : Sp12to4
    port map (
            O => \N__4209\,
            I => \N__4197\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__4202\,
            I => \N__4197\
        );

    \I__420\ : Odrv12
    port map (
            O => \N__4197\,
            I => \A_c_7\
        );

    \I__419\ : InMux
    port map (
            O => \N__4194\,
            I => \N__4185\
        );

    \I__418\ : InMux
    port map (
            O => \N__4193\,
            I => \N__4185\
        );

    \I__417\ : InMux
    port map (
            O => \N__4192\,
            I => \N__4185\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__4185\,
            I => \N__4181\
        );

    \I__415\ : CascadeMux
    port map (
            O => \N__4184\,
            I => \N__4178\
        );

    \I__414\ : Span4Mux_v
    port map (
            O => \N__4181\,
            I => \N__4175\
        );

    \I__413\ : InMux
    port map (
            O => \N__4178\,
            I => \N__4172\
        );

    \I__412\ : Sp12to4
    port map (
            O => \N__4175\,
            I => \N__4167\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__4172\,
            I => \N__4167\
        );

    \I__410\ : Odrv12
    port map (
            O => \N__4167\,
            I => \A_c_6\
        );

    \I__409\ : CascadeMux
    port map (
            O => \N__4164\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4_cascade_\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__4161\,
            I => \N__4157\
        );

    \I__407\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4154\
        );

    \I__406\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4151\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__4154\,
            I => \N__4146\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__4151\,
            I => \N__4146\
        );

    \I__403\ : Sp12to4
    port map (
            O => \N__4146\,
            I => \N__4143\
        );

    \I__402\ : Span12Mux_v
    port map (
            O => \N__4143\,
            I => \N__4140\
        );

    \I__401\ : Odrv12
    port map (
            O => \N__4140\,
            I => \A_c_24\
        );

    \I__400\ : InMux
    port map (
            O => \N__4137\,
            I => \N__4131\
        );

    \I__399\ : InMux
    port map (
            O => \N__4136\,
            I => \N__4131\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__4131\,
            I => \N__4128\
        );

    \I__397\ : Sp12to4
    port map (
            O => \N__4128\,
            I => \N__4125\
        );

    \I__396\ : Span12Mux_v
    port map (
            O => \N__4125\,
            I => \N__4122\
        );

    \I__395\ : Odrv12
    port map (
            O => \N__4122\,
            I => \A_c_26\
        );

    \I__394\ : InMux
    port map (
            O => \N__4119\,
            I => \N__4113\
        );

    \I__393\ : InMux
    port map (
            O => \N__4118\,
            I => \N__4113\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__4113\,
            I => \N__4110\
        );

    \I__391\ : Span4Mux_v
    port map (
            O => \N__4110\,
            I => \N__4107\
        );

    \I__390\ : Sp12to4
    port map (
            O => \N__4107\,
            I => \N__4104\
        );

    \I__389\ : Odrv12
    port map (
            O => \N__4104\,
            I => \A_c_27\
        );

    \I__388\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4098\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__4098\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_5\
        );

    \I__386\ : InMux
    port map (
            O => \N__4095\,
            I => \N__4092\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__4092\,
            I => \N__4089\
        );

    \I__384\ : Odrv4
    port map (
            O => \N__4089\,
            I => \U409_AUTOCONFIG.N_42\
        );

    \I__383\ : CascadeMux
    port map (
            O => \N__4086\,
            I => \U409_AUTOCONFIG.N_111_cascade_\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__4083\,
            I => \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_a3_0Z0Z_2_cascade_\
        );

    \I__381\ : IoInMux
    port map (
            O => \N__4080\,
            I => \N__4077\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__4077\,
            I => \N__4074\
        );

    \I__379\ : IoSpan4Mux
    port map (
            O => \N__4074\,
            I => \N__4071\
        );

    \I__378\ : Span4Mux_s3_h
    port map (
            O => \N__4071\,
            I => \N__4068\
        );

    \I__377\ : Sp12to4
    port map (
            O => \N__4068\,
            I => \N__4065\
        );

    \I__376\ : Span12Mux_h
    port map (
            O => \N__4065\,
            I => \N__4062\
        );

    \I__375\ : Span12Mux_h
    port map (
            O => \N__4062\,
            I => \N__4059\
        );

    \I__374\ : Odrv12
    port map (
            O => \N__4059\,
            I => \A_c_15\
        );

    \I__373\ : IoInMux
    port map (
            O => \N__4056\,
            I => \N__4053\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__4053\,
            I => \N__4050\
        );

    \I__371\ : Span4Mux_s3_h
    port map (
            O => \N__4050\,
            I => \N__4047\
        );

    \I__370\ : Span4Mux_v
    port map (
            O => \N__4047\,
            I => \N__4044\
        );

    \I__369\ : Sp12to4
    port map (
            O => \N__4044\,
            I => \N__4041\
        );

    \I__368\ : Span12Mux_h
    port map (
            O => \N__4041\,
            I => \N__4038\
        );

    \I__367\ : Span12Mux_h
    port map (
            O => \N__4038\,
            I => \N__4035\
        );

    \I__366\ : Odrv12
    port map (
            O => \N__4035\,
            I => \A_c_14\
        );

    \I__365\ : ClkMux
    port map (
            O => \N__4032\,
            I => \N__3990\
        );

    \I__364\ : ClkMux
    port map (
            O => \N__4031\,
            I => \N__3990\
        );

    \I__363\ : ClkMux
    port map (
            O => \N__4030\,
            I => \N__3990\
        );

    \I__362\ : ClkMux
    port map (
            O => \N__4029\,
            I => \N__3990\
        );

    \I__361\ : ClkMux
    port map (
            O => \N__4028\,
            I => \N__3990\
        );

    \I__360\ : ClkMux
    port map (
            O => \N__4027\,
            I => \N__3990\
        );

    \I__359\ : ClkMux
    port map (
            O => \N__4026\,
            I => \N__3990\
        );

    \I__358\ : ClkMux
    port map (
            O => \N__4025\,
            I => \N__3990\
        );

    \I__357\ : ClkMux
    port map (
            O => \N__4024\,
            I => \N__3990\
        );

    \I__356\ : ClkMux
    port map (
            O => \N__4023\,
            I => \N__3990\
        );

    \I__355\ : ClkMux
    port map (
            O => \N__4022\,
            I => \N__3990\
        );

    \I__354\ : ClkMux
    port map (
            O => \N__4021\,
            I => \N__3990\
        );

    \I__353\ : ClkMux
    port map (
            O => \N__4020\,
            I => \N__3990\
        );

    \I__352\ : ClkMux
    port map (
            O => \N__4019\,
            I => \N__3990\
        );

    \I__351\ : GlobalMux
    port map (
            O => \N__3990\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            I => \N__4029\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            I => \N__4021\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            I => \N__4026\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            I => \N__4024\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            I => \N__4022\
        );

    \INVU409_TRANSFER_ACK.CIA_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            I => \N__4020\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__4019\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            I => \N__4027\
        );

    \INVU409_TRANSFER_ACK.TACK_OUTnC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            I => \N__4025\
        );

    \INVU409_TRANSFER_ACK.TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            I => \N__4023\
        );

    \INVU409_TRANSFER_ACK.ROMENn_nessC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROMENn_nessC_net\,
            I => \N__4032\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            I => \N__4028\
        );

    \INVU409_AUTOCONFIG.ATA_BASE_2C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.ATA_BASE_2C_net\,
            I => \N__8262\
        );

    \INVU409_AUTOCONFIG.ATA_BASE_4C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.ATA_BASE_4C_net\,
            I => \N__8263\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            I => \N__4031\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            I => \N__4030\
        );

    \INVU409_AUTOCONFIG.CONFIGENnC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            I => \N__8267\
        );

    \INVU409_AUTOCONFIG.LIDE_CONFC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            I => \N__8266\
        );

    \INVU409_AUTOCONFIG.BRIDGE_OUT_1C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net\,
            I => \N__8268\
        );

    \INVU409_AUTOCONFIG.BRIDGE_OUT_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            I => \N__8270\
        );

    \INVU409_AUTOCONFIG.LIDE_OUT_3C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_OUT_3C_net\,
            I => \N__8269\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_16_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_7_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8169\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_4_0_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4192\,
            in1 => \N__4212\,
            in2 => \_gnd_net_\,
            in3 => \N__4725\,
            lcout => \U409_AUTOCONFIG.N_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_11_3_i_o3_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4214\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4194\,
            lcout => \U409_AUTOCONFIG.N_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_a3_0_2_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__4726\,
            in1 => \N__6342\,
            in2 => \N__4872\,
            in3 => \N__4948\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_a3_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0_0_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__4294\,
            in1 => \N__4949\,
            in2 => \N__4083\,
            in3 => \N__10187\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4241\,
            in1 => \N__4293\,
            in2 => \N__4871\,
            in3 => \N__4947\,
            lcout => \U409_AUTOCONFIG.N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_1_sqmuxa_0_a2_0_2_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4193\,
            in1 => \N__4782\,
            in2 => \N__4739\,
            in3 => \N__4213\,
            lcout => \U409_AUTOCONFIG.LIDE_CONF_1_sqmuxa_0_a2_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_5_0_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__4221\,
            in1 => \N__6341\,
            in2 => \N__4184\,
            in3 => \N__4724\,
            lcout => \U409_AUTOCONFIG.N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7027\,
            in1 => \N__5852\,
            in2 => \_gnd_net_\,
            in3 => \N__4160\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_3_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__4397\,
            in1 => \N__10191\,
            in2 => \N__4164\,
            in3 => \N__4101\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_7_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4119\,
            in1 => \N__4422\,
            in2 => \N__4161\,
            in3 => \N__4137\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_5_LC_3_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4136\,
            in1 => \N__5980\,
            in2 => \N__5903\,
            in3 => \N__4118\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_4_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__6114\,
            in1 => \N__5610\,
            in2 => \N__6032\,
            in3 => \N__4626\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_o2_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100110011"
        )
    port map (
            in0 => \N__6359\,
            in1 => \N__10148\,
            in2 => \N__5001\,
            in3 => \N__4769\,
            lcout => \U409_AUTOCONFIG.N_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_6_0_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4873\,
            in1 => \N__4311\,
            in2 => \_gnd_net_\,
            in3 => \N__4295\,
            lcout => \U409_AUTOCONFIG.N_111\,
            ltout => \U409_AUTOCONFIG.N_111_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__6358\,
            in1 => \N__4095\,
            in2 => \N__4086\,
            in3 => \N__4960\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__4768\,
            in1 => \N__4477\,
            in2 => \N__4314\,
            in3 => \N__4310\,
            lcout => \U409_AUTOCONFIG.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_3_1_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__4296\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4874\,
            lcout => \U409_AUTOCONFIG.N_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_2_i_o3_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6481\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7150\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.N_54_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6115\,
            in1 => \N__6924\,
            in2 => \N__4299\,
            in3 => \N__6574\,
            lcout => \U409_ADDRESS_DECODE.HIROMZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__4705\,
            in1 => \N__6352\,
            in2 => \N__4862\,
            in3 => \N__4959\,
            lcout => \U409_AUTOCONFIG.N_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__4478\,
            in1 => \N__4278\,
            in2 => \N__4251\,
            in3 => \N__4843\,
            lcout => \U409_AUTOCONFIG.N_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_0_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4844\,
            in1 => \N__4279\,
            in2 => \_gnd_net_\,
            in3 => \N__4958\,
            lcout => \U409_AUTOCONFIG.N_86\,
            ltout => \U409_AUTOCONFIG.N_86_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110011"
        )
    port map (
            in0 => \N__4250\,
            in1 => \N__10149\,
            in2 => \N__4230\,
            in3 => \N__4227\,
            lcout => \U409_AUTOCONFIG.N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_3_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4494\,
            in1 => \N__6351\,
            in2 => \_gnd_net_\,
            in3 => \N__4904\,
            lcout => \U409_AUTOCONFIG.N_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_3_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6480\,
            in1 => \N__4652\,
            in2 => \N__7166\,
            in3 => \N__4634\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_1_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6573\,
            in2 => \_gnd_net_\,
            in3 => \N__6925\,
            lcout => \N_89_1\,
            ltout => \N_89_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4653\,
            in1 => \N__6479\,
            in2 => \N__4410\,
            in3 => \N__7146\,
            lcout => \U409_ADDRESS_DECODE.N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_11_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4407\,
            in1 => \N__10176\,
            in2 => \N__4341\,
            in3 => \N__4398\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_9_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5902\,
            in1 => \N__4371\,
            in2 => \N__4359\,
            in3 => \N__5981\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_0_3_163_i_i_o2_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__4778\,
            in1 => \N__10169\,
            in2 => \_gnd_net_\,
            in3 => \N__6372\,
            lcout => \U409_AUTOCONFIG.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__4329\,
            in1 => \N__4461\,
            in2 => \N__5193\,
            in3 => \N__5234\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000010001"
        )
    port map (
            in0 => \N__4788\,
            in1 => \N__4328\,
            in2 => \N__5285\,
            in3 => \N__5188\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__4320\,
            in1 => \N__4659\,
            in2 => \N__5192\,
            in3 => \N__4541\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001000"
        )
    port map (
            in0 => \N__6353\,
            in1 => \N__4490\,
            in2 => \N__4974\,
            in3 => \N__4479\,
            lcout => \U409_AUTOCONFIG.N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4964\,
            in1 => \N__4878\,
            in2 => \N__6379\,
            in3 => \N__4723\,
            lcout => \U409_AUTOCONFIG.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110101010101"
        )
    port map (
            in0 => \N__10170\,
            in1 => \N__4455\,
            in2 => \N__4977\,
            in3 => \N__6357\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000101"
        )
    port map (
            in0 => \N__4428\,
            in1 => \N__5345\,
            in2 => \N__4449\,
            in3 => \N__5184\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a2_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6907\,
            in1 => \N__6487\,
            in2 => \_gnd_net_\,
            in3 => \N__7161\,
            lcout => \U409_ADDRESS_DECODE.N_112\,
            ltout => \U409_ADDRESS_DECODE.N_112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7189\,
            in1 => \N__4446\,
            in2 => \N__4440\,
            in3 => \N__6580\,
            lcout => \AUTOCONFIG_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3_0_2_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__6045\,
            in1 => \N__4437\,
            in2 => \_gnd_net_\,
            in3 => \N__6131\,
            lcout => \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4743\,
            in1 => \N__6362\,
            in2 => \N__4976\,
            in3 => \N__4852\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.N_74_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__6360\,
            in1 => \N__4770\,
            in2 => \N__4431\,
            in3 => \N__4740\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_0_114_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__4741\,
            in1 => \N__6361\,
            in2 => \N__4975\,
            in3 => \N__4851\,
            lcout => \U409_AUTOCONFIG.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__10147\,
            in1 => \N__4771\,
            in2 => \_gnd_net_\,
            in3 => \N__4742\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_cnst_0_a2_1_85_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un2_REGSPACEn_i_a2_0_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6046\,
            in1 => \N__6133\,
            in2 => \_gnd_net_\,
            in3 => \N__5617\,
            lcout => \N_121\,
            ltout => \N_121_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__6893\,
            in1 => \_gnd_net_\,
            in2 => \N__4641\,
            in3 => \N__4630\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4566\,
            in1 => \N__4560\,
            in2 => \N__5478\,
            in3 => \N__6485\,
            lcout => \CIA_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_2_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7159\,
            in1 => \N__5734\,
            in2 => \N__5665\,
            in3 => \N__6575\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13_10_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7032\,
            in1 => \N__4554\,
            in2 => \_gnd_net_\,
            in3 => \N__5845\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_13Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIA2DB1_0_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__4542\,
            in1 => \N__4505\,
            in2 => \N__6230\,
            in3 => \N__5710\,
            lcout => \U409_AUTOCONFIG_D_OUT_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000101010101"
        )
    port map (
            in0 => \N__4518\,
            in1 => \N__10153\,
            in2 => \N__4506\,
            in3 => \N__5018\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001100010011"
        )
    port map (
            in0 => \N__5019\,
            in1 => \N__5082\,
            in2 => \N__10177\,
            in3 => \N__5255\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000101010101"
        )
    port map (
            in0 => \N__5070\,
            in1 => \N__10160\,
            in2 => \N__5333\,
            in3 => \N__5016\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_0_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000011110000"
        )
    port map (
            in0 => \N__5791\,
            in1 => \N__5770\,
            in2 => \N__10180\,
            in3 => \N__5028\,
            lcout => \U409_AUTOCONFIG.STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5769\,
            in1 => \N__5058\,
            in2 => \_gnd_net_\,
            in3 => \N__5790\,
            lcout => \U409_AUTOCONFIG.N_122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001100010011"
        )
    port map (
            in0 => \N__5017\,
            in1 => \N__5049\,
            in2 => \N__10179\,
            in3 => \N__5303\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000001000"
        )
    port map (
            in0 => \N__5771\,
            in1 => \N__10167\,
            in2 => \N__5549\,
            in3 => \N__5792\,
            lcout => \U409_AUTOCONFIG.STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_ns_1_0__m2_0_o2_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__5040\,
            in1 => \N__5768\,
            in2 => \_gnd_net_\,
            in3 => \N__5118\,
            lcout => \U409_AUTOCONFIG.N_52\,
            ltout => \U409_AUTOCONFIG.N_52_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIBM2Q1_1_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__5543\,
            in1 => \_gnd_net_\,
            in2 => \N__5022\,
            in3 => \N__5789\,
            lcout => \U409_AUTOCONFIG.N_56\,
            ltout => \U409_AUTOCONFIG.N_56_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNI7U5N3_1_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__10168\,
            in1 => \N__5000\,
            in2 => \N__4980\,
            in3 => \N__5202\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_7_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.LOWROM_2_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7162\,
            in1 => \N__6584\,
            in2 => \N__6492\,
            in3 => \N__6923\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.LOWROMZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_ROMEN_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__5172\,
            in1 => \N__7077\,
            in2 => \N__5163\,
            in3 => \N__6132\,
            lcout => \U409_ADDRESS_DECODE_un1_ROMEN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.D_1_i_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5539\,
            in1 => \N__10268\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \D_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__10269\,
            in1 => \N__8349\,
            in2 => \_gnd_net_\,
            in3 => \N__5703\,
            lcout => \U409_AUTOCONFIG.AC_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_1_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5667\,
            in1 => \N__5750\,
            in2 => \N__6590\,
            in3 => \N__5625\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_4_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6134\,
            in1 => \N__6486\,
            in2 => \N__5112\,
            in3 => \N__6047\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_4\,
            ltout => \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5472\,
            in1 => \N__6906\,
            in2 => \N__5109\,
            in3 => \N__7160\,
            lcout => \N_120\,
            ltout => \N_120_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__5106\,
            in1 => \_gnd_net_\,
            in2 => \N__5097\,
            in3 => \N__5094\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_1_0_a2_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__5749\,
            in1 => \N__5666\,
            in2 => \_gnd_net_\,
            in3 => \N__5471\,
            lcout => \U409_ADDRESS_DECODE_ROMEN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111111111"
        )
    port map (
            in0 => \N__5364\,
            in1 => \N__5376\,
            in2 => \N__6589\,
            in3 => \N__5470\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100000"
        )
    port map (
            in0 => \N__5375\,
            in1 => \N__5363\,
            in2 => \N__5479\,
            in3 => \N__6576\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIC4DB1_1_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__5352\,
            in1 => \N__5334\,
            in2 => \N__6231\,
            in3 => \N__5712\,
            lcout => \U409_AUTOCONFIG_D_OUT_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIE6DB1_2_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__5304\,
            in1 => \N__5705\,
            in2 => \N__5292\,
            in3 => \N__6211\,
            lcout => \U409_AUTOCONFIG_D_OUT_0_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6383\,
            in1 => \N__6210\,
            in2 => \_gnd_net_\,
            in3 => \N__6163\,
            lcout => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIG8DB1_3_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__5256\,
            in1 => \N__5706\,
            in2 => \N__5244\,
            in3 => \N__6212\,
            lcout => \U409_AUTOCONFIG_D_OUT_0_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__6215\,
            in1 => \N__6371\,
            in2 => \_gnd_net_\,
            in3 => \N__6166\,
            lcout => \U409_AUTOCONFIG.LIDE_CONFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__9028\
        );

    \U409_AUTOCONFIG.CONFIGURED_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__6167\,
            in1 => \N__6216\,
            in2 => \N__6382\,
            in3 => \N__5704\,
            lcout => \CONFIGURED\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__9028\
        );

    \U409_AUTOCONFIG.AC_TACK_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001000"
        )
    port map (
            in0 => \N__5793\,
            in1 => \N__5772\,
            in2 => \N__5550\,
            in3 => \N__7544\,
            lcout => \AC_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__9028\
        );

    \U409_AUTOCONFIG.ATA_BASE_3_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7326\,
            in1 => \N__7292\,
            in2 => \N__6708\,
            in3 => \N__6063\,
            lcout => \ATA_BASE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__9028\
        );

    \U409_AUTOCONFIG.ATA_BASE_1_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7325\,
            in1 => \N__7291\,
            in2 => \N__7432\,
            in3 => \N__5568\,
            lcout => \ATA_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__9028\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__5751\,
            in1 => \_gnd_net_\,
            in2 => \N__5711\,
            in3 => \N__5656\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1\,
            ltout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__5624\,
            in1 => \N__5480\,
            in2 => \N__5571\,
            in3 => \N__5567\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6390\,
            in1 => \N__5994\,
            in2 => \N__5556\,
            in3 => \N__6846\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0\,
            ltout => \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001000000"
        )
    port map (
            in0 => \N__5544\,
            in1 => \N__10178\,
            in2 => \N__5553\,
            in3 => \N__6805\,
            lcout => \U409_ADDRESS_DECODE.ATA_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_0_a3_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__10279\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5545\,
            lcout => \un1_AUTOCONFIG_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.N_120_i_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__5490\,
            in1 => \N__7167\,
            in2 => \N__5484\,
            in3 => \N__6932\,
            lcout => \N_120_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_1_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7624\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7913\,
            lcout => \U409_TRANSFER_ACK.CO1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_3_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000000000"
        )
    port map (
            in0 => \N__6663\,
            in1 => \N__5988\,
            in2 => \N__5982\,
            in3 => \N__5820\,
            lcout => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_1_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7599\,
            in1 => \N__7622\,
            in2 => \N__7921\,
            in3 => \N__7865\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.LOWROM_3_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__6588\,
            in1 => \N__6491\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_ADDRESS_DECODE.LOWROMZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__7623\,
            in1 => \N__7598\,
            in2 => \N__7876\,
            in3 => \N__7909\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10231\,
            in1 => \N__10288\,
            in2 => \_gnd_net_\,
            in3 => \N__5937\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.PORTSIZEZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNI4345U_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111001111"
        )
    port map (
            in0 => \N__7760\,
            in1 => \N__7724\,
            in2 => \N__5931\,
            in3 => \N__6810\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_0_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__6648\,
            in1 => \N__5907\,
            in2 => \N__5862\,
            in3 => \N__6627\,
            lcout => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.CONFIGENn_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000101010101010"
        )
    port map (
            in0 => \N__5804\,
            in1 => \N__6384\,
            in2 => \N__6226\,
            in3 => \N__6171\,
            lcout => \CONFIGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            ce => 'H',
            sr => \N__9029\
        );

    \U409_AUTOCONFIG.ATA_BASE_7_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7346\,
            in1 => \N__7386\,
            in2 => \N__6697\,
            in3 => \N__6504\,
            lcout => \ATA_BASE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            ce => 'H',
            sr => \N__9029\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7352\,
            in1 => \N__6609\,
            in2 => \N__6698\,
            in3 => \N__6659\,
            lcout => \BRIDGE_BASE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            ce => 'H',
            sr => \N__9029\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__7264\,
            in1 => \N__7351\,
            in2 => \N__6644\,
            in3 => \N__6608\,
            lcout => \BRIDGE_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            ce => 'H',
            sr => \N__9029\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__6606\,
            in1 => \N__7439\,
            in2 => \N__7356\,
            in3 => \N__6620\,
            lcout => \BRIDGE_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            ce => 'H',
            sr => \N__9029\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__7484\,
            in1 => \N__7347\,
            in2 => \N__6986\,
            in3 => \N__6607\,
            lcout => \BRIDGE_BASE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            ce => 'H',
            sr => \N__9029\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__6591\,
            in1 => \N__6503\,
            in2 => \N__6478\,
            in3 => \N__7367\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_1_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6381\,
            in1 => \N__6214\,
            in2 => \_gnd_net_\,
            in3 => \N__6165\,
            lcout => \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6380\,
            in1 => \N__6213\,
            in2 => \_gnd_net_\,
            in3 => \N__6164\,
            lcout => \U409_AUTOCONFIG.LIDE_CONF_RNIUPP42Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__6135\,
            in1 => \N__6062\,
            in2 => \N__6051\,
            in3 => \N__7232\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_1_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__7168\,
            in1 => \N__7397\,
            in2 => \N__6936\,
            in3 => \N__7460\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACE_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__7202\,
            in1 => \N__7066\,
            in2 => \N__7221\,
            in3 => \N__7169\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6819\,
            in1 => \N__8367\,
            in2 => \N__8306\,
            in3 => \N__7203\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNI206O6_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__7753\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6806\,
            lcout => \U409_ADDRESS_DECODE_un1_ATA_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__7601\,
            in1 => \N__6768\,
            in2 => \N__6720\,
            in3 => \N__7869\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__9023\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__6767\,
            in1 => \N__6716\,
            in2 => \_gnd_net_\,
            in3 => \N__7602\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__9023\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7914\,
            in2 => \_gnd_net_\,
            in3 => \N__7626\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__9023\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000101"
        )
    port map (
            in0 => \N__7925\,
            in1 => \N__6747\,
            in2 => \N__6735\,
            in3 => \N__6759\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__9019\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIL9Q68_1_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6758\,
            in1 => \N__6746\,
            in2 => \_gnd_net_\,
            in3 => \N__6731\,
            lcout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0\,
            ltout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_ness_RNO_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9033\,
            in1 => \_gnd_net_\,
            in2 => \N__7497\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.ATA_BASE_4_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7353\,
            in1 => \N__7383\,
            in2 => \N__7494\,
            in3 => \N__7461\,
            lcout => \ATA_BASE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_4C_net\,
            ce => 'H',
            sr => \N__9026\
        );

    \U409_AUTOCONFIG.ATA_BASE_5_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7354\,
            in1 => \N__7384\,
            in2 => \N__7449\,
            in3 => \N__7398\,
            lcout => \ATA_BASE_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_4C_net\,
            ce => 'H',
            sr => \N__9026\
        );

    \U409_AUTOCONFIG.ATA_BASE_6_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7355\,
            in1 => \N__7385\,
            in2 => \N__7277\,
            in3 => \N__7368\,
            lcout => \ATA_BASE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_4C_net\,
            ce => 'H',
            sr => \N__9026\
        );

    \U409_AUTOCONFIG.ATA_BASE_2_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7338\,
            in1 => \N__7293\,
            in2 => \N__7278\,
            in3 => \N__7233\,
            lcout => \ATA_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_2C_net\,
            ce => 'H',
            sr => \N__9024\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__7220\,
            in1 => \N__7196\,
            in2 => \N__7173\,
            in3 => \N__7073\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8303\,
            in1 => \N__8368\,
            in2 => \N__7817\,
            in3 => \N__7829\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111111111"
        )
    port map (
            in0 => \N__7031\,
            in1 => \N__10080\,
            in2 => \N__6990\,
            in3 => \N__6969\,
            lcout => \U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7625\,
            in2 => \_gnd_net_\,
            in3 => \N__7600\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_ness_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7878\,
            lcout => \ROMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROMENn_nessC_net\,
            ce => \N__7560\,
            sr => \N__9016\
        );

    \U409_TRANSFER_ACK.TACK_EN_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000001110001"
        )
    port map (
            in0 => \N__7515\,
            in1 => \N__8004\,
            in2 => \N__10324\,
            in3 => \N__7527\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            ce => 'H',
            sr => \N__9025\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__7946\,
            in1 => \_gnd_net_\,
            in2 => \N__10146\,
            in3 => \N__7932\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__8002\,
            in1 => \_gnd_net_\,
            in2 => \N__10145\,
            in3 => \N__7513\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001010000"
        )
    port map (
            in0 => \N__8003\,
            in1 => \N__7514\,
            in2 => \N__10144\,
            in3 => \N__7526\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8153\,
            in2 => \_gnd_net_\,
            in3 => \N__7793\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7548\,
            in1 => \N__7841\,
            in2 => \N__7530\,
            in3 => \N__8015\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER6\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111011101"
        )
    port map (
            in0 => \N__7512\,
            in1 => \N__8001\,
            in2 => \N__7986\,
            in3 => \N__7945\,
            lcout => \U409_TRANSFER_ACK.TACK_OUTn_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__7842\,
            in1 => \N__7926\,
            in2 => \N__7887\,
            in3 => \N__7877\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9017\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__7689\,
            in1 => \N__7830\,
            in2 => \N__7818\,
            in3 => \N__7794\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9017\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__7782\,
            in1 => \N__10094\,
            in2 => \N__7737\,
            in3 => \N__7713\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.LV_SPACE_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7764\,
            in1 => \N__10295\,
            in2 => \N__7736\,
            in3 => \N__7712\,
            lcout => \BUFENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8369\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8301\,
            lcout => \U409_TRANSFER_ACK.N_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8305\,
            lcout => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8585\,
            in2 => \_gnd_net_\,
            in3 => \N__8421\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9606\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__9369\,
            in1 => \N__8385\,
            in2 => \N__9336\,
            in3 => \N__9399\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9608\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__8519\,
            in1 => \_gnd_net_\,
            in2 => \N__8562\,
            in3 => \N__8304\,
            lcout => \U409_TRANSFER_ACK.N_17_mux\,
            ltout => \U409_TRANSFER_ACK.N_17_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100111111"
        )
    port map (
            in0 => \N__8536\,
            in1 => \N__8057\,
            in2 => \N__8091\,
            in3 => \N__8548\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010010001100"
        )
    port map (
            in0 => \N__8033\,
            in1 => \N__10061\,
            in2 => \N__8088\,
            in3 => \N__8082\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011111"
        )
    port map (
            in0 => \N__8549\,
            in1 => \N__8537\,
            in2 => \N__8066\,
            in3 => \N__8076\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.N_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101000001000"
        )
    port map (
            in0 => \N__10062\,
            in1 => \N__8032\,
            in2 => \N__8085\,
            in3 => \N__8064\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__8550\,
            in1 => \N__8535\,
            in2 => \N__8067\,
            in3 => \N__8075\,
            lcout => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8558\,
            in2 => \_gnd_net_\,
            in3 => \N__8518\,
            lcout => \U409_TRANSFER_ACK.N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111100001000"
        )
    port map (
            in0 => \N__8065\,
            in1 => \N__8040\,
            in2 => \N__8034\,
            in3 => \N__8016\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9018\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__8205\,
            in1 => \N__8154\,
            in2 => \_gnd_net_\,
            in3 => \N__8118\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            ce => 'H',
            sr => \N__8773\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8964\,
            in1 => \N__8945\,
            in2 => \N__8192\,
            in3 => \N__8101\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8924\,
            in2 => \_gnd_net_\,
            in3 => \N__8865\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__8965\,
            in1 => \N__8946\,
            in2 => \N__8193\,
            in3 => \N__8102\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__8893\,
            in1 => \N__8798\,
            in2 => \N__8142\,
            in3 => \N__8135\,
            lcout => \U409_TRANSFER_ACK.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8797\,
            in1 => \N__8892\,
            in2 => \N__8139\,
            in3 => \N__8127\,
            lcout => \U409_TRANSFER_ACK.N_87\,
            ltout => \U409_TRANSFER_ACK.N_87_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011111111"
        )
    port map (
            in0 => \N__8370\,
            in1 => \N__8302\,
            in2 => \N__8121\,
            in3 => \N__8117\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__8190\,
            in1 => \N__8103\,
            in2 => \N__8106\,
            in3 => \N__8982\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7C_net\,
            ce => 'H',
            sr => \N__8777\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__8928\,
            in1 => \N__8899\,
            in2 => \_gnd_net_\,
            in3 => \N__8832\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__8766\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8927\,
            in2 => \N__8904\,
            in3 => \N__8868\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__8766\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110000110011"
        )
    port map (
            in0 => \N__8348\,
            in1 => \N__8898\,
            in2 => \N__8307\,
            in3 => \N__8204\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__8766\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__8981\,
            in1 => \N__8191\,
            in2 => \_gnd_net_\,
            in3 => \N__8831\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__8766\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10027\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9736\,
            in1 => \N__9783\,
            in2 => \N__9690\,
            in3 => \N__9069\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9054\,
            in1 => \N__8729\,
            in2 => \N__9093\,
            in3 => \N__9227\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__9735\,
            in1 => \N__9686\,
            in2 => \N__9128\,
            in3 => \N__9784\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8419\,
            in2 => \N__8589\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8447\,
            in2 => \_gnd_net_\,
            in3 => \N__8157\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__9600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8603\,
            in2 => \_gnd_net_\,
            in3 => \N__8403\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__9600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8643\,
            in2 => \_gnd_net_\,
            in3 => \N__8400\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8654\,
            in2 => \_gnd_net_\,
            in3 => \N__8397\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__9600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9507\,
            in2 => \_gnd_net_\,
            in3 => \N__8394\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8708\,
            in2 => \_gnd_net_\,
            in3 => \N__8391\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__9600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9416\,
            in2 => \_gnd_net_\,
            in3 => \N__8388\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9518\,
            in2 => \_gnd_net_\,
            in3 => \N__8379\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8696\,
            in2 => \_gnd_net_\,
            in3 => \N__8376\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__9602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8621\,
            in2 => \_gnd_net_\,
            in3 => \N__8373\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__9602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8462\,
            in2 => \_gnd_net_\,
            in3 => \N__8505\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__9602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8681\,
            in2 => \_gnd_net_\,
            in3 => \N__8502\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__9602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9482\,
            in2 => \_gnd_net_\,
            in3 => \N__8499\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8669\,
            in2 => \_gnd_net_\,
            in3 => \N__8496\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8435\,
            in2 => \_gnd_net_\,
            in3 => \N__8493\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9395\,
            in1 => \N__9365\,
            in2 => \N__9334\,
            in3 => \N__8490\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__9363\,
            in1 => \N__9393\,
            in2 => \N__8481\,
            in3 => \N__9325\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9394\,
            in1 => \N__9364\,
            in2 => \N__9333\,
            in3 => \N__8472\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8463\,
            in1 => \N__8451\,
            in2 => \N__8436\,
            in3 => \N__8420\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8712\,
            in1 => \N__8697\,
            in2 => \N__8685\,
            in3 => \N__8670\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__8658\,
            in1 => \N__8642\,
            in2 => \_gnd_net_\,
            in3 => \N__8583\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8628\,
            in1 => \N__8622\,
            in2 => \N__8610\,
            in3 => \N__8607\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__9362\,
            in1 => \N__9318\,
            in2 => \N__8592\,
            in3 => \N__8584\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8520\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \N__9027\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8538\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \N__9027\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10060\,
            in2 => \_gnd_net_\,
            in3 => \N__9974\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \N__9027\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9200\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \N__9027\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8966\,
            in1 => \N__8866\,
            in2 => \N__8805\,
            in3 => \N__8947\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8894\,
            in2 => \N__8985\,
            in3 => \N__8925\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8948\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8802\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__8967\,
            in1 => \N__8834\,
            in2 => \N__8970\,
            in3 => \N__8846\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__8778\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__8949\,
            in1 => \N__8804\,
            in2 => \N__8847\,
            in3 => \N__8833\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__8778\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__8926\,
            in1 => \_gnd_net_\,
            in2 => \N__8903\,
            in3 => \N__8867\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010000010100"
        )
    port map (
            in0 => \N__8835\,
            in1 => \N__8803\,
            in2 => \N__8808\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__8778\
        );

    \U409_TICK.COUNTER50_1_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9120\,
            in2 => \_gnd_net_\,
            in3 => \N__8730\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9599\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8728\,
            in2 => \N__9124\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9089\,
            in2 => \_gnd_net_\,
            in3 => \N__9078\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__9601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9140\,
            in2 => \_gnd_net_\,
            in3 => \N__9075\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__9601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9851\,
            in2 => \_gnd_net_\,
            in3 => \N__9072\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__9601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9164\,
            in3 => \N__9063\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9878\,
            in2 => \_gnd_net_\,
            in3 => \N__9060\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9866\,
            in2 => \_gnd_net_\,
            in3 => \N__9057\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__9601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9053\,
            in2 => \_gnd_net_\,
            in3 => \N__9042\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__9601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9263\,
            in2 => \_gnd_net_\,
            in3 => \N__9039\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9560\,
            in2 => \_gnd_net_\,
            in3 => \N__9036\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__9603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9620\,
            in2 => \_gnd_net_\,
            in3 => \N__9246\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9533\,
            in2 => \_gnd_net_\,
            in3 => \N__9243\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__9603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9833\,
            in2 => \_gnd_net_\,
            in3 => \N__9240\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9797\,
            in2 => \_gnd_net_\,
            in3 => \N__9237\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9815\,
            in2 => \_gnd_net_\,
            in3 => \N__9234\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9228\,
            in2 => \_gnd_net_\,
            in3 => \N__9231\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_1_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011000"
        )
    port map (
            in0 => \N__10587\,
            in1 => \N__10473\,
            in2 => \N__9199\,
            in3 => \N__10449\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA_r_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001101010"
        )
    port map (
            in0 => \N__9192\,
            in1 => \N__9567\,
            in2 => \N__9216\,
            in3 => \N__10423\,
            lcout => \CLK_CIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__9168\,
            in1 => \_gnd_net_\,
            in2 => \N__9147\,
            in3 => \N__9129\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__9561\,
            in1 => \N__9549\,
            in2 => \N__9537\,
            in3 => \N__9534\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9522\,
            in1 => \N__9506\,
            in2 => \N__9417\,
            in3 => \N__9483\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9366\,
            in1 => \N__9396\,
            in2 => \N__9492\,
            in3 => \N__9489\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9609\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__9684\,
            in1 => \N__9734\,
            in2 => \N__9471\,
            in3 => \N__9786\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9609\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__9685\,
            in1 => \N__9443\,
            in2 => \N__9741\,
            in3 => \N__9785\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9609\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__9367\,
            in1 => \N__9397\,
            in2 => \N__9432\,
            in3 => \N__9329\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9609\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__9398\,
            in1 => \N__9368\,
            in2 => \N__9335\,
            in3 => \N__9275\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9609\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9621\,
            in1 => \N__9264\,
            in2 => \N__9882\,
            in3 => \N__9834\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9778\,
            in1 => \N__9740\,
            in2 => \N__9891\,
            in3 => \N__9888\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__9798\,
            in1 => \N__9867\,
            in2 => \N__9855\,
            in3 => \N__9816\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9730\,
            in1 => \N__9781\,
            in2 => \N__9682\,
            in3 => \N__9840\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9780\,
            in1 => \N__9733\,
            in2 => \N__9681\,
            in3 => \N__9822\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9731\,
            in1 => \N__9782\,
            in2 => \N__9683\,
            in3 => \N__9804\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9779\,
            in1 => \N__9732\,
            in2 => \N__9680\,
            in3 => \N__9627\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_0_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10392\,
            in1 => \N__10546\,
            in2 => \N__10518\,
            in3 => \N__9917\,
            lcout => \U409_CIA.CLK_CIA6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__9919\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10393\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__10547\,
            in1 => \N__10582\,
            in2 => \N__10517\,
            in3 => \N__9918\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_3\,
            ltout => \U409_CIA.CIA_CLK_COUNT11_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100101010"
        )
    port map (
            in0 => \N__10472\,
            in1 => \N__9942\,
            in2 => \N__9945\,
            in3 => \N__10596\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__10471\,
            in1 => \N__10445\,
            in2 => \N__10425\,
            in3 => \N__10391\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_2_0\,
            ltout => \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__9936\,
            in1 => \N__10422\,
            in2 => \N__9930\,
            in3 => \N__10557\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_1_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10515\,
            in2 => \_gnd_net_\,
            in3 => \N__10545\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA6_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__10583\,
            in1 => \N__10365\,
            in2 => \N__9927\,
            in3 => \N__9920\,
            lcout => OPEN,
            ltout => \U409_CIA.VMA_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__9921\,
            in1 => \N__10248\,
            in2 => \N__9924\,
            in3 => \N__9961\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10394\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10490\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9916\,
            in2 => \N__10395\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_7_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10443\,
            in2 => \_gnd_net_\,
            in3 => \N__9894\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__10488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10469\,
            in2 => \_gnd_net_\,
            in3 => \N__10590\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10581\,
            in2 => \_gnd_net_\,
            in3 => \N__10560\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__10488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10418\,
            in2 => \_gnd_net_\,
            in3 => \N__10551\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_6_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10548\,
            in2 => \_gnd_net_\,
            in3 => \N__10524\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\,
            clk => \N__10488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_7_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10516\,
            in2 => \_gnd_net_\,
            in3 => \N__10521\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_2_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__10470\,
            in1 => \N__10444\,
            in2 => \N__10424\,
            in3 => \N__10390\,
            lcout => \U409_CIA.un1_CIA_CLK_COUNT_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__10337\,
            in1 => \N__10299\,
            in2 => \_gnd_net_\,
            in3 => \N__10238\,
            lcout => \TCIn_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNI692L_0_LC_22_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10005\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9975\,
            lcout => \CIA_ENABLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_24_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__10709\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10658\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_24_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10659\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10640\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

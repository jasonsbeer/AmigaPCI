-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Sep 14 2025 12:26:09

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    ROM_DELAY : in std_logic_vector(1 downto 0);
    TM : in std_logic_vector(2 downto 0);
    TT : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(31 downto 1);
    D : inout std_logic_vector(7 downto 4);
    RESETn : in std_logic;
    OVL : in std_logic;
    CONFIGENn : out std_logic;
    PPIO : out std_logic;
    PORTSIZE : out std_logic;
    TICK60 : out std_logic;
    PCS1 : out std_logic;
    CIACS0n : out std_logic;
    SCS0 : out std_logic;
    CPUCONFn : in std_logic;
    CLK6 : in std_logic;
    AGNUS_CLK : out std_logic;
    CLK_CIA : out std_logic;
    BUFENn : out std_logic;
    AUTOBOOT : in std_logic;
    RnW : in std_logic;
    XCLK : in std_logic;
    CIACS1n : out std_logic;
    PPIO_J : in std_logic;
    TICK50 : out std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : out std_logic;
    PCS0 : out std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    XCLK_ENn : in std_logic;
    SCS1 : out std_logic;
    REGSPACEn : out std_logic;
    F_ENn : out std_logic;
    TSn : in std_logic;
    SPIO_J : in std_logic;
    SPIO : out std_logic;
    RTC_ENn : out std_logic;
    ATA_ENn : out std_logic;
    TACKn : inout std_logic;
    ROMENn : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__11848\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \PPIO_c\ : std_logic;
signal \GNDG0\ : std_logic;
signal \SPIO_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_27\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_5_cascade_\ : std_logic;
signal \A_c_25\ : std_logic;
signal \A_c_24\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_31\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_28\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RTC_ENn_i\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.HIROMZ0Z_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0Z0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_BASE_3C_net\ : std_logic;
signal \LIDE_BASE_6\ : std_logic;
signal \U409_AUTOCONFIG.N_99_cascade_\ : std_logic;
signal \LIDE_BASE_5\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_BASE_5C_net\ : std_logic;
signal \D_in_4\ : std_logic;
signal \U409_AUTOCONFIG.N_101\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn_i\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_5\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0Z0Z_3_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.HIROMZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.N_121_cascade_\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U409_AUTOCONFIG.N_121\ : std_logic;
signal \U409_AUTOCONFIG.N_123\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_15\ : std_logic;
signal \D_1_i\ : std_logic;
signal \U409_AUTOCONFIG.N_103\ : std_logic;
signal \LIDE_BASE_4\ : std_logic;
signal \LIDE_BASE_3\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\ : std_logic;
signal \D_in_7\ : std_logic;
signal \U409_ADDRESS_DECODE.PORTSIZEZ0Z_1\ : std_logic;
signal \U409_ADDRESS_DECODE.PORTSIZEZ0Z_0_cascade_\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \BUFENn_c\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_ATA_ENn_i\ : std_logic;
signal \A_c_18\ : std_logic;
signal \LIDE_BASE_2\ : std_logic;
signal \A_c_17\ : std_logic;
signal \LIDE_BASE_1\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_ENZ0\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUT_cnst_i_i_0_0_2\ : std_logic;
signal \INVU409_AUTOCONFIG.PR_OUT_2C_net\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1_cascade_\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U409_AUTOCONFIG.N_84\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.LOWROMZ0Z_3\ : std_logic;
signal \A_c_21\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUTZ0Z_2\ : std_logic;
signal \D_OUT_2\ : std_logic;
signal \U409_AUTOCONFIG.N_97\ : std_logic;
signal \U409_AUTOCONFIG.STATE_d_2_cascade_\ : std_logic;
signal \D_in_6\ : std_logic;
signal \U409_AUTOCONFIG.N_105\ : std_logic;
signal \U409_AUTOCONFIG.N_49\ : std_logic;
signal \D_in_5\ : std_logic;
signal \U409_AUTOCONFIG.N_49_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_107\ : std_logic;
signal \U409_AUTOCONFIG.N_95\ : std_logic;
signal \U409_AUTOCONFIG.N_48_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.un1_A_13\ : std_logic;
signal \U409_AUTOCONFIG.STATE_d_2\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_BASE_7C_net\ : std_logic;
signal \LIDE_BASE_7\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_6_0\ : std_logic;
signal \U409_AUTOCONFIG.N_48\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONFZ0\ : std_logic;
signal \INVU409_AUTOCONFIG.STATE_0C_net\ : std_logic;
signal \U409_AUTOCONFIG.STATE_ns_1_cascade_\ : std_logic;
signal \A_c_22\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1\ : std_logic;
signal \OVL_c\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\ : std_logic;
signal \U409_AUTOCONFIG.STATEZ0Z_1\ : std_logic;
signal \RnW_c\ : std_logic;
signal \CPUCONFn_c\ : std_logic;
signal \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_1_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_227_3_cascade_\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_OUT_2C_net\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.N_129\ : std_logic;
signal \U409_AUTOCONFIG.N_133_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_127\ : std_logic;
signal \U409_AUTOCONFIG.N_110\ : std_logic;
signal \A_c_4\ : std_logic;
signal \D_OUT_1\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3\ : std_logic;
signal \D_OUT_3\ : std_logic;
signal \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa\ : std_logic;
signal \CONFIGENn_c\ : std_logic;
signal \INVU409_AUTOCONFIG.CONFIGUREDC_net\ : std_logic;
signal \U409_AUTOCONFIG.N_4\ : std_logic;
signal \D_OUT_0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNI7DMPZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_CONFZ0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNI5BMPZ0Z_0\ : std_logic;
signal \AUTOCONFIG_SPACE\ : std_logic;
signal \CONFIGURED\ : std_logic;
signal \U409_AUTOCONFIG.AC_STARTZ0\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.N_82\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0Z0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUTZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.N_131\ : std_logic;
signal \U409_AUTOCONFIG.N_93\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.N_116\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.N_78\ : std_logic;
signal \U409_AUTOCONFIG.N_92\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUTZ0Z_0\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_7_i_a3_1_0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_7_i_a3_0_0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\ : std_logic;
signal \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\ : std_logic;
signal \U409_AUTOCONFIG.N_133\ : std_logic;
signal \A_c_1\ : std_logic;
signal \AUTOBOOT_c\ : std_logic;
signal \U409_AUTOCONFIG.N_126\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_7_i_1_0\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn\ : std_logic;
signal \U409_AUTOCONFIG.STATEZ0Z_0\ : std_logic;
signal \INVU409_AUTOCONFIG.AC_TACK_nesrC_net\ : std_logic;
signal \U409_AUTOCONFIG.STATE_ns_0_0_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_EN8\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_STATE_ns_1_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_STATEZ0Z_1\ : std_logic;
signal \U409_ADDRESS_DECODE_Z2_SPACE\ : std_logic;
signal \U409_ADDRESS_DECODE_HIROM\ : std_logic;
signal \TACK_OUT\ : std_logic;
signal \U409_ADDRESS_DECODE_LOWROM\ : std_logic;
signal \U409_TRANSFER_ACK_un1_TACK_OUT_0_i\ : std_logic;
signal \GB_BUFFER_CLK40_IN_c_g_THRU_CO\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_6\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\ : std_logic;
signal \U409_CIA.CLK_CIA6_4\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_\ : std_logic;
signal \CIA_SPACE\ : std_logic;
signal \U409_CIA.VMA_RNOZ0Z_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RTC_ENn\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOVECTOR_10\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_2_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_5\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTOR_4Z0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOVECTOR_11\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \CIA_ENABLE\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \U409_TRANSFER_ACK.N_5_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_1\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_2\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_3\ : std_logic;
signal \AC_TACK\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_START_2_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_STARTZ0\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_0\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_RST_0_i\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_6\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_7\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \U409_CIA.CLK_CIA6_3_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CLK_CIA_r_1_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_17_mux\ : std_logic;
signal \U409_TRANSFER_ACK.N_17_mux_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_3_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_3_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.N_7_cascade_\ : std_logic;
signal \ROM_DELAY_c_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \ROM_DELAY_c_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_19_mux\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.TICK603_8_cascade_\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \bfn_15_6_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \CLK_CIA_c\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_11\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z5\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0\ : std_logic;
signal \ROMENn_c\ : std_logic;
signal \CLK40_IN_c_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \bfn_17_5_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \bfn_17_6_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \PCS1_c\ : std_logic;
signal \SCS0_c\ : std_logic;
signal \U409_ADDRESS_DECODE.CSZ0Z0\ : std_logic;
signal \PCS0_c\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U409_ADDRESS_DECODE.CSZ0Z1\ : std_logic;
signal \SCS1_c\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \XCLK_c\ : std_logic;
signal \XCLK_ENn_c\ : std_logic;
signal \AGNUS_CLK_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK6_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \CLK28_IN_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \ROM_DELAY_wire\ : std_logic_vector(1 downto 0);
signal \CPUCONFn_wire\ : std_logic;
signal \RTC_ENn_wire\ : std_logic;
signal \SPIO_J_wire\ : std_logic;
signal \PPIO_wire\ : std_logic;
signal \PPIO_J_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \AUTOBOOT_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \F_ENn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \SCS1_wire\ : std_logic;
signal \AGNUS_CLK_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \XCLK_ENn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CONFIGENn_wire\ : std_logic;
signal \SPIO_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \ATA_ENn_wire\ : std_logic;
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \PCS0_wire\ : std_logic;
signal \CLK_CIA_wire\ : std_logic;
signal \PCS1_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \SCS0_wire\ : std_logic;
signal \XCLK_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK6_wire\ <= CLK6;
    \CLK40_IN_wire\ <= CLK40_IN;
    \CLK28_IN_wire\ <= CLK28_IN;
    \A_wire\ <= A;
    \TT_wire\ <= TT;
    \ROM_DELAY_wire\ <= ROM_DELAY;
    \CPUCONFn_wire\ <= CPUCONFn;
    RTC_ENn <= \RTC_ENn_wire\;
    \SPIO_J_wire\ <= SPIO_J;
    PPIO <= \PPIO_wire\;
    \PPIO_J_wire\ <= PPIO_J;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    TBIn <= \TBIn_wire\;
    \AUTOBOOT_wire\ <= AUTOBOOT;
    \TSn_wire\ <= TSn;
    PORTSIZE <= \PORTSIZE_wire\;
    F_ENn <= \F_ENn_wire\;
    \RESETn_wire\ <= RESETn;
    SCS1 <= \SCS1_wire\;
    AGNUS_CLK <= \AGNUS_CLK_wire\;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TCIn <= \TCIn_wire\;
    \XCLK_ENn_wire\ <= XCLK_ENn;
    \RnW_wire\ <= RnW;
    CONFIGENn <= \CONFIGENn_wire\;
    SPIO <= \SPIO_wire\;
    TICK60 <= \TICK60_wire\;
    ATA_ENn <= \ATA_ENn_wire\;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    PCS0 <= \PCS0_wire\;
    CLK_CIA <= \CLK_CIA_wire\;
    PCS1 <= \PCS1_wire\;
    BUFENn <= \BUFENn_wire\;
    SCS0 <= \SCS0_wire\;
    \XCLK_wire\ <= XCLK;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__7523\,
            RESETB => \N__11186\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11846\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11848\,
            DIN => \N__11847\,
            DOUT => \N__11846\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11848\,
            PADOUT => \N__11847\,
            PADIN => \N__11846\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11836\,
            GLOBALBUFFEROUTPUT => \CLK40_IN_c_g\
        );

    \CLK40_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11838\,
            DIN => \N__11837\,
            DOUT => \N__11836\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11838\,
            PADOUT => \N__11837\,
            PADIN => \N__11836\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11826\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11828\,
            DIN => \N__11827\,
            DOUT => \N__11826\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11828\,
            PADOUT => \N__11827\,
            PADIN => \N__11826\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11817\,
            DIN => \N__11816\,
            DOUT => \N__11815\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11817\,
            PADOUT => \N__11816\,
            PADIN => \N__11815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11808\,
            DIN => \N__11807\,
            DOUT => \N__11806\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11808\,
            PADOUT => \N__11807\,
            PADIN => \N__11806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROM_DELAY_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11799\,
            DIN => \N__11798\,
            DOUT => \N__11797\,
            PACKAGEPIN => \ROM_DELAY_wire\(1)
        );

    \ROM_DELAY_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11799\,
            PADOUT => \N__11798\,
            PADIN => \N__11797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ROM_DELAY_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11790\,
            DIN => \N__11789\,
            DOUT => \N__11788\,
            PACKAGEPIN => D(7)
        );

    \D_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11790\,
            PADOUT => \N__11789\,
            PADIN => \N__11788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4757\,
            DIN0 => \D_in_7\,
            DOUT0 => \N__6326\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11781\,
            DIN => \N__11780\,
            DOUT => \N__11779\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11781\,
            PADOUT => \N__11780\,
            PADIN => \N__11779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUCONFn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11772\,
            DIN => \N__11771\,
            DOUT => \N__11770\,
            PACKAGEPIN => \CPUCONFn_wire\
        );

    \CPUCONFn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11772\,
            PADOUT => \N__11771\,
            PADIN => \N__11770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CPUCONFn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RTC_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11763\,
            DIN => \N__11762\,
            DOUT => \N__11761\,
            PACKAGEPIN => \RTC_ENn_wire\
        );

    \RTC_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11763\,
            PADOUT => \N__11762\,
            PADIN => \N__11761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4352\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11754\,
            DIN => \N__11753\,
            DOUT => \N__11752\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11754\,
            PADOUT => \N__11753\,
            PADIN => \N__11752\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SPIO_J_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11745\,
            DIN => \N__11744\,
            DOUT => \N__11743\,
            PACKAGEPIN => \SPIO_J_wire\
        );

    \SPIO_J_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11745\,
            PADOUT => \N__11744\,
            PADIN => \N__11743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SPIO_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11736\,
            DIN => \N__11735\,
            DOUT => \N__11734\,
            PACKAGEPIN => D(4)
        );

    \D_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11736\,
            PADOUT => \N__11735\,
            PADIN => \N__11734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4742\,
            DIN0 => \D_in_4\,
            DOUT0 => \N__7022\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PPIO_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11727\,
            DIN => \N__11726\,
            DOUT => \N__11725\,
            PACKAGEPIN => \PPIO_wire\
        );

    \PPIO_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11727\,
            PADOUT => \N__11726\,
            PADIN => \N__11725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4253\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11718\,
            DIN => \N__11717\,
            DOUT => \N__11716\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11718\,
            PADOUT => \N__11717\,
            PADIN => \N__11716\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11709\,
            DIN => \N__11708\,
            DOUT => \N__11707\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11709\,
            PADOUT => \N__11708\,
            PADIN => \N__11707\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PPIO_J_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11700\,
            DIN => \N__11699\,
            DOUT => \N__11698\,
            PACKAGEPIN => \PPIO_J_wire\
        );

    \PPIO_J_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11700\,
            PADOUT => \N__11699\,
            PADIN => \N__11698\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PPIO_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11691\,
            DIN => \N__11690\,
            DOUT => \N__11689\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11691\,
            PADOUT => \N__11690\,
            PADIN => \N__11689\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6068\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11682\,
            DIN => \N__11681\,
            DOUT => \N__11680\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11682\,
            PADOUT => \N__11681\,
            PADIN => \N__11680\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11673\,
            DIN => \N__11672\,
            DOUT => \N__11671\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11673\,
            PADOUT => \N__11672\,
            PADIN => \N__11671\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9899\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11664\,
            DIN => \N__11663\,
            DOUT => \N__11662\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11664\,
            PADOUT => \N__11663\,
            PADIN => \N__11662\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9108\,
            DIN0 => OPEN,
            DOUT0 => \N__7615\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AUTOBOOT_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11655\,
            DIN => \N__11654\,
            DOUT => \N__11653\,
            PACKAGEPIN => \AUTOBOOT_wire\
        );

    \AUTOBOOT_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11655\,
            PADOUT => \N__11654\,
            PADIN => \N__11653\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AUTOBOOT_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11646\,
            DIN => \N__11645\,
            DOUT => \N__11644\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11646\,
            PADOUT => \N__11645\,
            PADIN => \N__11644\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11637\,
            DIN => \N__11636\,
            DOUT => \N__11635\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11637\,
            PADOUT => \N__11636\,
            PADIN => \N__11635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5255\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11628\,
            DIN => \N__11627\,
            DOUT => \N__11626\,
            PACKAGEPIN => \F_ENn_wire\
        );

    \F_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11628\,
            PADOUT => \N__11627\,
            PADIN => \N__11626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11176\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11619\,
            DIN => \N__11618\,
            DOUT => \N__11617\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11619\,
            PADOUT => \N__11618\,
            PADIN => \N__11617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11610\,
            DIN => \N__11609\,
            DOUT => \N__11608\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11610\,
            PADOUT => \N__11609\,
            PADIN => \N__11608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11601\,
            DIN => \N__11600\,
            DOUT => \N__11599\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11601\,
            PADOUT => \N__11600\,
            PADIN => \N__11599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11592\,
            DIN => \N__11591\,
            DOUT => \N__11590\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11592\,
            PADOUT => \N__11591\,
            PADIN => \N__11590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11583\,
            DIN => \N__11582\,
            DOUT => \N__11581\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11583\,
            PADOUT => \N__11582\,
            PADIN => \N__11581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROM_DELAY_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11574\,
            DIN => \N__11573\,
            DOUT => \N__11572\,
            PACKAGEPIN => \ROM_DELAY_wire\(0)
        );

    \ROM_DELAY_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11574\,
            PADOUT => \N__11573\,
            PADIN => \N__11572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ROM_DELAY_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11565\,
            DIN => \N__11564\,
            DOUT => \N__11563\,
            PACKAGEPIN => \SCS1_wire\
        );

    \SCS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11565\,
            PADOUT => \N__11564\,
            PADIN => \N__11563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10703\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11556\,
            DIN => \N__11555\,
            DOUT => \N__11554\,
            PACKAGEPIN => \AGNUS_CLK_wire\
        );

    \AGNUS_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11556\,
            PADOUT => \N__11555\,
            PADIN => \N__11554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11102\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11547\,
            DIN => \N__11546\,
            DOUT => \N__11545\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11547\,
            PADOUT => \N__11546\,
            PADIN => \N__11545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11538\,
            DIN => \N__11537\,
            DOUT => \N__11536\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11538\,
            PADOUT => \N__11537\,
            PADIN => \N__11536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8417\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11529\,
            DIN => \N__11528\,
            DOUT => \N__11527\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11529\,
            PADOUT => \N__11528\,
            PADIN => \N__11527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9383\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11520\,
            DIN => \N__11519\,
            DOUT => \N__11518\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11520\,
            PADOUT => \N__11519\,
            PADIN => \N__11518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11511\,
            DIN => \N__11510\,
            DOUT => \N__11509\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11511\,
            PADOUT => \N__11510\,
            PADIN => \N__11509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11502\,
            DIN => \N__11501\,
            DOUT => \N__11500\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11502\,
            PADOUT => \N__11501\,
            PADIN => \N__11500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11493\,
            DIN => \N__11492\,
            DOUT => \N__11491\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11493\,
            PADOUT => \N__11492\,
            PADIN => \N__11491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11484\,
            DIN => \N__11483\,
            DOUT => \N__11482\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11484\,
            PADOUT => \N__11483\,
            PADIN => \N__11482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9122\,
            DIN0 => OPEN,
            DOUT0 => \N__7544\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11475\,
            DIN => \N__11474\,
            DOUT => \N__11473\,
            PACKAGEPIN => D(5)
        );

    \D_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11475\,
            PADOUT => \N__11474\,
            PADIN => \N__11473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4752\,
            DIN0 => \D_in_5\,
            DOUT0 => \N__6359\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \XCLK_ENn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11466\,
            DIN => \N__11465\,
            DOUT => \N__11464\,
            PACKAGEPIN => \XCLK_ENn_wire\
        );

    \XCLK_ENn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11466\,
            PADOUT => \N__11465\,
            PADIN => \N__11464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \XCLK_ENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11457\,
            DIN => \N__11456\,
            DOUT => \N__11455\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11457\,
            PADOUT => \N__11456\,
            PADIN => \N__11455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11448\,
            DIN => \N__11447\,
            DOUT => \N__11446\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11448\,
            PADOUT => \N__11447\,
            PADIN => \N__11446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11439\,
            DIN => \N__11438\,
            DOUT => \N__11437\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11439\,
            PADOUT => \N__11438\,
            PADIN => \N__11437\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CONFIGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11430\,
            DIN => \N__11429\,
            DOUT => \N__11428\,
            PACKAGEPIN => \CONFIGENn_wire\
        );

    \CONFIGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11430\,
            PADOUT => \N__11429\,
            PADIN => \N__11428\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6299\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SPIO_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11421\,
            DIN => \N__11420\,
            DOUT => \N__11419\,
            PACKAGEPIN => \SPIO_wire\
        );

    \SPIO_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11421\,
            PADOUT => \N__11420\,
            PADIN => \N__11419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4316\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11412\,
            DIN => \N__11411\,
            DOUT => \N__11410\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11412\,
            PADOUT => \N__11411\,
            PADIN => \N__11410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9413\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11403\,
            DIN => \N__11402\,
            DOUT => \N__11401\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11403\,
            PADOUT => \N__11402\,
            PADIN => \N__11401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11394\,
            DIN => \N__11393\,
            DOUT => \N__11392\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11394\,
            PADOUT => \N__11393\,
            PADIN => \N__11392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11385\,
            DIN => \N__11384\,
            DOUT => \N__11383\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11385\,
            PADOUT => \N__11384\,
            PADIN => \N__11383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ATA_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11376\,
            DIN => \N__11375\,
            DOUT => \N__11374\,
            PACKAGEPIN => \ATA_ENn_wire\
        );

    \ATA_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11376\,
            PADOUT => \N__11375\,
            PADIN => \N__11374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5213\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11367\,
            DIN => \N__11366\,
            DOUT => \N__11365\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11367\,
            PADOUT => \N__11366\,
            PADIN => \N__11365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11358\,
            DIN => \N__11357\,
            DOUT => \N__11356\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11358\,
            PADOUT => \N__11357\,
            PADIN => \N__11356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8342\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11349\,
            DIN => \N__11348\,
            DOUT => \N__11347\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11349\,
            PADOUT => \N__11348\,
            PADIN => \N__11347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4571\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCS0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11340\,
            DIN => \N__11339\,
            DOUT => \N__11338\,
            PACKAGEPIN => \PCS0_wire\
        );

    \PCS0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11340\,
            PADOUT => \N__11339\,
            PADIN => \N__11338\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10787\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11331\,
            DIN => \N__11330\,
            DOUT => \N__11329\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11331\,
            PADOUT => \N__11330\,
            PADIN => \N__11329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_CIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11322\,
            DIN => \N__11321\,
            DOUT => \N__11320\,
            PACKAGEPIN => \CLK_CIA_wire\
        );

    \CLK_CIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11322\,
            PADOUT => \N__11321\,
            PADIN => \N__11320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9641\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11313\,
            DIN => \N__11312\,
            DOUT => \N__11311\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11313\,
            PADOUT => \N__11312\,
            PADIN => \N__11311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11304\,
            DIN => \N__11303\,
            DOUT => \N__11302\,
            PACKAGEPIN => \PCS1_wire\
        );

    \PCS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11304\,
            PADOUT => \N__11303\,
            PADIN => \N__11302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10841\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11295\,
            DIN => \N__11294\,
            DOUT => \N__11293\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11295\,
            PADOUT => \N__11294\,
            PADIN => \N__11293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9121\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__7622\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11286\,
            DIN => \N__11285\,
            DOUT => \N__11284\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11286\,
            PADOUT => \N__11285\,
            PADIN => \N__11284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11277\,
            DIN => \N__11276\,
            DOUT => \N__11275\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11277\,
            PADOUT => \N__11276\,
            PADIN => \N__11275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5234\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11268\,
            DIN => \N__11267\,
            DOUT => \N__11266\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11268\,
            PADOUT => \N__11267\,
            PADIN => \N__11266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11259\,
            DIN => \N__11258\,
            DOUT => \N__11257\,
            PACKAGEPIN => D(6)
        );

    \D_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11259\,
            PADOUT => \N__11258\,
            PADIN => \N__11257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4753\,
            DIN0 => \D_in_6\,
            DOUT0 => \N__5462\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11250\,
            DIN => \N__11249\,
            DOUT => \N__11248\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11250\,
            PADOUT => \N__11249\,
            PADIN => \N__11248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11241\,
            DIN => \N__11240\,
            DOUT => \N__11239\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11241\,
            PADOUT => \N__11240\,
            PADIN => \N__11239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCS0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11232\,
            DIN => \N__11231\,
            DOUT => \N__11230\,
            PACKAGEPIN => \SCS0_wire\
        );

    \SCS0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11232\,
            PADOUT => \N__11231\,
            PADIN => \N__11230\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10823\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \XCLK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11223\,
            DIN => \N__11222\,
            DOUT => \N__11221\,
            PACKAGEPIN => \XCLK_wire\
        );

    \XCLK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11223\,
            PADOUT => \N__11222\,
            PADIN => \N__11221\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \XCLK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11214\,
            DIN => \N__11213\,
            DOUT => \N__11212\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11214\,
            PADOUT => \N__11213\,
            PADIN => \N__11212\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11205\,
            DIN => \N__11204\,
            DOUT => \N__11203\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11205\,
            PADOUT => \N__11204\,
            PADIN => \N__11203\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2688\ : IoInMux
    port map (
            O => \N__11186\,
            I => \N__11183\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__11183\,
            I => \N__11180\
        );

    \I__2686\ : Span4Mux_s2_v
    port map (
            O => \N__11180\,
            I => \N__11177\
        );

    \I__2685\ : Sp12to4
    port map (
            O => \N__11177\,
            I => \N__11173\
        );

    \I__2684\ : IoInMux
    port map (
            O => \N__11176\,
            I => \N__11170\
        );

    \I__2683\ : Span12Mux_h
    port map (
            O => \N__11173\,
            I => \N__11167\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__11170\,
            I => \N__11164\
        );

    \I__2681\ : Span12Mux_v
    port map (
            O => \N__11167\,
            I => \N__11161\
        );

    \I__2680\ : Span12Mux_s6_h
    port map (
            O => \N__11164\,
            I => \N__11158\
        );

    \I__2679\ : Odrv12
    port map (
            O => \N__11161\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2678\ : Odrv12
    port map (
            O => \N__11158\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2677\ : InMux
    port map (
            O => \N__11153\,
            I => \N__11150\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__11150\,
            I => \N__11143\
        );

    \I__2675\ : ClkMux
    port map (
            O => \N__11149\,
            I => \N__11132\
        );

    \I__2674\ : ClkMux
    port map (
            O => \N__11148\,
            I => \N__11132\
        );

    \I__2673\ : ClkMux
    port map (
            O => \N__11147\,
            I => \N__11132\
        );

    \I__2672\ : ClkMux
    port map (
            O => \N__11146\,
            I => \N__11132\
        );

    \I__2671\ : Glb2LocalMux
    port map (
            O => \N__11143\,
            I => \N__11132\
        );

    \I__2670\ : GlobalMux
    port map (
            O => \N__11132\,
            I => \N__11129\
        );

    \I__2669\ : gio2CtrlBuf
    port map (
            O => \N__11129\,
            I => \CLK28_IN_c_g\
        );

    \I__2668\ : InMux
    port map (
            O => \N__11126\,
            I => \N__11123\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__11123\,
            I => \N__11120\
        );

    \I__2666\ : Span4Mux_v
    port map (
            O => \N__11120\,
            I => \N__11117\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__11117\,
            I => \XCLK_c\
        );

    \I__2664\ : InMux
    port map (
            O => \N__11114\,
            I => \N__11111\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__11111\,
            I => \N__11108\
        );

    \I__2662\ : Span12Mux_v
    port map (
            O => \N__11108\,
            I => \N__11105\
        );

    \I__2661\ : Odrv12
    port map (
            O => \N__11105\,
            I => \XCLK_ENn_c\
        );

    \I__2660\ : IoInMux
    port map (
            O => \N__11102\,
            I => \N__11099\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__11099\,
            I => \N__11096\
        );

    \I__2658\ : Span4Mux_s3_h
    port map (
            O => \N__11096\,
            I => \N__11093\
        );

    \I__2657\ : Odrv4
    port map (
            O => \N__11093\,
            I => \AGNUS_CLK_c\
        );

    \I__2656\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11086\
        );

    \I__2655\ : InMux
    port map (
            O => \N__11089\,
            I => \N__11083\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__11086\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__11083\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2652\ : InMux
    port map (
            O => \N__11078\,
            I => \N__11075\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__11075\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__2650\ : InMux
    port map (
            O => \N__11072\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__2649\ : InMux
    port map (
            O => \N__11069\,
            I => \N__11065\
        );

    \I__2648\ : InMux
    port map (
            O => \N__11068\,
            I => \N__11062\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__11065\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__11062\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__2645\ : InMux
    port map (
            O => \N__11057\,
            I => \N__11054\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__11054\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__2643\ : InMux
    port map (
            O => \N__11051\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__2642\ : InMux
    port map (
            O => \N__11048\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__2641\ : InMux
    port map (
            O => \N__11045\,
            I => \N__11041\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11044\,
            I => \N__11038\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__11041\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__11038\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__11033\,
            I => \N__11025\
        );

    \I__2636\ : InMux
    port map (
            O => \N__11032\,
            I => \N__11018\
        );

    \I__2635\ : InMux
    port map (
            O => \N__11031\,
            I => \N__11018\
        );

    \I__2634\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11015\
        );

    \I__2633\ : InMux
    port map (
            O => \N__11029\,
            I => \N__11012\
        );

    \I__2632\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11003\
        );

    \I__2631\ : InMux
    port map (
            O => \N__11025\,
            I => \N__11003\
        );

    \I__2630\ : InMux
    port map (
            O => \N__11024\,
            I => \N__11003\
        );

    \I__2629\ : InMux
    port map (
            O => \N__11023\,
            I => \N__11003\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__11018\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__11015\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__11012\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__11003\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__10994\,
            I => \N__10990\
        );

    \I__2623\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10984\
        );

    \I__2622\ : InMux
    port map (
            O => \N__10990\,
            I => \N__10978\
        );

    \I__2621\ : InMux
    port map (
            O => \N__10989\,
            I => \N__10975\
        );

    \I__2620\ : InMux
    port map (
            O => \N__10988\,
            I => \N__10972\
        );

    \I__2619\ : InMux
    port map (
            O => \N__10987\,
            I => \N__10969\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__10984\,
            I => \N__10966\
        );

    \I__2617\ : InMux
    port map (
            O => \N__10983\,
            I => \N__10959\
        );

    \I__2616\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10959\
        );

    \I__2615\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10959\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__10978\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__10975\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__10972\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__10969\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__10966\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__10959\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__10946\,
            I => \N__10942\
        );

    \I__2607\ : InMux
    port map (
            O => \N__10945\,
            I => \N__10936\
        );

    \I__2606\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10936\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__10941\,
            I => \N__10933\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__10936\,
            I => \N__10925\
        );

    \I__2603\ : InMux
    port map (
            O => \N__10933\,
            I => \N__10922\
        );

    \I__2602\ : InMux
    port map (
            O => \N__10932\,
            I => \N__10911\
        );

    \I__2601\ : InMux
    port map (
            O => \N__10931\,
            I => \N__10911\
        );

    \I__2600\ : InMux
    port map (
            O => \N__10930\,
            I => \N__10911\
        );

    \I__2599\ : InMux
    port map (
            O => \N__10929\,
            I => \N__10911\
        );

    \I__2598\ : InMux
    port map (
            O => \N__10928\,
            I => \N__10911\
        );

    \I__2597\ : Span4Mux_h
    port map (
            O => \N__10925\,
            I => \N__10908\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__10922\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__10911\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__10908\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2593\ : InMux
    port map (
            O => \N__10901\,
            I => \N__10898\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__10898\,
            I => \N__10895\
        );

    \I__2591\ : Odrv4
    port map (
            O => \N__10895\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__2590\ : InMux
    port map (
            O => \N__10892\,
            I => \N__10888\
        );

    \I__2589\ : InMux
    port map (
            O => \N__10891\,
            I => \N__10885\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__10888\,
            I => \N__10882\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__10885\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2586\ : Odrv12
    port map (
            O => \N__10882\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2585\ : ClkMux
    port map (
            O => \N__10877\,
            I => \N__10847\
        );

    \I__2584\ : ClkMux
    port map (
            O => \N__10876\,
            I => \N__10847\
        );

    \I__2583\ : ClkMux
    port map (
            O => \N__10875\,
            I => \N__10847\
        );

    \I__2582\ : ClkMux
    port map (
            O => \N__10874\,
            I => \N__10847\
        );

    \I__2581\ : ClkMux
    port map (
            O => \N__10873\,
            I => \N__10847\
        );

    \I__2580\ : ClkMux
    port map (
            O => \N__10872\,
            I => \N__10847\
        );

    \I__2579\ : ClkMux
    port map (
            O => \N__10871\,
            I => \N__10847\
        );

    \I__2578\ : ClkMux
    port map (
            O => \N__10870\,
            I => \N__10847\
        );

    \I__2577\ : ClkMux
    port map (
            O => \N__10869\,
            I => \N__10847\
        );

    \I__2576\ : ClkMux
    port map (
            O => \N__10868\,
            I => \N__10847\
        );

    \I__2575\ : GlobalMux
    port map (
            O => \N__10847\,
            I => \N__10844\
        );

    \I__2574\ : gio2CtrlBuf
    port map (
            O => \N__10844\,
            I => \CLK6_c_g\
        );

    \I__2573\ : IoInMux
    port map (
            O => \N__10841\,
            I => \N__10838\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__10838\,
            I => \N__10835\
        );

    \I__2571\ : Span4Mux_s3_h
    port map (
            O => \N__10835\,
            I => \N__10832\
        );

    \I__2570\ : Span4Mux_v
    port map (
            O => \N__10832\,
            I => \N__10829\
        );

    \I__2569\ : Span4Mux_h
    port map (
            O => \N__10829\,
            I => \N__10826\
        );

    \I__2568\ : Odrv4
    port map (
            O => \N__10826\,
            I => \PCS1_c\
        );

    \I__2567\ : IoInMux
    port map (
            O => \N__10823\,
            I => \N__10820\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__10820\,
            I => \N__10817\
        );

    \I__2565\ : IoSpan4Mux
    port map (
            O => \N__10817\,
            I => \N__10814\
        );

    \I__2564\ : Span4Mux_s3_h
    port map (
            O => \N__10814\,
            I => \N__10811\
        );

    \I__2563\ : Span4Mux_h
    port map (
            O => \N__10811\,
            I => \N__10808\
        );

    \I__2562\ : Odrv4
    port map (
            O => \N__10808\,
            I => \SCS0_c\
        );

    \I__2561\ : InMux
    port map (
            O => \N__10805\,
            I => \N__10801\
        );

    \I__2560\ : InMux
    port map (
            O => \N__10804\,
            I => \N__10798\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__10801\,
            I => \N__10793\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__10798\,
            I => \N__10793\
        );

    \I__2557\ : Span12Mux_s10_h
    port map (
            O => \N__10793\,
            I => \N__10790\
        );

    \I__2556\ : Odrv12
    port map (
            O => \N__10790\,
            I => \U409_ADDRESS_DECODE.CSZ0Z0\
        );

    \I__2555\ : IoInMux
    port map (
            O => \N__10787\,
            I => \N__10784\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__10784\,
            I => \N__10781\
        );

    \I__2553\ : IoSpan4Mux
    port map (
            O => \N__10781\,
            I => \N__10778\
        );

    \I__2552\ : Span4Mux_s3_v
    port map (
            O => \N__10778\,
            I => \N__10775\
        );

    \I__2551\ : Span4Mux_v
    port map (
            O => \N__10775\,
            I => \N__10772\
        );

    \I__2550\ : Odrv4
    port map (
            O => \N__10772\,
            I => \PCS0_c\
        );

    \I__2549\ : InMux
    port map (
            O => \N__10769\,
            I => \N__10763\
        );

    \I__2548\ : InMux
    port map (
            O => \N__10768\,
            I => \N__10760\
        );

    \I__2547\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10757\
        );

    \I__2546\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10754\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__10763\,
            I => \N__10749\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__10760\,
            I => \N__10749\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__10757\,
            I => \N__10744\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__10754\,
            I => \N__10744\
        );

    \I__2541\ : Span4Mux_v
    port map (
            O => \N__10749\,
            I => \N__10741\
        );

    \I__2540\ : Span4Mux_v
    port map (
            O => \N__10744\,
            I => \N__10738\
        );

    \I__2539\ : Sp12to4
    port map (
            O => \N__10741\,
            I => \N__10735\
        );

    \I__2538\ : Span4Mux_h
    port map (
            O => \N__10738\,
            I => \N__10732\
        );

    \I__2537\ : Span12Mux_h
    port map (
            O => \N__10735\,
            I => \N__10727\
        );

    \I__2536\ : Sp12to4
    port map (
            O => \N__10732\,
            I => \N__10727\
        );

    \I__2535\ : Span12Mux_h
    port map (
            O => \N__10727\,
            I => \N__10724\
        );

    \I__2534\ : Odrv12
    port map (
            O => \N__10724\,
            I => \A_c_14\
        );

    \I__2533\ : InMux
    port map (
            O => \N__10721\,
            I => \N__10717\
        );

    \I__2532\ : InMux
    port map (
            O => \N__10720\,
            I => \N__10714\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__10717\,
            I => \N__10709\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__10714\,
            I => \N__10709\
        );

    \I__2529\ : Span12Mux_h
    port map (
            O => \N__10709\,
            I => \N__10706\
        );

    \I__2528\ : Odrv12
    port map (
            O => \N__10706\,
            I => \U409_ADDRESS_DECODE.CSZ0Z1\
        );

    \I__2527\ : IoInMux
    port map (
            O => \N__10703\,
            I => \N__10700\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__2525\ : IoSpan4Mux
    port map (
            O => \N__10697\,
            I => \N__10694\
        );

    \I__2524\ : IoSpan4Mux
    port map (
            O => \N__10694\,
            I => \N__10691\
        );

    \I__2523\ : Span4Mux_s3_h
    port map (
            O => \N__10691\,
            I => \N__10688\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__10688\,
            I => \SCS1_c\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__10685\,
            I => \N__10682\
        );

    \I__2520\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10678\
        );

    \I__2519\ : InMux
    port map (
            O => \N__10681\,
            I => \N__10675\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__10678\,
            I => \N__10670\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__10675\,
            I => \N__10670\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__10670\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2515\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10664\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__10664\,
            I => \N__10661\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__10661\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__2512\ : InMux
    port map (
            O => \N__10658\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10655\,
            I => \N__10651\
        );

    \I__2510\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10648\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__10651\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10648\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__2507\ : InMux
    port map (
            O => \N__10643\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10640\,
            I => \N__10636\
        );

    \I__2505\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10633\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__10636\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10633\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2502\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10625\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__10625\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10622\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__2499\ : InMux
    port map (
            O => \N__10619\,
            I => \N__10615\
        );

    \I__2498\ : InMux
    port map (
            O => \N__10618\,
            I => \N__10612\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__10615\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10612\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2495\ : CascadeMux
    port map (
            O => \N__10607\,
            I => \N__10604\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10604\,
            I => \N__10601\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__10601\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10598\,
            I => \bfn_17_6_0_\
        );

    \I__2491\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10591\
        );

    \I__2490\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10588\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__10591\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__10588\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__2487\ : InMux
    port map (
            O => \N__10583\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__2486\ : InMux
    port map (
            O => \N__10580\,
            I => \N__10577\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__10577\,
            I => \N__10574\
        );

    \I__2484\ : Span4Mux_h
    port map (
            O => \N__10574\,
            I => \N__10570\
        );

    \I__2483\ : InMux
    port map (
            O => \N__10573\,
            I => \N__10567\
        );

    \I__2482\ : Odrv4
    port map (
            O => \N__10570\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__10567\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__2480\ : InMux
    port map (
            O => \N__10562\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__2479\ : InMux
    port map (
            O => \N__10559\,
            I => \N__10555\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10558\,
            I => \N__10552\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__10555\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__10552\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__2475\ : InMux
    port map (
            O => \N__10547\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__10544\,
            I => \N__10541\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10541\,
            I => \N__10537\
        );

    \I__2472\ : InMux
    port map (
            O => \N__10540\,
            I => \N__10534\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__10537\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__10534\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__2469\ : InMux
    port map (
            O => \N__10529\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__2468\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10523\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__10523\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__2466\ : InMux
    port map (
            O => \N__10520\,
            I => \N__10516\
        );

    \I__2465\ : InMux
    port map (
            O => \N__10519\,
            I => \N__10513\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__10516\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__10513\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2462\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10504\
        );

    \I__2461\ : InMux
    port map (
            O => \N__10507\,
            I => \N__10501\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__10504\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__10501\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__10496\,
            I => \N__10493\
        );

    \I__2457\ : InMux
    port map (
            O => \N__10493\,
            I => \N__10489\
        );

    \I__2456\ : InMux
    port map (
            O => \N__10492\,
            I => \N__10486\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__10489\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__10486\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10481\,
            I => \N__10477\
        );

    \I__2452\ : InMux
    port map (
            O => \N__10480\,
            I => \N__10474\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__10477\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10474\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__2449\ : CascadeMux
    port map (
            O => \N__10469\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__2448\ : InMux
    port map (
            O => \N__10466\,
            I => \N__10463\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__10463\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__2446\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10456\
        );

    \I__2445\ : InMux
    port map (
            O => \N__10459\,
            I => \N__10453\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__10456\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__10453\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__10448\,
            I => \N__10444\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10447\,
            I => \N__10438\
        );

    \I__2440\ : InMux
    port map (
            O => \N__10444\,
            I => \N__10438\
        );

    \I__2439\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10435\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__10438\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10435\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2436\ : CascadeMux
    port map (
            O => \N__10430\,
            I => \N__10426\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__10429\,
            I => \N__10421\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10426\,
            I => \N__10416\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10425\,
            I => \N__10416\
        );

    \I__2432\ : InMux
    port map (
            O => \N__10424\,
            I => \N__10413\
        );

    \I__2431\ : InMux
    port map (
            O => \N__10421\,
            I => \N__10410\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__10416\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__10413\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__10410\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2427\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10399\
        );

    \I__2426\ : InMux
    port map (
            O => \N__10402\,
            I => \N__10396\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10399\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__10396\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__2423\ : InMux
    port map (
            O => \N__10391\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__10385\,
            I => \N__10381\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10384\,
            I => \N__10378\
        );

    \I__2419\ : Odrv4
    port map (
            O => \N__10381\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__10378\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10373\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10363\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10366\,
            I => \N__10360\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__10363\,
            I => \N__10357\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__10360\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__2411\ : Odrv12
    port map (
            O => \N__10357\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__10349\,
            I => \N__10346\
        );

    \I__2408\ : Odrv4
    port map (
            O => \N__10346\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10343\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__2406\ : InMux
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__10337\,
            I => \N__10333\
        );

    \I__2404\ : InMux
    port map (
            O => \N__10336\,
            I => \N__10330\
        );

    \I__2403\ : Odrv4
    port map (
            O => \N__10333\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__10330\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__2401\ : InMux
    port map (
            O => \N__10325\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__10322\,
            I => \N__10314\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__10321\,
            I => \N__10311\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10320\,
            I => \N__10303\
        );

    \I__2397\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10303\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10318\,
            I => \N__10303\
        );

    \I__2395\ : InMux
    port map (
            O => \N__10317\,
            I => \N__10294\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10314\,
            I => \N__10294\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10311\,
            I => \N__10294\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10294\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__10303\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__10294\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10289\,
            I => \N__10272\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10288\,
            I => \N__10272\
        );

    \I__2387\ : InMux
    port map (
            O => \N__10287\,
            I => \N__10272\
        );

    \I__2386\ : InMux
    port map (
            O => \N__10286\,
            I => \N__10272\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10285\,
            I => \N__10272\
        );

    \I__2384\ : InMux
    port map (
            O => \N__10284\,
            I => \N__10267\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10267\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__10272\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10267\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__10262\,
            I => \N__10259\
        );

    \I__2379\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10250\
        );

    \I__2378\ : InMux
    port map (
            O => \N__10258\,
            I => \N__10247\
        );

    \I__2377\ : InMux
    port map (
            O => \N__10257\,
            I => \N__10236\
        );

    \I__2376\ : InMux
    port map (
            O => \N__10256\,
            I => \N__10236\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10255\,
            I => \N__10236\
        );

    \I__2374\ : InMux
    port map (
            O => \N__10254\,
            I => \N__10236\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10236\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10250\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10247\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__10236\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__10229\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10226\,
            I => \N__10222\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10225\,
            I => \N__10219\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__10222\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__10219\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10214\,
            I => \N__10211\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10211\,
            I => \N__10208\
        );

    \I__2362\ : Odrv12
    port map (
            O => \N__10208\,
            I => \U409_TICK.TICK503_11\
        );

    \I__2361\ : InMux
    port map (
            O => \N__10205\,
            I => \N__10201\
        );

    \I__2360\ : InMux
    port map (
            O => \N__10204\,
            I => \N__10198\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10201\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__10198\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2357\ : CascadeMux
    port map (
            O => \N__10193\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__2356\ : InMux
    port map (
            O => \N__10190\,
            I => \N__10186\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10189\,
            I => \N__10183\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__10186\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__10183\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__10178\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__2351\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10172\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10172\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10166\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__10166\,
            I => \N__10161\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__10165\,
            I => \N__10158\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__10164\,
            I => \N__10154\
        );

    \I__2345\ : Span4Mux_h
    port map (
            O => \N__10161\,
            I => \N__10151\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10158\,
            I => \N__10146\
        );

    \I__2343\ : InMux
    port map (
            O => \N__10157\,
            I => \N__10146\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10143\
        );

    \I__2341\ : Odrv4
    port map (
            O => \N__10151\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__10146\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10143\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10133\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__10133\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__2336\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10126\
        );

    \I__2335\ : InMux
    port map (
            O => \N__10129\,
            I => \N__10123\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__10126\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__10123\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__2332\ : InMux
    port map (
            O => \N__10118\,
            I => \N__10114\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10117\,
            I => \N__10111\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__10114\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10111\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2328\ : CascadeMux
    port map (
            O => \N__10106\,
            I => \N__10103\
        );

    \I__2327\ : InMux
    port map (
            O => \N__10103\,
            I => \N__10099\
        );

    \I__2326\ : InMux
    port map (
            O => \N__10102\,
            I => \N__10096\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10099\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__10096\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__10091\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10088\,
            I => \N__10085\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__10085\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__2320\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10077\
        );

    \I__2319\ : InMux
    port map (
            O => \N__10081\,
            I => \N__10072\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10080\,
            I => \N__10072\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__10077\,
            I => \U409_TRANSFER_ACK.N_11\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__10072\,
            I => \U409_TRANSFER_ACK.N_11\
        );

    \I__2315\ : InMux
    port map (
            O => \N__10067\,
            I => \N__10064\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__10064\,
            I => \N__10059\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10063\,
            I => \N__10053\
        );

    \I__2312\ : InMux
    port map (
            O => \N__10062\,
            I => \N__10053\
        );

    \I__2311\ : Span4Mux_h
    port map (
            O => \N__10059\,
            I => \N__10050\
        );

    \I__2310\ : InMux
    port map (
            O => \N__10058\,
            I => \N__10047\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__10053\,
            I => \N__10044\
        );

    \I__2308\ : Odrv4
    port map (
            O => \N__10050\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__10047\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__2306\ : Odrv12
    port map (
            O => \N__10044\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10037\,
            I => \N__10027\
        );

    \I__2304\ : InMux
    port map (
            O => \N__10036\,
            I => \N__10027\
        );

    \I__2303\ : InMux
    port map (
            O => \N__10035\,
            I => \N__10027\
        );

    \I__2302\ : InMux
    port map (
            O => \N__10034\,
            I => \N__10024\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10027\,
            I => \N__10020\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__10024\,
            I => \N__10017\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__10023\,
            I => \N__10012\
        );

    \I__2298\ : Span4Mux_v
    port map (
            O => \N__10020\,
            I => \N__10006\
        );

    \I__2297\ : Span4Mux_v
    port map (
            O => \N__10017\,
            I => \N__10006\
        );

    \I__2296\ : InMux
    port map (
            O => \N__10016\,
            I => \N__10003\
        );

    \I__2295\ : InMux
    port map (
            O => \N__10015\,
            I => \N__10000\
        );

    \I__2294\ : InMux
    port map (
            O => \N__10012\,
            I => \N__9995\
        );

    \I__2293\ : InMux
    port map (
            O => \N__10011\,
            I => \N__9995\
        );

    \I__2292\ : Odrv4
    port map (
            O => \N__10006\,
            I => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_1\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__10003\,
            I => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_1\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__10000\,
            I => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_1\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__9995\,
            I => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_1\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__9986\,
            I => \N__9983\
        );

    \I__2287\ : InMux
    port map (
            O => \N__9983\,
            I => \N__9979\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__9982\,
            I => \N__9976\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__9979\,
            I => \N__9973\
        );

    \I__2284\ : InMux
    port map (
            O => \N__9976\,
            I => \N__9970\
        );

    \I__2283\ : Span4Mux_h
    port map (
            O => \N__9973\,
            I => \N__9965\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__9970\,
            I => \N__9965\
        );

    \I__2281\ : Span4Mux_h
    port map (
            O => \N__9965\,
            I => \N__9962\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__9962\,
            I => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z5\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__9959\,
            I => \N__9953\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__9958\,
            I => \N__9950\
        );

    \I__2277\ : InMux
    port map (
            O => \N__9957\,
            I => \N__9940\
        );

    \I__2276\ : InMux
    port map (
            O => \N__9956\,
            I => \N__9940\
        );

    \I__2275\ : InMux
    port map (
            O => \N__9953\,
            I => \N__9940\
        );

    \I__2274\ : InMux
    port map (
            O => \N__9950\,
            I => \N__9940\
        );

    \I__2273\ : InMux
    port map (
            O => \N__9949\,
            I => \N__9937\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__9940\,
            I => \N__9927\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__9937\,
            I => \N__9927\
        );

    \I__2270\ : InMux
    port map (
            O => \N__9936\,
            I => \N__9924\
        );

    \I__2269\ : InMux
    port map (
            O => \N__9935\,
            I => \N__9921\
        );

    \I__2268\ : InMux
    port map (
            O => \N__9934\,
            I => \N__9918\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9933\,
            I => \N__9913\
        );

    \I__2266\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9913\
        );

    \I__2265\ : Span4Mux_h
    port map (
            O => \N__9927\,
            I => \N__9910\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__9924\,
            I => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__9921\,
            I => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__9918\,
            I => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__9913\,
            I => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__9910\,
            I => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0\
        );

    \I__2259\ : IoInMux
    port map (
            O => \N__9899\,
            I => \N__9896\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__9896\,
            I => \N__9893\
        );

    \I__2257\ : Span4Mux_s1_v
    port map (
            O => \N__9893\,
            I => \N__9890\
        );

    \I__2256\ : Span4Mux_v
    port map (
            O => \N__9890\,
            I => \N__9887\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__9887\,
            I => \N__9884\
        );

    \I__2254\ : Span4Mux_v
    port map (
            O => \N__9884\,
            I => \N__9880\
        );

    \I__2253\ : InMux
    port map (
            O => \N__9883\,
            I => \N__9877\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__9880\,
            I => \ROMENn_c\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__9877\,
            I => \ROMENn_c\
        );

    \I__2250\ : CascadeMux
    port map (
            O => \N__9872\,
            I => \N__9866\
        );

    \I__2249\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9861\
        );

    \I__2248\ : InMux
    port map (
            O => \N__9870\,
            I => \N__9858\
        );

    \I__2247\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9855\
        );

    \I__2246\ : InMux
    port map (
            O => \N__9866\,
            I => \N__9852\
        );

    \I__2245\ : InMux
    port map (
            O => \N__9865\,
            I => \N__9847\
        );

    \I__2244\ : InMux
    port map (
            O => \N__9864\,
            I => \N__9847\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__9861\,
            I => \N__9843\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__9858\,
            I => \N__9834\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__9855\,
            I => \N__9827\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__9852\,
            I => \N__9815\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__9847\,
            I => \N__9812\
        );

    \I__2238\ : ClkMux
    port map (
            O => \N__9846\,
            I => \N__9761\
        );

    \I__2237\ : Glb2LocalMux
    port map (
            O => \N__9843\,
            I => \N__9761\
        );

    \I__2236\ : ClkMux
    port map (
            O => \N__9842\,
            I => \N__9761\
        );

    \I__2235\ : ClkMux
    port map (
            O => \N__9841\,
            I => \N__9761\
        );

    \I__2234\ : ClkMux
    port map (
            O => \N__9840\,
            I => \N__9761\
        );

    \I__2233\ : ClkMux
    port map (
            O => \N__9839\,
            I => \N__9761\
        );

    \I__2232\ : ClkMux
    port map (
            O => \N__9838\,
            I => \N__9761\
        );

    \I__2231\ : ClkMux
    port map (
            O => \N__9837\,
            I => \N__9761\
        );

    \I__2230\ : Glb2LocalMux
    port map (
            O => \N__9834\,
            I => \N__9761\
        );

    \I__2229\ : ClkMux
    port map (
            O => \N__9833\,
            I => \N__9761\
        );

    \I__2228\ : ClkMux
    port map (
            O => \N__9832\,
            I => \N__9761\
        );

    \I__2227\ : ClkMux
    port map (
            O => \N__9831\,
            I => \N__9761\
        );

    \I__2226\ : ClkMux
    port map (
            O => \N__9830\,
            I => \N__9761\
        );

    \I__2225\ : Glb2LocalMux
    port map (
            O => \N__9827\,
            I => \N__9761\
        );

    \I__2224\ : ClkMux
    port map (
            O => \N__9826\,
            I => \N__9761\
        );

    \I__2223\ : ClkMux
    port map (
            O => \N__9825\,
            I => \N__9761\
        );

    \I__2222\ : ClkMux
    port map (
            O => \N__9824\,
            I => \N__9761\
        );

    \I__2221\ : ClkMux
    port map (
            O => \N__9823\,
            I => \N__9761\
        );

    \I__2220\ : ClkMux
    port map (
            O => \N__9822\,
            I => \N__9761\
        );

    \I__2219\ : ClkMux
    port map (
            O => \N__9821\,
            I => \N__9761\
        );

    \I__2218\ : ClkMux
    port map (
            O => \N__9820\,
            I => \N__9761\
        );

    \I__2217\ : ClkMux
    port map (
            O => \N__9819\,
            I => \N__9761\
        );

    \I__2216\ : ClkMux
    port map (
            O => \N__9818\,
            I => \N__9761\
        );

    \I__2215\ : Glb2LocalMux
    port map (
            O => \N__9815\,
            I => \N__9761\
        );

    \I__2214\ : Glb2LocalMux
    port map (
            O => \N__9812\,
            I => \N__9761\
        );

    \I__2213\ : GlobalMux
    port map (
            O => \N__9761\,
            I => \N__9758\
        );

    \I__2212\ : gio2CtrlBuf
    port map (
            O => \N__9758\,
            I => \CLK40_IN_c_g\
        );

    \I__2211\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9752\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9752\,
            I => \N__9740\
        );

    \I__2209\ : SRMux
    port map (
            O => \N__9751\,
            I => \N__9692\
        );

    \I__2208\ : SRMux
    port map (
            O => \N__9750\,
            I => \N__9692\
        );

    \I__2207\ : SRMux
    port map (
            O => \N__9749\,
            I => \N__9692\
        );

    \I__2206\ : SRMux
    port map (
            O => \N__9748\,
            I => \N__9692\
        );

    \I__2205\ : SRMux
    port map (
            O => \N__9747\,
            I => \N__9692\
        );

    \I__2204\ : SRMux
    port map (
            O => \N__9746\,
            I => \N__9692\
        );

    \I__2203\ : SRMux
    port map (
            O => \N__9745\,
            I => \N__9692\
        );

    \I__2202\ : SRMux
    port map (
            O => \N__9744\,
            I => \N__9692\
        );

    \I__2201\ : SRMux
    port map (
            O => \N__9743\,
            I => \N__9692\
        );

    \I__2200\ : Glb2LocalMux
    port map (
            O => \N__9740\,
            I => \N__9692\
        );

    \I__2199\ : SRMux
    port map (
            O => \N__9739\,
            I => \N__9692\
        );

    \I__2198\ : SRMux
    port map (
            O => \N__9738\,
            I => \N__9692\
        );

    \I__2197\ : SRMux
    port map (
            O => \N__9737\,
            I => \N__9692\
        );

    \I__2196\ : SRMux
    port map (
            O => \N__9736\,
            I => \N__9692\
        );

    \I__2195\ : SRMux
    port map (
            O => \N__9735\,
            I => \N__9692\
        );

    \I__2194\ : SRMux
    port map (
            O => \N__9734\,
            I => \N__9692\
        );

    \I__2193\ : SRMux
    port map (
            O => \N__9733\,
            I => \N__9692\
        );

    \I__2192\ : SRMux
    port map (
            O => \N__9732\,
            I => \N__9692\
        );

    \I__2191\ : SRMux
    port map (
            O => \N__9731\,
            I => \N__9692\
        );

    \I__2190\ : GlobalMux
    port map (
            O => \N__9692\,
            I => \N__9689\
        );

    \I__2189\ : gio2CtrlBuf
    port map (
            O => \N__9689\,
            I => \RESETn_c_i_g\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9686\,
            I => \N__9683\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__9683\,
            I => \U409_TICK.TICK603_11\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9680\,
            I => \bfn_15_7_0_\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9677\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9674\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9671\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9668\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__2181\ : InMux
    port map (
            O => \N__9665\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9662\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9659\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__2178\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9652\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9655\,
            I => \N__9649\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9652\,
            I => \N__9646\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__9649\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__9646\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__2173\ : IoInMux
    port map (
            O => \N__9641\,
            I => \N__9638\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9638\,
            I => \N__9635\
        );

    \I__2171\ : IoSpan4Mux
    port map (
            O => \N__9635\,
            I => \N__9632\
        );

    \I__2170\ : Span4Mux_s0_v
    port map (
            O => \N__9632\,
            I => \N__9629\
        );

    \I__2169\ : Sp12to4
    port map (
            O => \N__9629\,
            I => \N__9624\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9621\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__9627\,
            I => \N__9617\
        );

    \I__2166\ : Span12Mux_s11_v
    port map (
            O => \N__9624\,
            I => \N__9614\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9621\,
            I => \N__9611\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9606\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9606\
        );

    \I__2162\ : Odrv12
    port map (
            O => \N__9614\,
            I => \CLK_CIA_c\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__9611\,
            I => \CLK_CIA_c\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__9606\,
            I => \CLK_CIA_c\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9594\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9598\,
            I => \N__9589\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9597\,
            I => \N__9589\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__9594\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9589\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9584\,
            I => \N__9579\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9583\,
            I => \N__9576\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9582\,
            I => \N__9573\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__9579\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__9576\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9573\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9562\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9565\,
            I => \N__9559\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__9562\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__9559\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9554\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9551\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9548\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__2141\ : InMux
    port map (
            O => \N__9545\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__9542\,
            I => \N__9539\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9536\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9536\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9533\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9530\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__2135\ : CascadeMux
    port map (
            O => \N__9527\,
            I => \N__9524\
        );

    \I__2134\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9520\
        );

    \I__2133\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9517\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9520\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9517\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9512\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__9509\,
            I => \N__9505\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9508\,
            I => \N__9500\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9505\,
            I => \N__9500\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__9500\,
            I => \N__9497\
        );

    \I__2125\ : Span4Mux_v
    port map (
            O => \N__9497\,
            I => \N__9494\
        );

    \I__2124\ : Sp12to4
    port map (
            O => \N__9494\,
            I => \N__9491\
        );

    \I__2123\ : Span12Mux_v
    port map (
            O => \N__9491\,
            I => \N__9488\
        );

    \I__2122\ : Span12Mux_h
    port map (
            O => \N__9488\,
            I => \N__9485\
        );

    \I__2121\ : Odrv12
    port map (
            O => \N__9485\,
            I => \ROM_DELAY_c_0\
        );

    \I__2120\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9475\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9475\
        );

    \I__2118\ : InMux
    port map (
            O => \N__9480\,
            I => \N__9472\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9475\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__9472\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__9467\,
            I => \N__9464\
        );

    \I__2114\ : InMux
    port map (
            O => \N__9464\,
            I => \N__9458\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9463\,
            I => \N__9458\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__2111\ : Span4Mux_h
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__2110\ : Span4Mux_v
    port map (
            O => \N__9452\,
            I => \N__9449\
        );

    \I__2109\ : Sp12to4
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__2108\ : Span12Mux_h
    port map (
            O => \N__9446\,
            I => \N__9443\
        );

    \I__2107\ : Span12Mux_v
    port map (
            O => \N__9443\,
            I => \N__9440\
        );

    \I__2106\ : Odrv12
    port map (
            O => \N__9440\,
            I => \ROM_DELAY_c_1\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9432\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9436\,
            I => \N__9427\
        );

    \I__2103\ : InMux
    port map (
            O => \N__9435\,
            I => \N__9427\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__9432\,
            I => \N__9424\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9427\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__9424\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9416\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__9416\,
            I => \U409_TRANSFER_ACK.N_19_mux\
        );

    \I__2097\ : IoInMux
    port map (
            O => \N__9413\,
            I => \N__9410\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__9410\,
            I => \N__9407\
        );

    \I__2095\ : IoSpan4Mux
    port map (
            O => \N__9407\,
            I => \N__9404\
        );

    \I__2094\ : Span4Mux_s2_v
    port map (
            O => \N__9404\,
            I => \N__9401\
        );

    \I__2093\ : Sp12to4
    port map (
            O => \N__9401\,
            I => \N__9398\
        );

    \I__2092\ : Span12Mux_s10_v
    port map (
            O => \N__9398\,
            I => \N__9394\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9391\
        );

    \I__2090\ : Odrv12
    port map (
            O => \N__9394\,
            I => \TICK60_c\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__9391\,
            I => \TICK60_c\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__9386\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__2087\ : IoInMux
    port map (
            O => \N__9383\,
            I => \N__9380\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9380\,
            I => \N__9377\
        );

    \I__2085\ : Span4Mux_s1_v
    port map (
            O => \N__9377\,
            I => \N__9374\
        );

    \I__2084\ : Sp12to4
    port map (
            O => \N__9374\,
            I => \N__9371\
        );

    \I__2083\ : Span12Mux_h
    port map (
            O => \N__9371\,
            I => \N__9367\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9364\
        );

    \I__2081\ : Odrv12
    port map (
            O => \N__9367\,
            I => \TICK50_c\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9364\,
            I => \TICK50_c\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__9359\,
            I => \U409_TICK.TICK603_8_cascade_\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__9356\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9353\,
            I => \N__9350\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9350\,
            I => \U409_TRANSFER_ACK.N_17_mux\
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__9347\,
            I => \U409_TRANSFER_ACK.N_17_mux_cascade_\
        );

    \I__2074\ : InMux
    port map (
            O => \N__9344\,
            I => \N__9341\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__9341\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0\
        );

    \I__2072\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9335\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__9335\,
            I => \U409_TRANSFER_ACK.N_3_0\
        );

    \I__2070\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9326\
        );

    \I__2069\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9323\
        );

    \I__2068\ : InMux
    port map (
            O => \N__9330\,
            I => \N__9318\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9318\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9326\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9323\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__9318\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9306\
        );

    \I__2062\ : InMux
    port map (
            O => \N__9310\,
            I => \N__9301\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9309\,
            I => \N__9301\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__9306\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9301\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__9296\,
            I => \U409_TRANSFER_ACK.N_3_0_cascade_\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9293\,
            I => \N__9287\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9292\,
            I => \N__9284\
        );

    \I__2055\ : InMux
    port map (
            O => \N__9291\,
            I => \N__9279\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9279\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9287\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9284\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__9279\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__2050\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9269\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9269\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9266\,
            I => \N__9260\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9265\,
            I => \N__9260\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__9260\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9253\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9256\,
            I => \N__9250\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__9253\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9250\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9241\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9238\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__9241\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__9238\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__9233\,
            I => \U409_TRANSFER_ACK.N_7_cascade_\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9230\,
            I => \N__9227\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9227\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_3\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9221\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9221\,
            I => \N__9218\
        );

    \I__2032\ : Span4Mux_v
    port map (
            O => \N__9218\,
            I => \N__9215\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__9215\,
            I => \AC_TACK\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9212\,
            I => \N__9208\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9211\,
            I => \N__9205\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9208\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__9205\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__9197\,
            I => \U409_TRANSFER_ACK.TACK_START_2_1\
        );

    \I__2024\ : InMux
    port map (
            O => \N__9194\,
            I => \N__9189\
        );

    \I__2023\ : CascadeMux
    port map (
            O => \N__9193\,
            I => \N__9186\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__9192\,
            I => \N__9182\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9189\,
            I => \N__9179\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9186\,
            I => \N__9174\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9174\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9171\
        );

    \I__2017\ : Span4Mux_v
    port map (
            O => \N__9179\,
            I => \N__9166\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9174\,
            I => \N__9166\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9171\,
            I => \U409_TRANSFER_ACK.TACK_STARTZ0\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__9166\,
            I => \U409_TRANSFER_ACK.TACK_STARTZ0\
        );

    \I__2013\ : ClkMux
    port map (
            O => \N__9161\,
            I => \N__9134\
        );

    \I__2012\ : ClkMux
    port map (
            O => \N__9160\,
            I => \N__9134\
        );

    \I__2011\ : ClkMux
    port map (
            O => \N__9159\,
            I => \N__9134\
        );

    \I__2010\ : ClkMux
    port map (
            O => \N__9158\,
            I => \N__9134\
        );

    \I__2009\ : ClkMux
    port map (
            O => \N__9157\,
            I => \N__9134\
        );

    \I__2008\ : ClkMux
    port map (
            O => \N__9156\,
            I => \N__9134\
        );

    \I__2007\ : ClkMux
    port map (
            O => \N__9155\,
            I => \N__9134\
        );

    \I__2006\ : ClkMux
    port map (
            O => \N__9154\,
            I => \N__9134\
        );

    \I__2005\ : ClkMux
    port map (
            O => \N__9153\,
            I => \N__9134\
        );

    \I__2004\ : GlobalMux
    port map (
            O => \N__9134\,
            I => \CLK80_OUT\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9128\,
            I => \N__9125\
        );

    \I__2001\ : Odrv4
    port map (
            O => \N__9125\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_0\
        );

    \I__2000\ : IoInMux
    port map (
            O => \N__9122\,
            I => \N__9118\
        );

    \I__1999\ : IoInMux
    port map (
            O => \N__9121\,
            I => \N__9115\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__9118\,
            I => \N__9112\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__9115\,
            I => \N__9109\
        );

    \I__1996\ : IoSpan4Mux
    port map (
            O => \N__9112\,
            I => \N__9103\
        );

    \I__1995\ : IoSpan4Mux
    port map (
            O => \N__9109\,
            I => \N__9103\
        );

    \I__1994\ : IoInMux
    port map (
            O => \N__9108\,
            I => \N__9100\
        );

    \I__1993\ : Span4Mux_s3_v
    port map (
            O => \N__9103\,
            I => \N__9097\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__9100\,
            I => \N__9093\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__9097\,
            I => \N__9090\
        );

    \I__1990\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9087\
        );

    \I__1989\ : Span12Mux_s7_v
    port map (
            O => \N__9093\,
            I => \N__9082\
        );

    \I__1988\ : Sp12to4
    port map (
            O => \N__9090\,
            I => \N__9082\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__9087\,
            I => \N__9079\
        );

    \I__1986\ : Span12Mux_h
    port map (
            O => \N__9082\,
            I => \N__9075\
        );

    \I__1985\ : Span4Mux_v
    port map (
            O => \N__9079\,
            I => \N__9072\
        );

    \I__1984\ : InMux
    port map (
            O => \N__9078\,
            I => \N__9069\
        );

    \I__1983\ : Odrv12
    port map (
            O => \N__9075\,
            I => \TACK_EN\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__9072\,
            I => \TACK_EN\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__9069\,
            I => \TACK_EN\
        );

    \I__1980\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__9059\,
            I => \N__9055\
        );

    \I__1978\ : InMux
    port map (
            O => \N__9058\,
            I => \N__9052\
        );

    \I__1977\ : Span4Mux_v
    port map (
            O => \N__9055\,
            I => \N__9049\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__9052\,
            I => \N__9042\
        );

    \I__1975\ : Span4Mux_h
    port map (
            O => \N__9049\,
            I => \N__9037\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__9048\,
            I => \N__9031\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__9047\,
            I => \N__9028\
        );

    \I__1972\ : InMux
    port map (
            O => \N__9046\,
            I => \N__9016\
        );

    \I__1971\ : InMux
    port map (
            O => \N__9045\,
            I => \N__9016\
        );

    \I__1970\ : Span4Mux_v
    port map (
            O => \N__9042\,
            I => \N__9013\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9041\,
            I => \N__9008\
        );

    \I__1968\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9008\
        );

    \I__1967\ : Span4Mux_h
    port map (
            O => \N__9037\,
            I => \N__9004\
        );

    \I__1966\ : InMux
    port map (
            O => \N__9036\,
            I => \N__9001\
        );

    \I__1965\ : InMux
    port map (
            O => \N__9035\,
            I => \N__8998\
        );

    \I__1964\ : InMux
    port map (
            O => \N__9034\,
            I => \N__8985\
        );

    \I__1963\ : InMux
    port map (
            O => \N__9031\,
            I => \N__8985\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9028\,
            I => \N__8985\
        );

    \I__1961\ : InMux
    port map (
            O => \N__9027\,
            I => \N__8985\
        );

    \I__1960\ : InMux
    port map (
            O => \N__9026\,
            I => \N__8985\
        );

    \I__1959\ : InMux
    port map (
            O => \N__9025\,
            I => \N__8985\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__9024\,
            I => \N__8980\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__9023\,
            I => \N__8977\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__9022\,
            I => \N__8973\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__9021\,
            I => \N__8970\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__9016\,
            I => \N__8966\
        );

    \I__1953\ : Span4Mux_v
    port map (
            O => \N__9013\,
            I => \N__8961\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__9008\,
            I => \N__8961\
        );

    \I__1951\ : InMux
    port map (
            O => \N__9007\,
            I => \N__8958\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__9004\,
            I => \N__8949\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__9001\,
            I => \N__8949\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__8998\,
            I => \N__8949\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8985\,
            I => \N__8949\
        );

    \I__1946\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8945\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8983\,
            I => \N__8940\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8980\,
            I => \N__8940\
        );

    \I__1943\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8937\
        );

    \I__1942\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8934\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8973\,
            I => \N__8929\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8929\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8969\,
            I => \N__8925\
        );

    \I__1938\ : Span4Mux_h
    port map (
            O => \N__8966\,
            I => \N__8918\
        );

    \I__1937\ : Span4Mux_h
    port map (
            O => \N__8961\,
            I => \N__8918\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8958\,
            I => \N__8918\
        );

    \I__1935\ : Span4Mux_v
    port map (
            O => \N__8949\,
            I => \N__8915\
        );

    \I__1934\ : InMux
    port map (
            O => \N__8948\,
            I => \N__8912\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__8945\,
            I => \N__8901\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__8940\,
            I => \N__8901\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__8937\,
            I => \N__8901\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__8934\,
            I => \N__8901\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__8929\,
            I => \N__8901\
        );

    \I__1928\ : InMux
    port map (
            O => \N__8928\,
            I => \N__8898\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__8925\,
            I => \N__8895\
        );

    \I__1926\ : Span4Mux_v
    port map (
            O => \N__8918\,
            I => \N__8892\
        );

    \I__1925\ : Span4Mux_h
    port map (
            O => \N__8915\,
            I => \N__8887\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8912\,
            I => \N__8887\
        );

    \I__1923\ : Span4Mux_v
    port map (
            O => \N__8901\,
            I => \N__8882\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__8898\,
            I => \N__8882\
        );

    \I__1921\ : Span12Mux_v
    port map (
            O => \N__8895\,
            I => \N__8879\
        );

    \I__1920\ : Sp12to4
    port map (
            O => \N__8892\,
            I => \N__8876\
        );

    \I__1919\ : Span4Mux_v
    port map (
            O => \N__8887\,
            I => \N__8871\
        );

    \I__1918\ : Span4Mux_v
    port map (
            O => \N__8882\,
            I => \N__8871\
        );

    \I__1917\ : Span12Mux_v
    port map (
            O => \N__8879\,
            I => \N__8868\
        );

    \I__1916\ : Span12Mux_h
    port map (
            O => \N__8876\,
            I => \N__8865\
        );

    \I__1915\ : Sp12to4
    port map (
            O => \N__8871\,
            I => \N__8862\
        );

    \I__1914\ : Span12Mux_h
    port map (
            O => \N__8868\,
            I => \N__8857\
        );

    \I__1913\ : Span12Mux_v
    port map (
            O => \N__8865\,
            I => \N__8857\
        );

    \I__1912\ : Span12Mux_h
    port map (
            O => \N__8862\,
            I => \N__8854\
        );

    \I__1911\ : Odrv12
    port map (
            O => \N__8857\,
            I => \RESETn_c\
        );

    \I__1910\ : Odrv12
    port map (
            O => \N__8854\,
            I => \RESETn_c\
        );

    \I__1909\ : SRMux
    port map (
            O => \N__8849\,
            I => \N__8846\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8846\,
            I => \N__8843\
        );

    \I__1907\ : Span4Mux_v
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__1906\ : Span4Mux_v
    port map (
            O => \N__8840\,
            I => \N__8837\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__8837\,
            I => \U409_TRANSFER_ACK.TACK_RST_0_i\
        );

    \I__1904\ : InMux
    port map (
            O => \N__8834\,
            I => \N__8829\
        );

    \I__1903\ : InMux
    port map (
            O => \N__8833\,
            I => \N__8825\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8822\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__8829\,
            I => \N__8819\
        );

    \I__1900\ : InMux
    port map (
            O => \N__8828\,
            I => \N__8816\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__8825\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__8822\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1897\ : Odrv12
    port map (
            O => \N__8819\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__8816\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8803\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__8806\,
            I => \N__8796\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__8803\,
            I => \N__8793\
        );

    \I__1892\ : InMux
    port map (
            O => \N__8802\,
            I => \N__8788\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8801\,
            I => \N__8788\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8783\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8799\,
            I => \N__8783\
        );

    \I__1888\ : InMux
    port map (
            O => \N__8796\,
            I => \N__8780\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__8793\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__8788\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8783\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__8780\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__8771\,
            I => \N__8768\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8764\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8767\,
            I => \N__8759\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8764\,
            I => \N__8756\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8753\
        );

    \I__1878\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8750\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8759\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__8756\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8753\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__8750\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8738\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8738\,
            I => \N__8731\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8737\,
            I => \N__8723\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8736\,
            I => \N__8723\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8735\,
            I => \N__8723\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8734\,
            I => \N__8720\
        );

    \I__1867\ : Span4Mux_v
    port map (
            O => \N__8731\,
            I => \N__8717\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8730\,
            I => \N__8714\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8723\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8720\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__8717\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8714\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__8705\,
            I => \U409_CIA.CLK_CIA6_3_cascade_\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8697\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__8701\,
            I => \N__8692\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__8700\,
            I => \N__8689\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__8697\,
            I => \N__8686\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8696\,
            I => \N__8683\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8695\,
            I => \N__8678\
        );

    \I__1854\ : InMux
    port map (
            O => \N__8692\,
            I => \N__8678\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8689\,
            I => \N__8675\
        );

    \I__1852\ : Odrv12
    port map (
            O => \N__8686\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8683\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8678\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8675\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8662\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__8665\,
            I => \N__8658\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__8662\,
            I => \N__8654\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8661\,
            I => \N__8651\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8658\,
            I => \N__8648\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8657\,
            I => \N__8645\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__8654\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8651\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8648\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8645\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8636\,
            I => \N__8633\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8633\,
            I => \N__8626\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8632\,
            I => \N__8623\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8631\,
            I => \N__8620\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8615\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8629\,
            I => \N__8615\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__8626\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8623\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8620\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__8615\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8606\,
            I => \N__8603\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8603\,
            I => \N__8597\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8602\,
            I => \N__8594\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8601\,
            I => \N__8591\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8600\,
            I => \N__8588\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__8597\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8594\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8591\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8588\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8576\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__8576\,
            I => \U409_CIA.CLK_CIA_r_1_0\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__8573\,
            I => \N__8569\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__8572\,
            I => \N__8565\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8562\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8559\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8565\,
            I => \N__8556\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8562\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__8559\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8556\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8546\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8546\,
            I => \N__8541\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8545\,
            I => \N__8538\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8535\
        );

    \I__1805\ : Odrv4
    port map (
            O => \N__8541\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8538\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8535\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1802\ : InMux
    port map (
            O => \N__8528\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_0\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8525\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_1\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8522\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_2\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8516\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8516\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_2\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8510\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8510\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_1\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8507\,
            I => \N__8503\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8506\,
            I => \N__8500\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8503\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__8500\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8491\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8494\,
            I => \N__8488\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8491\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8488\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8480\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8480\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_2\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8471\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8476\,
            I => \N__8471\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8471\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__8468\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_cascade_\
        );

    \I__1781\ : IoInMux
    port map (
            O => \N__8465\,
            I => \N__8462\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8462\,
            I => \N__8459\
        );

    \I__1779\ : Odrv12
    port map (
            O => \N__8459\,
            I => \RESETn_c_i\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8452\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__8455\,
            I => \N__8448\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8452\,
            I => \N__8445\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8451\,
            I => \N__8442\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8448\,
            I => \N__8439\
        );

    \I__1773\ : Span4Mux_v
    port map (
            O => \N__8445\,
            I => \N__8436\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8442\,
            I => \N__8431\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__8439\,
            I => \N__8431\
        );

    \I__1770\ : Span4Mux_h
    port map (
            O => \N__8436\,
            I => \N__8428\
        );

    \I__1769\ : Span4Mux_v
    port map (
            O => \N__8431\,
            I => \N__8425\
        );

    \I__1768\ : Sp12to4
    port map (
            O => \N__8428\,
            I => \N__8420\
        );

    \I__1767\ : Sp12to4
    port map (
            O => \N__8425\,
            I => \N__8420\
        );

    \I__1766\ : Odrv12
    port map (
            O => \N__8420\,
            I => \A_c_12\
        );

    \I__1765\ : IoInMux
    port map (
            O => \N__8417\,
            I => \N__8414\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8414\,
            I => \N__8411\
        );

    \I__1763\ : IoSpan4Mux
    port map (
            O => \N__8411\,
            I => \N__8408\
        );

    \I__1762\ : IoSpan4Mux
    port map (
            O => \N__8408\,
            I => \N__8405\
        );

    \I__1761\ : Sp12to4
    port map (
            O => \N__8405\,
            I => \N__8402\
        );

    \I__1760\ : Span12Mux_s7_h
    port map (
            O => \N__8402\,
            I => \N__8399\
        );

    \I__1759\ : Odrv12
    port map (
            O => \N__8399\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8396\,
            I => \N__8392\
        );

    \I__1757\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8389\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8392\,
            I => \CIA_ENABLE\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__8389\,
            I => \CIA_ENABLE\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8384\,
            I => \N__8380\
        );

    \I__1753\ : CascadeMux
    port map (
            O => \N__8383\,
            I => \N__8376\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8380\,
            I => \N__8373\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8379\,
            I => \N__8370\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8367\
        );

    \I__1749\ : Sp12to4
    port map (
            O => \N__8373\,
            I => \N__8364\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8370\,
            I => \N__8359\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8367\,
            I => \N__8359\
        );

    \I__1746\ : Span12Mux_v
    port map (
            O => \N__8364\,
            I => \N__8356\
        );

    \I__1745\ : Span4Mux_v
    port map (
            O => \N__8359\,
            I => \N__8353\
        );

    \I__1744\ : Span12Mux_h
    port map (
            O => \N__8356\,
            I => \N__8350\
        );

    \I__1743\ : Sp12to4
    port map (
            O => \N__8353\,
            I => \N__8347\
        );

    \I__1742\ : Odrv12
    port map (
            O => \N__8350\,
            I => \A_c_13\
        );

    \I__1741\ : Odrv12
    port map (
            O => \N__8347\,
            I => \A_c_13\
        );

    \I__1740\ : IoInMux
    port map (
            O => \N__8342\,
            I => \N__8339\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8339\,
            I => \N__8336\
        );

    \I__1738\ : IoSpan4Mux
    port map (
            O => \N__8336\,
            I => \N__8333\
        );

    \I__1737\ : Span4Mux_s1_h
    port map (
            O => \N__8333\,
            I => \N__8330\
        );

    \I__1736\ : Sp12to4
    port map (
            O => \N__8330\,
            I => \N__8327\
        );

    \I__1735\ : Span12Mux_h
    port map (
            O => \N__8327\,
            I => \N__8324\
        );

    \I__1734\ : Odrv12
    port map (
            O => \N__8324\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8318\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8318\,
            I => \U409_TRANSFER_ACK.N_5_0\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8315\,
            I => \N__8304\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8314\,
            I => \N__8304\
        );

    \I__1729\ : InMux
    port map (
            O => \N__8313\,
            I => \N__8304\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8312\,
            I => \N__8301\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8311\,
            I => \N__8298\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__8304\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8301\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8298\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8291\,
            I => \N__8285\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8282\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8289\,
            I => \N__8277\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8288\,
            I => \N__8277\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8285\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__8282\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8277\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__8270\,
            I => \N__8264\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8269\,
            I => \N__8261\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8268\,
            I => \N__8258\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8267\,
            I => \N__8253\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8264\,
            I => \N__8253\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8261\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8258\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__8253\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8246\,
            I => \N__8241\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8236\
        );

    \I__1706\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8236\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__8241\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__8236\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__8231\,
            I => \N__8225\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8220\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8229\,
            I => \N__8220\
        );

    \I__1700\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8215\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8225\,
            I => \N__8215\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__8220\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8215\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__8210\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\
        );

    \I__1695\ : InMux
    port map (
            O => \N__8207\,
            I => \N__8200\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8191\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8191\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8204\,
            I => \N__8191\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8203\,
            I => \N__8191\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__8200\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8191\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__8186\,
            I => \N__8181\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8185\,
            I => \N__8177\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8184\,
            I => \N__8170\
        );

    \I__1685\ : InMux
    port map (
            O => \N__8181\,
            I => \N__8170\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8180\,
            I => \N__8170\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8177\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__8170\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1681\ : InMux
    port map (
            O => \N__8165\,
            I => \N__8159\
        );

    \I__1680\ : InMux
    port map (
            O => \N__8164\,
            I => \N__8159\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8159\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__8156\,
            I => \N__8152\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8149\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8146\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__8149\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8146\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8141\,
            I => \N__8134\
        );

    \I__1672\ : InMux
    port map (
            O => \N__8140\,
            I => \N__8134\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8131\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8134\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8131\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__1668\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8121\
        );

    \I__1667\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8114\
        );

    \I__1666\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8111\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8121\,
            I => \N__8108\
        );

    \I__1664\ : InMux
    port map (
            O => \N__8120\,
            I => \N__8099\
        );

    \I__1663\ : InMux
    port map (
            O => \N__8119\,
            I => \N__8099\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8099\
        );

    \I__1661\ : InMux
    port map (
            O => \N__8117\,
            I => \N__8099\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__8114\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__8111\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__8108\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__8099\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1656\ : SRMux
    port map (
            O => \N__8090\,
            I => \N__8087\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__8087\,
            I => \N__8082\
        );

    \I__1654\ : SRMux
    port map (
            O => \N__8086\,
            I => \N__8079\
        );

    \I__1653\ : SRMux
    port map (
            O => \N__8085\,
            I => \N__8076\
        );

    \I__1652\ : Span4Mux_h
    port map (
            O => \N__8082\,
            I => \N__8073\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8079\,
            I => \N__8070\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__8076\,
            I => \N__8067\
        );

    \I__1649\ : Span4Mux_h
    port map (
            O => \N__8073\,
            I => \N__8062\
        );

    \I__1648\ : Span4Mux_h
    port map (
            O => \N__8070\,
            I => \N__8062\
        );

    \I__1647\ : Span4Mux_v
    port map (
            O => \N__8067\,
            I => \N__8059\
        );

    \I__1646\ : Odrv4
    port map (
            O => \N__8062\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1645\ : Odrv4
    port map (
            O => \N__8059\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1644\ : InMux
    port map (
            O => \N__8054\,
            I => \N__8051\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__8051\,
            I => \N__8048\
        );

    \I__1642\ : Span4Mux_v
    port map (
            O => \N__8048\,
            I => \N__8044\
        );

    \I__1641\ : InMux
    port map (
            O => \N__8047\,
            I => \N__8041\
        );

    \I__1640\ : Span4Mux_h
    port map (
            O => \N__8044\,
            I => \N__8036\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__8041\,
            I => \N__8036\
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__8036\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__8033\,
            I => \N__8030\
        );

    \I__1636\ : InMux
    port map (
            O => \N__8030\,
            I => \N__8027\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__8027\,
            I => \N__8024\
        );

    \I__1634\ : Span4Mux_v
    port map (
            O => \N__8024\,
            I => \N__8021\
        );

    \I__1633\ : Span4Mux_v
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1632\ : Span4Mux_v
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__1631\ : Span4Mux_h
    port map (
            O => \N__8015\,
            I => \N__8012\
        );

    \I__1630\ : Odrv4
    port map (
            O => \N__8012\,
            I => \U409_ADDRESS_DECODE_AUTOVECTOR_10\
        );

    \I__1629\ : InMux
    port map (
            O => \N__8009\,
            I => \N__8004\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8008\,
            I => \N__8001\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8007\,
            I => \N__7998\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__8004\,
            I => \N__7994\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__8001\,
            I => \N__7991\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7998\,
            I => \N__7988\
        );

    \I__1623\ : InMux
    port map (
            O => \N__7997\,
            I => \N__7984\
        );

    \I__1622\ : Span4Mux_v
    port map (
            O => \N__7994\,
            I => \N__7981\
        );

    \I__1621\ : Span4Mux_v
    port map (
            O => \N__7991\,
            I => \N__7976\
        );

    \I__1620\ : Span4Mux_v
    port map (
            O => \N__7988\,
            I => \N__7976\
        );

    \I__1619\ : InMux
    port map (
            O => \N__7987\,
            I => \N__7973\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__7984\,
            I => \N__7964\
        );

    \I__1617\ : Sp12to4
    port map (
            O => \N__7981\,
            I => \N__7964\
        );

    \I__1616\ : Sp12to4
    port map (
            O => \N__7976\,
            I => \N__7964\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__7973\,
            I => \N__7964\
        );

    \I__1614\ : Span12Mux_h
    port map (
            O => \N__7964\,
            I => \N__7961\
        );

    \I__1613\ : Span12Mux_v
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__1612\ : Odrv12
    port map (
            O => \N__7958\,
            I => \TSn_c\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__7955\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_2_cascade_\
        );

    \I__1610\ : InMux
    port map (
            O => \N__7952\,
            I => \N__7949\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__7949\,
            I => \N__7943\
        );

    \I__1608\ : InMux
    port map (
            O => \N__7948\,
            I => \N__7938\
        );

    \I__1607\ : InMux
    port map (
            O => \N__7947\,
            I => \N__7938\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7935\
        );

    \I__1605\ : Odrv12
    port map (
            O => \N__7943\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_5\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__7938\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_5\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__7935\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_5\
        );

    \I__1602\ : InMux
    port map (
            O => \N__7928\,
            I => \N__7925\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__7925\,
            I => \N__7922\
        );

    \I__1600\ : Odrv12
    port map (
            O => \N__7922\,
            I => \U409_ADDRESS_DECODE.AUTOVECTOR_4Z0Z_0\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7916\,
            I => \N__7913\
        );

    \I__1597\ : Span4Mux_v
    port map (
            O => \N__7913\,
            I => \N__7910\
        );

    \I__1596\ : Span4Mux_v
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__1595\ : Sp12to4
    port map (
            O => \N__7907\,
            I => \N__7904\
        );

    \I__1594\ : Odrv12
    port map (
            O => \N__7904\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7901\,
            I => \N__7898\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__7898\,
            I => \U409_ADDRESS_DECODE_AUTOVECTOR_11\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7892\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__7892\,
            I => \U409_CIA.CLK_CIA6_4\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__7889\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__7883\,
            I => \N__7880\
        );

    \I__1586\ : Span4Mux_v
    port map (
            O => \N__7880\,
            I => \N__7877\
        );

    \I__1585\ : Span4Mux_h
    port map (
            O => \N__7877\,
            I => \N__7873\
        );

    \I__1584\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7870\
        );

    \I__1583\ : Odrv4
    port map (
            O => \N__7873\,
            I => \CIA_SPACE\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7870\,
            I => \CIA_SPACE\
        );

    \I__1581\ : CascadeMux
    port map (
            O => \N__7865\,
            I => \U409_CIA.VMA_RNOZ0Z_0_cascade_\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7862\,
            I => \N__7853\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7861\,
            I => \N__7853\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7860\,
            I => \N__7853\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7853\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__7850\,
            I => \N__7844\
        );

    \I__1575\ : InMux
    port map (
            O => \N__7849\,
            I => \N__7840\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7848\,
            I => \N__7833\
        );

    \I__1573\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7833\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7833\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7843\,
            I => \N__7830\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7840\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7833\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7830\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__7823\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\
        );

    \I__1566\ : InMux
    port map (
            O => \N__7820\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7817\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7814\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7808\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__7808\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7805\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7802\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\
        );

    \I__1559\ : InMux
    port map (
            O => \N__7799\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\
        );

    \I__1558\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7793\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7793\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__7790\,
            I => \N__7787\
        );

    \I__1555\ : InMux
    port map (
            O => \N__7787\,
            I => \N__7783\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7786\,
            I => \N__7780\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__7783\,
            I => \U409_CIA.CIA_CLK_COUNT11_3\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7780\,
            I => \U409_CIA.CIA_CLK_COUNT11_3\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7772\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7772\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__7769\,
            I => \N__7766\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7766\,
            I => \N__7763\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7763\,
            I => \U409_TRANSFER_ACK.TACK_EN8\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7760\,
            I => \N__7757\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7757\,
            I => \U409_TRANSFER_ACK.TACK_STATE_ns_1_0\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7754\,
            I => \N__7748\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7743\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7752\,
            I => \N__7743\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7751\,
            I => \N__7740\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7748\,
            I => \U409_TRANSFER_ACK.TACK_STATEZ0Z_0\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7743\,
            I => \U409_TRANSFER_ACK.TACK_STATEZ0Z_0\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7740\,
            I => \U409_TRANSFER_ACK.TACK_STATEZ0Z_0\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__7733\,
            I => \N__7728\
        );

    \I__1536\ : InMux
    port map (
            O => \N__7732\,
            I => \N__7721\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7731\,
            I => \N__7721\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7728\,
            I => \N__7721\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7721\,
            I => \U409_TRANSFER_ACK.TACK_STATEZ0Z_1\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7718\,
            I => \N__7714\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7711\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7714\,
            I => \N__7705\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__7711\,
            I => \N__7705\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7700\
        );

    \I__1527\ : Span4Mux_v
    port map (
            O => \N__7705\,
            I => \N__7697\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7704\,
            I => \N__7694\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7691\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7700\,
            I => \N__7687\
        );

    \I__1523\ : Span4Mux_h
    port map (
            O => \N__7697\,
            I => \N__7680\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7694\,
            I => \N__7680\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7691\,
            I => \N__7680\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7690\,
            I => \N__7677\
        );

    \I__1519\ : Span4Mux_v
    port map (
            O => \N__7687\,
            I => \N__7674\
        );

    \I__1518\ : Span4Mux_h
    port map (
            O => \N__7680\,
            I => \N__7671\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__7677\,
            I => \N__7668\
        );

    \I__1516\ : Span4Mux_v
    port map (
            O => \N__7674\,
            I => \N__7665\
        );

    \I__1515\ : Span4Mux_v
    port map (
            O => \N__7671\,
            I => \N__7662\
        );

    \I__1514\ : Span12Mux_h
    port map (
            O => \N__7668\,
            I => \N__7659\
        );

    \I__1513\ : Span4Mux_v
    port map (
            O => \N__7665\,
            I => \N__7656\
        );

    \I__1512\ : Span4Mux_v
    port map (
            O => \N__7662\,
            I => \N__7653\
        );

    \I__1511\ : Odrv12
    port map (
            O => \N__7659\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__1510\ : Odrv4
    port map (
            O => \N__7656\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__1509\ : Odrv4
    port map (
            O => \N__7653\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__7646\,
            I => \N__7642\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7645\,
            I => \N__7639\
        );

    \I__1506\ : InMux
    port map (
            O => \N__7642\,
            I => \N__7636\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7639\,
            I => \N__7631\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7636\,
            I => \N__7631\
        );

    \I__1503\ : Span4Mux_v
    port map (
            O => \N__7631\,
            I => \N__7628\
        );

    \I__1502\ : Span4Mux_h
    port map (
            O => \N__7628\,
            I => \N__7625\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__7625\,
            I => \U409_ADDRESS_DECODE_HIROM\
        );

    \I__1500\ : IoInMux
    port map (
            O => \N__7622\,
            I => \N__7619\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__7619\,
            I => \N__7616\
        );

    \I__1498\ : IoSpan4Mux
    port map (
            O => \N__7616\,
            I => \N__7612\
        );

    \I__1497\ : IoInMux
    port map (
            O => \N__7615\,
            I => \N__7609\
        );

    \I__1496\ : Span4Mux_s2_v
    port map (
            O => \N__7612\,
            I => \N__7606\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7609\,
            I => \N__7602\
        );

    \I__1494\ : Span4Mux_v
    port map (
            O => \N__7606\,
            I => \N__7599\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__7605\,
            I => \N__7596\
        );

    \I__1492\ : Span12Mux_s8_v
    port map (
            O => \N__7602\,
            I => \N__7593\
        );

    \I__1491\ : Sp12to4
    port map (
            O => \N__7599\,
            I => \N__7590\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7596\,
            I => \N__7587\
        );

    \I__1489\ : Span12Mux_h
    port map (
            O => \N__7593\,
            I => \N__7583\
        );

    \I__1488\ : Span12Mux_v
    port map (
            O => \N__7590\,
            I => \N__7580\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7587\,
            I => \N__7577\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7586\,
            I => \N__7574\
        );

    \I__1485\ : Odrv12
    port map (
            O => \N__7583\,
            I => \TACK_OUT\
        );

    \I__1484\ : Odrv12
    port map (
            O => \N__7580\,
            I => \TACK_OUT\
        );

    \I__1483\ : Odrv4
    port map (
            O => \N__7577\,
            I => \TACK_OUT\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7574\,
            I => \TACK_OUT\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7562\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7562\,
            I => \N__7558\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7561\,
            I => \N__7555\
        );

    \I__1478\ : Span4Mux_h
    port map (
            O => \N__7558\,
            I => \N__7552\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__7555\,
            I => \N__7549\
        );

    \I__1476\ : Odrv4
    port map (
            O => \N__7552\,
            I => \U409_ADDRESS_DECODE_LOWROM\
        );

    \I__1475\ : Odrv12
    port map (
            O => \N__7549\,
            I => \U409_ADDRESS_DECODE_LOWROM\
        );

    \I__1474\ : IoInMux
    port map (
            O => \N__7544\,
            I => \N__7541\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7541\,
            I => \N__7538\
        );

    \I__1472\ : Span4Mux_s2_v
    port map (
            O => \N__7538\,
            I => \N__7535\
        );

    \I__1471\ : Sp12to4
    port map (
            O => \N__7535\,
            I => \N__7532\
        );

    \I__1470\ : Span12Mux_h
    port map (
            O => \N__7532\,
            I => \N__7529\
        );

    \I__1469\ : Span12Mux_v
    port map (
            O => \N__7529\,
            I => \N__7526\
        );

    \I__1468\ : Odrv12
    port map (
            O => \N__7526\,
            I => \U409_TRANSFER_ACK_un1_TACK_OUT_0_i\
        );

    \I__1467\ : IoInMux
    port map (
            O => \N__7523\,
            I => \N__7520\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7520\,
            I => \N__7517\
        );

    \I__1465\ : Span4Mux_s2_v
    port map (
            O => \N__7517\,
            I => \N__7514\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__7514\,
            I => \N__7511\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__7511\,
            I => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__7508\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__7505\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__7502\,
            I => \N__7499\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7499\,
            I => \N__7496\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7496\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__7493\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__7490\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7487\,
            I => \N__7481\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7486\,
            I => \N__7481\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7481\,
            I => \N__7478\
        );

    \I__1452\ : Span4Mux_v
    port map (
            O => \N__7478\,
            I => \N__7474\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7477\,
            I => \N__7471\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__7474\,
            I => \U409_AUTOCONFIG.N_78\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7471\,
            I => \U409_AUTOCONFIG.N_78\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7460\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7465\,
            I => \N__7460\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7460\,
            I => \N__7457\
        );

    \I__1445\ : Odrv12
    port map (
            O => \N__7457\,
            I => \U409_AUTOCONFIG.N_92\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7454\,
            I => \N__7451\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7451\,
            I => \N__7448\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__7448\,
            I => \U409_AUTOCONFIG.PR_OUTZ0Z_0\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7445\,
            I => \N__7442\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__7442\,
            I => \N__7439\
        );

    \I__1439\ : Odrv12
    port map (
            O => \N__7439\,
            I => \U409_AUTOCONFIG.LIDE_OUT_7_i_a3_1_0\
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__7436\,
            I => \N__7433\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7433\,
            I => \N__7430\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7430\,
            I => \N__7427\
        );

    \I__1435\ : Span12Mux_h
    port map (
            O => \N__7427\,
            I => \N__7424\
        );

    \I__1434\ : Odrv12
    port map (
            O => \N__7424\,
            I => \U409_AUTOCONFIG.LIDE_OUT_7_i_a3_0_0\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7421\,
            I => \N__7418\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7418\,
            I => \N__7415\
        );

    \I__1431\ : Odrv12
    port map (
            O => \N__7415\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\
        );

    \I__1430\ : CEMux
    port map (
            O => \N__7412\,
            I => \N__7408\
        );

    \I__1429\ : CEMux
    port map (
            O => \N__7411\,
            I => \N__7403\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__7408\,
            I => \N__7400\
        );

    \I__1427\ : CEMux
    port map (
            O => \N__7407\,
            I => \N__7397\
        );

    \I__1426\ : CEMux
    port map (
            O => \N__7406\,
            I => \N__7394\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7403\,
            I => \N__7391\
        );

    \I__1424\ : Span4Mux_v
    port map (
            O => \N__7400\,
            I => \N__7385\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__7397\,
            I => \N__7385\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7394\,
            I => \N__7382\
        );

    \I__1421\ : Span4Mux_v
    port map (
            O => \N__7391\,
            I => \N__7379\
        );

    \I__1420\ : CEMux
    port map (
            O => \N__7390\,
            I => \N__7376\
        );

    \I__1419\ : Span4Mux_v
    port map (
            O => \N__7385\,
            I => \N__7371\
        );

    \I__1418\ : Span4Mux_v
    port map (
            O => \N__7382\,
            I => \N__7371\
        );

    \I__1417\ : Span4Mux_h
    port map (
            O => \N__7379\,
            I => \N__7368\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7376\,
            I => \N__7365\
        );

    \I__1415\ : Span4Mux_h
    port map (
            O => \N__7371\,
            I => \N__7362\
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__7368\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\
        );

    \I__1413\ : Odrv12
    port map (
            O => \N__7365\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\
        );

    \I__1412\ : Odrv4
    port map (
            O => \N__7362\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7355\,
            I => \N__7352\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__7352\,
            I => \N__7348\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7351\,
            I => \N__7345\
        );

    \I__1408\ : Odrv4
    port map (
            O => \N__7348\,
            I => \U409_AUTOCONFIG.N_133\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7345\,
            I => \U409_AUTOCONFIG.N_133\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__7340\,
            I => \N__7334\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7339\,
            I => \N__7329\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7338\,
            I => \N__7326\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__7337\,
            I => \N__7317\
        );

    \I__1402\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7308\
        );

    \I__1401\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7308\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7305\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7329\,
            I => \N__7300\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__7326\,
            I => \N__7300\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7297\
        );

    \I__1396\ : InMux
    port map (
            O => \N__7324\,
            I => \N__7294\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7323\,
            I => \N__7291\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7288\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7321\,
            I => \N__7285\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7282\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7317\,
            I => \N__7275\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7316\,
            I => \N__7275\
        );

    \I__1389\ : InMux
    port map (
            O => \N__7315\,
            I => \N__7275\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7314\,
            I => \N__7272\
        );

    \I__1387\ : InMux
    port map (
            O => \N__7313\,
            I => \N__7269\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7308\,
            I => \N__7266\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7305\,
            I => \N__7263\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__7300\,
            I => \N__7250\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__7297\,
            I => \N__7250\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__7294\,
            I => \N__7250\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__7291\,
            I => \N__7250\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7288\,
            I => \N__7250\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__7285\,
            I => \N__7250\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__7282\,
            I => \N__7247\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7275\,
            I => \N__7240\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__7272\,
            I => \N__7240\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7269\,
            I => \N__7240\
        );

    \I__1374\ : Span4Mux_v
    port map (
            O => \N__7266\,
            I => \N__7235\
        );

    \I__1373\ : Span4Mux_v
    port map (
            O => \N__7263\,
            I => \N__7235\
        );

    \I__1372\ : Span4Mux_v
    port map (
            O => \N__7250\,
            I => \N__7232\
        );

    \I__1371\ : Span4Mux_v
    port map (
            O => \N__7247\,
            I => \N__7227\
        );

    \I__1370\ : Span4Mux_v
    port map (
            O => \N__7240\,
            I => \N__7227\
        );

    \I__1369\ : Sp12to4
    port map (
            O => \N__7235\,
            I => \N__7220\
        );

    \I__1368\ : Sp12to4
    port map (
            O => \N__7232\,
            I => \N__7220\
        );

    \I__1367\ : Sp12to4
    port map (
            O => \N__7227\,
            I => \N__7220\
        );

    \I__1366\ : Span12Mux_h
    port map (
            O => \N__7220\,
            I => \N__7217\
        );

    \I__1365\ : Span12Mux_v
    port map (
            O => \N__7217\,
            I => \N__7214\
        );

    \I__1364\ : Odrv12
    port map (
            O => \N__7214\,
            I => \A_c_1\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__7211\,
            I => \N__7208\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7208\,
            I => \N__7205\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7205\,
            I => \N__7202\
        );

    \I__1360\ : Span4Mux_v
    port map (
            O => \N__7202\,
            I => \N__7199\
        );

    \I__1359\ : Span4Mux_h
    port map (
            O => \N__7199\,
            I => \N__7196\
        );

    \I__1358\ : Sp12to4
    port map (
            O => \N__7196\,
            I => \N__7193\
        );

    \I__1357\ : Span12Mux_h
    port map (
            O => \N__7193\,
            I => \N__7190\
        );

    \I__1356\ : Span12Mux_v
    port map (
            O => \N__7190\,
            I => \N__7187\
        );

    \I__1355\ : Odrv12
    port map (
            O => \N__7187\,
            I => \AUTOBOOT_c\
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__7184\,
            I => \N__7180\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7183\,
            I => \N__7175\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7180\,
            I => \N__7175\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7175\,
            I => \N__7171\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7174\,
            I => \N__7168\
        );

    \I__1349\ : Odrv4
    port map (
            O => \N__7171\,
            I => \U409_AUTOCONFIG.N_126\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__7168\,
            I => \U409_AUTOCONFIG.N_126\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7163\,
            I => \N__7160\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7160\,
            I => \U409_AUTOCONFIG.LIDE_OUT_7_i_1_0\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7157\,
            I => \N__7154\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7154\,
            I => \N__7151\
        );

    \I__1343\ : Span12Mux_h
    port map (
            O => \N__7151\,
            I => \N__7148\
        );

    \I__1342\ : Span12Mux_v
    port map (
            O => \N__7148\,
            I => \N__7145\
        );

    \I__1341\ : Odrv12
    port map (
            O => \N__7145\,
            I => \TACKn_in\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7142\,
            I => \N__7139\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__7139\,
            I => \N__7134\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7138\,
            I => \N__7129\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7137\,
            I => \N__7129\
        );

    \I__1336\ : Odrv12
    port map (
            O => \N__7134\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__7129\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__7124\,
            I => \N__7121\
        );

    \I__1333\ : InMux
    port map (
            O => \N__7121\,
            I => \N__7118\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__7118\,
            I => \N__7114\
        );

    \I__1331\ : InMux
    port map (
            O => \N__7117\,
            I => \N__7111\
        );

    \I__1330\ : Span4Mux_v
    port map (
            O => \N__7114\,
            I => \N__7108\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__7111\,
            I => \N__7105\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__7108\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__7105\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7096\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7099\,
            I => \N__7090\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__7096\,
            I => \N__7085\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7095\,
            I => \N__7082\
        );

    \I__1322\ : InMux
    port map (
            O => \N__7094\,
            I => \N__7077\
        );

    \I__1321\ : InMux
    port map (
            O => \N__7093\,
            I => \N__7077\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__7090\,
            I => \N__7074\
        );

    \I__1319\ : InMux
    port map (
            O => \N__7089\,
            I => \N__7069\
        );

    \I__1318\ : InMux
    port map (
            O => \N__7088\,
            I => \N__7069\
        );

    \I__1317\ : Span4Mux_h
    port map (
            O => \N__7085\,
            I => \N__7064\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__7082\,
            I => \N__7064\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__7077\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__7074\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__7069\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__1312\ : Odrv4
    port map (
            O => \N__7064\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__1311\ : CEMux
    port map (
            O => \N__7055\,
            I => \N__7052\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__7052\,
            I => \N__7049\
        );

    \I__1309\ : Odrv4
    port map (
            O => \N__7049\,
            I => \U409_AUTOCONFIG.STATE_ns_0_0_1\
        );

    \I__1308\ : CascadeMux
    port map (
            O => \N__7046\,
            I => \N__7041\
        );

    \I__1307\ : InMux
    port map (
            O => \N__7045\,
            I => \N__7037\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7044\,
            I => \N__7032\
        );

    \I__1305\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7032\
        );

    \I__1304\ : InMux
    port map (
            O => \N__7040\,
            I => \N__7029\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__7037\,
            I => \U409_AUTOCONFIG.N_4\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__7032\,
            I => \U409_AUTOCONFIG.N_4\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__7029\,
            I => \U409_AUTOCONFIG.N_4\
        );

    \I__1300\ : IoInMux
    port map (
            O => \N__7022\,
            I => \N__7019\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__7019\,
            I => \N__7016\
        );

    \I__1298\ : IoSpan4Mux
    port map (
            O => \N__7016\,
            I => \N__7013\
        );

    \I__1297\ : Sp12to4
    port map (
            O => \N__7013\,
            I => \N__7010\
        );

    \I__1296\ : Span12Mux_s9_v
    port map (
            O => \N__7010\,
            I => \N__7007\
        );

    \I__1295\ : Odrv12
    port map (
            O => \N__7007\,
            I => \D_OUT_0\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7004\,
            I => \N__7001\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7001\,
            I => \N__6998\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__6998\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNI7DMPZ0Z_1\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6991\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6994\,
            I => \N__6988\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6991\,
            I => \N__6976\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6988\,
            I => \N__6976\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6987\,
            I => \N__6971\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6986\,
            I => \N__6971\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6985\,
            I => \N__6966\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6984\,
            I => \N__6966\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6983\,
            I => \N__6963\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6982\,
            I => \N__6958\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6981\,
            I => \N__6958\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__6976\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6971\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__6966\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6963\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__6958\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6947\,
            I => \N__6944\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__6944\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNI5BMPZ0Z_0\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__6941\,
            I => \N__6932\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__6940\,
            I => \N__6929\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__6939\,
            I => \N__6925\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6938\,
            I => \N__6921\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6916\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6936\,
            I => \N__6916\
        );

    \I__1267\ : CascadeMux
    port map (
            O => \N__6935\,
            I => \N__6913\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6906\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6929\,
            I => \N__6906\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6928\,
            I => \N__6906\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6903\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__6924\,
            I => \N__6899\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6921\,
            I => \N__6896\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6916\,
            I => \N__6893\
        );

    \I__1259\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6890\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__6906\,
            I => \N__6885\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6903\,
            I => \N__6885\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6902\,
            I => \N__6880\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6899\,
            I => \N__6880\
        );

    \I__1254\ : Span4Mux_v
    port map (
            O => \N__6896\,
            I => \N__6876\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__6893\,
            I => \N__6871\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6890\,
            I => \N__6871\
        );

    \I__1251\ : Span4Mux_h
    port map (
            O => \N__6885\,
            I => \N__6866\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__6880\,
            I => \N__6866\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6863\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__6876\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1247\ : Odrv4
    port map (
            O => \N__6871\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1246\ : Odrv4
    port map (
            O => \N__6866\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6863\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__6854\,
            I => \N__6849\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6853\,
            I => \N__6843\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6852\,
            I => \N__6839\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6836\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6831\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6847\,
            I => \N__6831\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6828\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6843\,
            I => \N__6825\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6822\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6839\,
            I => \CONFIGURED\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6836\,
            I => \CONFIGURED\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6831\,
            I => \CONFIGURED\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6828\,
            I => \CONFIGURED\
        );

    \I__1231\ : Odrv4
    port map (
            O => \N__6825\,
            I => \CONFIGURED\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__6822\,
            I => \CONFIGURED\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6805\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6808\,
            I => \N__6802\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6805\,
            I => \U409_AUTOCONFIG.AC_STARTZ0\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6802\,
            I => \U409_AUTOCONFIG.AC_STARTZ0\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6797\,
            I => \N__6794\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6794\,
            I => \N__6791\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__6791\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__6785\,
            I => \U409_AUTOCONFIG.N_82\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6779\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6779\,
            I => \N__6776\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__6776\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__6773\,
            I => \N__6770\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6767\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__6767\,
            I => \N__6764\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__6764\,
            I => \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0Z0Z_3\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6761\,
            I => \N__6758\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6758\,
            I => \N__6755\
        );

    \I__1211\ : Odrv12
    port map (
            O => \N__6755\,
            I => \U409_AUTOCONFIG.PR_OUTZ0Z_3\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__6752\,
            I => \N__6748\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6751\,
            I => \N__6743\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6743\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6743\,
            I => \N__6740\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__6740\,
            I => \U409_AUTOCONFIG.N_131\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6734\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6734\,
            I => \U409_AUTOCONFIG.N_93\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__6731\,
            I => \N__6728\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6725\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6725\,
            I => \N__6722\
        );

    \I__1200\ : Odrv12
    port map (
            O => \N__6722\,
            I => \U409_AUTOCONFIG.PR_OUTZ0Z_1\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6713\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6718\,
            I => \N__6713\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6713\,
            I => \N__6709\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6712\,
            I => \N__6706\
        );

    \I__1195\ : Span4Mux_v
    port map (
            O => \N__6709\,
            I => \N__6701\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__6706\,
            I => \N__6698\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6705\,
            I => \N__6693\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6704\,
            I => \N__6693\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__6701\,
            I => \U409_AUTOCONFIG.N_116\
        );

    \I__1190\ : Odrv4
    port map (
            O => \N__6698\,
            I => \U409_AUTOCONFIG.N_116\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__6693\,
            I => \U409_AUTOCONFIG.N_116\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6686\,
            I => \N__6679\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6685\,
            I => \N__6679\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6684\,
            I => \N__6676\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6679\,
            I => \N__6665\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6676\,
            I => \N__6665\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6660\
        );

    \I__1182\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6660\
        );

    \I__1181\ : CascadeMux
    port map (
            O => \N__6673\,
            I => \N__6657\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6672\,
            I => \N__6652\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6671\,
            I => \N__6649\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6670\,
            I => \N__6646\
        );

    \I__1177\ : Span4Mux_v
    port map (
            O => \N__6665\,
            I => \N__6641\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6660\,
            I => \N__6641\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6657\,
            I => \N__6636\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6636\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6655\,
            I => \N__6633\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6652\,
            I => \N__6627\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6649\,
            I => \N__6627\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6646\,
            I => \N__6620\
        );

    \I__1169\ : Span4Mux_v
    port map (
            O => \N__6641\,
            I => \N__6620\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6636\,
            I => \N__6620\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__6633\,
            I => \N__6617\
        );

    \I__1166\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6614\
        );

    \I__1165\ : Span4Mux_v
    port map (
            O => \N__6627\,
            I => \N__6611\
        );

    \I__1164\ : Span4Mux_h
    port map (
            O => \N__6620\,
            I => \N__6604\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__6617\,
            I => \N__6604\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6614\,
            I => \N__6604\
        );

    \I__1161\ : Span4Mux_v
    port map (
            O => \N__6611\,
            I => \N__6601\
        );

    \I__1160\ : Span4Mux_v
    port map (
            O => \N__6604\,
            I => \N__6598\
        );

    \I__1159\ : Sp12to4
    port map (
            O => \N__6601\,
            I => \N__6593\
        );

    \I__1158\ : Sp12to4
    port map (
            O => \N__6598\,
            I => \N__6593\
        );

    \I__1157\ : Span12Mux_h
    port map (
            O => \N__6593\,
            I => \N__6590\
        );

    \I__1156\ : Odrv12
    port map (
            O => \N__6590\,
            I => \A_c_2\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6587\,
            I => \N__6584\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6584\,
            I => \N__6581\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__6581\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6575\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__6575\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6569\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6569\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6566\,
            I => \N__6563\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6563\,
            I => \N__6560\
        );

    \I__1146\ : Odrv12
    port map (
            O => \N__6560\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6554\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6554\,
            I => \N__6550\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__6553\,
            I => \N__6547\
        );

    \I__1142\ : Span4Mux_v
    port map (
            O => \N__6550\,
            I => \N__6544\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6541\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__6544\,
            I => \U409_AUTOCONFIG.N_129\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6541\,
            I => \U409_AUTOCONFIG.N_129\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__6536\,
            I => \U409_AUTOCONFIG.N_133_cascade_\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6533\,
            I => \N__6527\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6532\,
            I => \N__6527\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6527\,
            I => \U409_AUTOCONFIG.N_127\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__6524\,
            I => \N__6521\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6521\,
            I => \N__6515\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6520\,
            I => \N__6515\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6515\,
            I => \N__6508\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6514\,
            I => \N__6505\
        );

    \I__1129\ : InMux
    port map (
            O => \N__6513\,
            I => \N__6502\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6512\,
            I => \N__6497\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6511\,
            I => \N__6497\
        );

    \I__1126\ : Span4Mux_v
    port map (
            O => \N__6508\,
            I => \N__6492\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6505\,
            I => \N__6489\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6502\,
            I => \N__6486\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6497\,
            I => \N__6483\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6480\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6495\,
            I => \N__6477\
        );

    \I__1120\ : Odrv4
    port map (
            O => \N__6492\,
            I => \U409_AUTOCONFIG.N_110\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__6489\,
            I => \U409_AUTOCONFIG.N_110\
        );

    \I__1118\ : Odrv12
    port map (
            O => \N__6486\,
            I => \U409_AUTOCONFIG.N_110\
        );

    \I__1117\ : Odrv12
    port map (
            O => \N__6483\,
            I => \U409_AUTOCONFIG.N_110\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6480\,
            I => \U409_AUTOCONFIG.N_110\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__6477\,
            I => \U409_AUTOCONFIG.N_110\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__6464\,
            I => \N__6458\
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__6463\,
            I => \N__6452\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__6462\,
            I => \N__6446\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__6461\,
            I => \N__6442\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6458\,
            I => \N__6439\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6457\,
            I => \N__6436\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6433\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6455\,
            I => \N__6428\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6452\,
            I => \N__6428\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__6451\,
            I => \N__6425\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__6450\,
            I => \N__6422\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6449\,
            I => \N__6417\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6417\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6445\,
            I => \N__6412\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6442\,
            I => \N__6412\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6439\,
            I => \N__6401\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__6436\,
            I => \N__6401\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__6433\,
            I => \N__6401\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__6428\,
            I => \N__6401\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6425\,
            I => \N__6396\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6422\,
            I => \N__6396\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6417\,
            I => \N__6391\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__6412\,
            I => \N__6391\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6386\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6410\,
            I => \N__6386\
        );

    \I__1089\ : Span4Mux_v
    port map (
            O => \N__6401\,
            I => \N__6383\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6396\,
            I => \N__6380\
        );

    \I__1087\ : Span4Mux_v
    port map (
            O => \N__6391\,
            I => \N__6375\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6386\,
            I => \N__6375\
        );

    \I__1085\ : Span4Mux_h
    port map (
            O => \N__6383\,
            I => \N__6372\
        );

    \I__1084\ : Span4Mux_v
    port map (
            O => \N__6380\,
            I => \N__6369\
        );

    \I__1083\ : Sp12to4
    port map (
            O => \N__6375\,
            I => \N__6362\
        );

    \I__1082\ : Sp12to4
    port map (
            O => \N__6372\,
            I => \N__6362\
        );

    \I__1081\ : Sp12to4
    port map (
            O => \N__6369\,
            I => \N__6362\
        );

    \I__1080\ : Odrv12
    port map (
            O => \N__6362\,
            I => \A_c_4\
        );

    \I__1079\ : IoInMux
    port map (
            O => \N__6359\,
            I => \N__6356\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6356\,
            I => \N__6353\
        );

    \I__1077\ : Span4Mux_s3_v
    port map (
            O => \N__6353\,
            I => \N__6350\
        );

    \I__1076\ : Span4Mux_v
    port map (
            O => \N__6350\,
            I => \N__6347\
        );

    \I__1075\ : Span4Mux_v
    port map (
            O => \N__6347\,
            I => \N__6344\
        );

    \I__1074\ : Odrv4
    port map (
            O => \N__6344\,
            I => \D_OUT_1\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6341\,
            I => \N__6338\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__6338\,
            I => \N__6335\
        );

    \I__1071\ : Span4Mux_v
    port map (
            O => \N__6335\,
            I => \N__6332\
        );

    \I__1070\ : Span4Mux_v
    port map (
            O => \N__6332\,
            I => \N__6329\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__6329\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3\
        );

    \I__1068\ : IoInMux
    port map (
            O => \N__6326\,
            I => \N__6323\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6323\,
            I => \N__6320\
        );

    \I__1066\ : IoSpan4Mux
    port map (
            O => \N__6320\,
            I => \N__6317\
        );

    \I__1065\ : Span4Mux_s3_v
    port map (
            O => \N__6317\,
            I => \N__6314\
        );

    \I__1064\ : Span4Mux_v
    port map (
            O => \N__6314\,
            I => \N__6311\
        );

    \I__1063\ : Odrv4
    port map (
            O => \N__6311\,
            I => \D_OUT_3\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6308\,
            I => \N__6302\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6302\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6302\,
            I => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa\
        );

    \I__1059\ : IoInMux
    port map (
            O => \N__6299\,
            I => \N__6296\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6296\,
            I => \N__6293\
        );

    \I__1057\ : Span4Mux_s0_v
    port map (
            O => \N__6293\,
            I => \N__6290\
        );

    \I__1056\ : Sp12to4
    port map (
            O => \N__6290\,
            I => \N__6287\
        );

    \I__1055\ : Span12Mux_h
    port map (
            O => \N__6287\,
            I => \N__6284\
        );

    \I__1054\ : Span12Mux_v
    port map (
            O => \N__6284\,
            I => \N__6280\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6283\,
            I => \N__6277\
        );

    \I__1052\ : Odrv12
    port map (
            O => \N__6280\,
            I => \CONFIGENn_c\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6277\,
            I => \CONFIGENn_c\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__6272\,
            I => \U409_AUTOCONFIG.STATE_ns_1_cascade_\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6263\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6260\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6257\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6266\,
            I => \N__6254\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6263\,
            I => \N__6248\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__6260\,
            I => \N__6248\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6257\,
            I => \N__6239\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6254\,
            I => \N__6239\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6253\,
            I => \N__6235\
        );

    \I__1040\ : Span4Mux_v
    port map (
            O => \N__6248\,
            I => \N__6232\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6225\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6225\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6225\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6244\,
            I => \N__6222\
        );

    \I__1035\ : Span4Mux_v
    port map (
            O => \N__6239\,
            I => \N__6219\
        );

    \I__1034\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6216\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6235\,
            I => \N__6203\
        );

    \I__1032\ : Sp12to4
    port map (
            O => \N__6232\,
            I => \N__6203\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6225\,
            I => \N__6203\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6222\,
            I => \N__6203\
        );

    \I__1029\ : Sp12to4
    port map (
            O => \N__6219\,
            I => \N__6203\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__6216\,
            I => \N__6203\
        );

    \I__1027\ : Span12Mux_h
    port map (
            O => \N__6203\,
            I => \N__6200\
        );

    \I__1026\ : Span12Mux_v
    port map (
            O => \N__6200\,
            I => \N__6197\
        );

    \I__1025\ : Odrv12
    port map (
            O => \N__6197\,
            I => \A_c_22\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6191\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6191\,
            I => \N__6188\
        );

    \I__1022\ : Odrv4
    port map (
            O => \N__6188\,
            I => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__6185\,
            I => \N__6180\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6177\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6183\,
            I => \N__6174\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6180\,
            I => \N__6171\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__6177\,
            I => \N__6166\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6166\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6171\,
            I => \N__6163\
        );

    \I__1014\ : Span4Mux_v
    port map (
            O => \N__6166\,
            I => \N__6160\
        );

    \I__1013\ : Span4Mux_v
    port map (
            O => \N__6163\,
            I => \N__6157\
        );

    \I__1012\ : Sp12to4
    port map (
            O => \N__6160\,
            I => \N__6152\
        );

    \I__1011\ : Sp12to4
    port map (
            O => \N__6157\,
            I => \N__6152\
        );

    \I__1010\ : Span12Mux_h
    port map (
            O => \N__6152\,
            I => \N__6149\
        );

    \I__1009\ : Span12Mux_v
    port map (
            O => \N__6149\,
            I => \N__6146\
        );

    \I__1008\ : Odrv12
    port map (
            O => \N__6146\,
            I => \OVL_c\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__6143\,
            I => \N__6140\
        );

    \I__1006\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6132\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6139\,
            I => \N__6128\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6138\,
            I => \N__6121\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6137\,
            I => \N__6121\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6136\,
            I => \N__6121\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__6135\,
            I => \N__6118\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__6132\,
            I => \N__6114\
        );

    \I__999\ : InMux
    port map (
            O => \N__6131\,
            I => \N__6111\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__6128\,
            I => \N__6106\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__6121\,
            I => \N__6106\
        );

    \I__996\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6101\
        );

    \I__995\ : InMux
    port map (
            O => \N__6117\,
            I => \N__6101\
        );

    \I__994\ : Span4Mux_v
    port map (
            O => \N__6114\,
            I => \N__6098\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__6111\,
            I => \N__6095\
        );

    \I__992\ : Span4Mux_h
    port map (
            O => \N__6106\,
            I => \N__6090\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__6101\,
            I => \N__6090\
        );

    \I__990\ : Span4Mux_h
    port map (
            O => \N__6098\,
            I => \N__6085\
        );

    \I__989\ : Span4Mux_v
    port map (
            O => \N__6095\,
            I => \N__6085\
        );

    \I__988\ : Span4Mux_h
    port map (
            O => \N__6090\,
            I => \N__6082\
        );

    \I__987\ : Span4Mux_v
    port map (
            O => \N__6085\,
            I => \N__6079\
        );

    \I__986\ : Span4Mux_v
    port map (
            O => \N__6082\,
            I => \N__6076\
        );

    \I__985\ : Sp12to4
    port map (
            O => \N__6079\,
            I => \N__6071\
        );

    \I__984\ : Sp12to4
    port map (
            O => \N__6076\,
            I => \N__6071\
        );

    \I__983\ : Odrv12
    port map (
            O => \N__6071\,
            I => \A_c_23\
        );

    \I__982\ : IoInMux
    port map (
            O => \N__6068\,
            I => \N__6065\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__6065\,
            I => \N__6062\
        );

    \I__980\ : Span4Mux_s3_v
    port map (
            O => \N__6062\,
            I => \N__6059\
        );

    \I__979\ : Span4Mux_h
    port map (
            O => \N__6059\,
            I => \N__6056\
        );

    \I__978\ : Sp12to4
    port map (
            O => \N__6056\,
            I => \N__6053\
        );

    \I__977\ : Odrv12
    port map (
            O => \N__6053\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\
        );

    \I__976\ : InMux
    port map (
            O => \N__6050\,
            I => \N__6044\
        );

    \I__975\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6039\
        );

    \I__974\ : InMux
    port map (
            O => \N__6048\,
            I => \N__6036\
        );

    \I__973\ : InMux
    port map (
            O => \N__6047\,
            I => \N__6033\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__6044\,
            I => \N__6030\
        );

    \I__971\ : InMux
    port map (
            O => \N__6043\,
            I => \N__6025\
        );

    \I__970\ : InMux
    port map (
            O => \N__6042\,
            I => \N__6025\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6039\,
            I => \N__6022\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__6036\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__6033\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__966\ : Odrv4
    port map (
            O => \N__6030\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__6025\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__964\ : Odrv4
    port map (
            O => \N__6022\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__963\ : InMux
    port map (
            O => \N__6011\,
            I => \N__6002\
        );

    \I__962\ : InMux
    port map (
            O => \N__6010\,
            I => \N__6002\
        );

    \I__961\ : InMux
    port map (
            O => \N__6009\,
            I => \N__6002\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__6002\,
            I => \N__5996\
        );

    \I__959\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5993\
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__6000\,
            I => \N__5990\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__5999\,
            I => \N__5986\
        );

    \I__956\ : Span4Mux_v
    port map (
            O => \N__5996\,
            I => \N__5976\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5993\,
            I => \N__5976\
        );

    \I__954\ : InMux
    port map (
            O => \N__5990\,
            I => \N__5971\
        );

    \I__953\ : InMux
    port map (
            O => \N__5989\,
            I => \N__5971\
        );

    \I__952\ : InMux
    port map (
            O => \N__5986\,
            I => \N__5968\
        );

    \I__951\ : InMux
    port map (
            O => \N__5985\,
            I => \N__5965\
        );

    \I__950\ : InMux
    port map (
            O => \N__5984\,
            I => \N__5962\
        );

    \I__949\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5959\
        );

    \I__948\ : InMux
    port map (
            O => \N__5982\,
            I => \N__5954\
        );

    \I__947\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5954\
        );

    \I__946\ : Span4Mux_h
    port map (
            O => \N__5976\,
            I => \N__5949\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5971\,
            I => \N__5949\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5968\,
            I => \N__5938\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__5965\,
            I => \N__5938\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5962\,
            I => \N__5938\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5959\,
            I => \N__5938\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5954\,
            I => \N__5938\
        );

    \I__939\ : Span4Mux_v
    port map (
            O => \N__5949\,
            I => \N__5935\
        );

    \I__938\ : Span4Mux_v
    port map (
            O => \N__5938\,
            I => \N__5932\
        );

    \I__937\ : Span4Mux_v
    port map (
            O => \N__5935\,
            I => \N__5929\
        );

    \I__936\ : Sp12to4
    port map (
            O => \N__5932\,
            I => \N__5926\
        );

    \I__935\ : Sp12to4
    port map (
            O => \N__5929\,
            I => \N__5923\
        );

    \I__934\ : Span12Mux_h
    port map (
            O => \N__5926\,
            I => \N__5920\
        );

    \I__933\ : Span12Mux_h
    port map (
            O => \N__5923\,
            I => \N__5915\
        );

    \I__932\ : Span12Mux_v
    port map (
            O => \N__5920\,
            I => \N__5915\
        );

    \I__931\ : Odrv12
    port map (
            O => \N__5915\,
            I => \RnW_c\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__5912\,
            I => \N__5909\
        );

    \I__929\ : InMux
    port map (
            O => \N__5909\,
            I => \N__5906\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5906\,
            I => \N__5902\
        );

    \I__927\ : InMux
    port map (
            O => \N__5905\,
            I => \N__5899\
        );

    \I__926\ : Span4Mux_h
    port map (
            O => \N__5902\,
            I => \N__5894\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__5899\,
            I => \N__5894\
        );

    \I__924\ : Span4Mux_v
    port map (
            O => \N__5894\,
            I => \N__5891\
        );

    \I__923\ : Sp12to4
    port map (
            O => \N__5891\,
            I => \N__5888\
        );

    \I__922\ : Span12Mux_h
    port map (
            O => \N__5888\,
            I => \N__5885\
        );

    \I__921\ : Span12Mux_v
    port map (
            O => \N__5885\,
            I => \N__5882\
        );

    \I__920\ : Odrv12
    port map (
            O => \N__5882\,
            I => \CPUCONFn_c\
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__5879\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_1_cascade_\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__5876\,
            I => \U409_AUTOCONFIG.N_227_3_cascade_\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__5873\,
            I => \N__5870\
        );

    \I__916\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5867\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__5867\,
            I => \N__5864\
        );

    \I__914\ : Span4Mux_v
    port map (
            O => \N__5864\,
            I => \N__5861\
        );

    \I__913\ : Sp12to4
    port map (
            O => \N__5861\,
            I => \N__5857\
        );

    \I__912\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5854\
        );

    \I__911\ : Span12Mux_h
    port map (
            O => \N__5857\,
            I => \N__5849\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5854\,
            I => \N__5849\
        );

    \I__909\ : Span12Mux_v
    port map (
            O => \N__5849\,
            I => \N__5846\
        );

    \I__908\ : Odrv12
    port map (
            O => \N__5846\,
            I => \D_in_5\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__5843\,
            I => \U409_AUTOCONFIG.N_49_cascade_\
        );

    \I__906\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5837\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5837\,
            I => \U409_AUTOCONFIG.N_107\
        );

    \I__904\ : InMux
    port map (
            O => \N__5834\,
            I => \N__5831\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5831\,
            I => \U409_AUTOCONFIG.N_95\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__5828\,
            I => \U409_AUTOCONFIG.N_48_cascade_\
        );

    \I__901\ : InMux
    port map (
            O => \N__5825\,
            I => \N__5822\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__5822\,
            I => \N__5818\
        );

    \I__899\ : InMux
    port map (
            O => \N__5821\,
            I => \N__5815\
        );

    \I__898\ : Span4Mux_h
    port map (
            O => \N__5818\,
            I => \N__5810\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5815\,
            I => \N__5810\
        );

    \I__896\ : Span4Mux_v
    port map (
            O => \N__5810\,
            I => \N__5807\
        );

    \I__895\ : Odrv4
    port map (
            O => \N__5807\,
            I => \U409_AUTOCONFIG.un1_A_13\
        );

    \I__894\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5801\,
            I => \U409_AUTOCONFIG.STATE_d_2\
        );

    \I__892\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5792\
        );

    \I__891\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5792\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5792\,
            I => \LIDE_BASE_7\
        );

    \I__889\ : InMux
    port map (
            O => \N__5789\,
            I => \N__5786\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5786\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__5783\,
            I => \N__5776\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__5782\,
            I => \N__5773\
        );

    \I__885\ : CascadeMux
    port map (
            O => \N__5781\,
            I => \N__5770\
        );

    \I__884\ : CascadeMux
    port map (
            O => \N__5780\,
            I => \N__5766\
        );

    \I__883\ : InMux
    port map (
            O => \N__5779\,
            I => \N__5763\
        );

    \I__882\ : InMux
    port map (
            O => \N__5776\,
            I => \N__5757\
        );

    \I__881\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5757\
        );

    \I__880\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5750\
        );

    \I__879\ : InMux
    port map (
            O => \N__5769\,
            I => \N__5750\
        );

    \I__878\ : InMux
    port map (
            O => \N__5766\,
            I => \N__5750\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5763\,
            I => \N__5746\
        );

    \I__876\ : InMux
    port map (
            O => \N__5762\,
            I => \N__5743\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5757\,
            I => \N__5740\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5750\,
            I => \N__5737\
        );

    \I__873\ : InMux
    port map (
            O => \N__5749\,
            I => \N__5734\
        );

    \I__872\ : Span4Mux_v
    port map (
            O => \N__5746\,
            I => \N__5729\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5743\,
            I => \N__5729\
        );

    \I__870\ : Odrv4
    port map (
            O => \N__5740\,
            I => \U409_AUTOCONFIG.un1_STATE_6_0\
        );

    \I__869\ : Odrv4
    port map (
            O => \N__5737\,
            I => \U409_AUTOCONFIG.un1_STATE_6_0\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__5734\,
            I => \U409_AUTOCONFIG.un1_STATE_6_0\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__5729\,
            I => \U409_AUTOCONFIG.un1_STATE_6_0\
        );

    \I__866\ : InMux
    port map (
            O => \N__5720\,
            I => \N__5713\
        );

    \I__865\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5713\
        );

    \I__864\ : InMux
    port map (
            O => \N__5718\,
            I => \N__5706\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5713\,
            I => \N__5703\
        );

    \I__862\ : InMux
    port map (
            O => \N__5712\,
            I => \N__5698\
        );

    \I__861\ : InMux
    port map (
            O => \N__5711\,
            I => \N__5698\
        );

    \I__860\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5694\
        );

    \I__859\ : InMux
    port map (
            O => \N__5709\,
            I => \N__5691\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5706\,
            I => \N__5684\
        );

    \I__857\ : Span4Mux_v
    port map (
            O => \N__5703\,
            I => \N__5684\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__5698\,
            I => \N__5684\
        );

    \I__855\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5681\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5694\,
            I => \U409_AUTOCONFIG.N_48\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5691\,
            I => \U409_AUTOCONFIG.N_48\
        );

    \I__852\ : Odrv4
    port map (
            O => \N__5684\,
            I => \U409_AUTOCONFIG.N_48\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5681\,
            I => \U409_AUTOCONFIG.N_48\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__5672\,
            I => \N__5669\
        );

    \I__849\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5658\
        );

    \I__848\ : InMux
    port map (
            O => \N__5668\,
            I => \N__5658\
        );

    \I__847\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5658\
        );

    \I__846\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5655\
        );

    \I__845\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5652\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5658\,
            I => \N__5649\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__5655\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5652\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__841\ : Odrv4
    port map (
            O => \N__5649\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__840\ : InMux
    port map (
            O => \N__5642\,
            I => \N__5639\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__5639\,
            I => \N__5636\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__5636\,
            I => \U409_ADDRESS_DECODE.LOWROMZ0Z_3\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__5633\,
            I => \N__5628\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__5632\,
            I => \N__5625\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__5631\,
            I => \N__5620\
        );

    \I__834\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5614\
        );

    \I__833\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5609\
        );

    \I__832\ : InMux
    port map (
            O => \N__5624\,
            I => \N__5609\
        );

    \I__831\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5604\
        );

    \I__830\ : InMux
    port map (
            O => \N__5620\,
            I => \N__5604\
        );

    \I__829\ : InMux
    port map (
            O => \N__5619\,
            I => \N__5600\
        );

    \I__828\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5597\
        );

    \I__827\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5594\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5614\,
            I => \N__5587\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5609\,
            I => \N__5587\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5604\,
            I => \N__5587\
        );

    \I__823\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5584\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5600\,
            I => \N__5576\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5597\,
            I => \N__5576\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5594\,
            I => \N__5576\
        );

    \I__819\ : Span4Mux_v
    port map (
            O => \N__5587\,
            I => \N__5571\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5584\,
            I => \N__5571\
        );

    \I__817\ : InMux
    port map (
            O => \N__5583\,
            I => \N__5568\
        );

    \I__816\ : Span4Mux_v
    port map (
            O => \N__5576\,
            I => \N__5565\
        );

    \I__815\ : Span4Mux_h
    port map (
            O => \N__5571\,
            I => \N__5560\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__5568\,
            I => \N__5560\
        );

    \I__813\ : Span4Mux_v
    port map (
            O => \N__5565\,
            I => \N__5557\
        );

    \I__812\ : Span4Mux_v
    port map (
            O => \N__5560\,
            I => \N__5554\
        );

    \I__811\ : Sp12to4
    port map (
            O => \N__5557\,
            I => \N__5549\
        );

    \I__810\ : Sp12to4
    port map (
            O => \N__5554\,
            I => \N__5549\
        );

    \I__809\ : Odrv12
    port map (
            O => \N__5549\,
            I => \A_c_21\
        );

    \I__808\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5542\
        );

    \I__807\ : InMux
    port map (
            O => \N__5545\,
            I => \N__5537\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5542\,
            I => \N__5533\
        );

    \I__805\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5530\
        );

    \I__804\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5527\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5537\,
            I => \N__5524\
        );

    \I__802\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5521\
        );

    \I__801\ : Span4Mux_v
    port map (
            O => \N__5533\,
            I => \N__5512\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__5530\,
            I => \N__5512\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5527\,
            I => \N__5512\
        );

    \I__798\ : Span4Mux_h
    port map (
            O => \N__5524\,
            I => \N__5507\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5521\,
            I => \N__5507\
        );

    \I__796\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5504\
        );

    \I__795\ : InMux
    port map (
            O => \N__5519\,
            I => \N__5501\
        );

    \I__794\ : Span4Mux_v
    port map (
            O => \N__5512\,
            I => \N__5498\
        );

    \I__793\ : Span4Mux_v
    port map (
            O => \N__5507\,
            I => \N__5495\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5504\,
            I => \N__5492\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__5501\,
            I => \N__5489\
        );

    \I__790\ : Sp12to4
    port map (
            O => \N__5498\,
            I => \N__5482\
        );

    \I__789\ : Sp12to4
    port map (
            O => \N__5495\,
            I => \N__5482\
        );

    \I__788\ : Span12Mux_v
    port map (
            O => \N__5492\,
            I => \N__5482\
        );

    \I__787\ : Span12Mux_h
    port map (
            O => \N__5489\,
            I => \N__5479\
        );

    \I__786\ : Odrv12
    port map (
            O => \N__5482\,
            I => \A_c_20\
        );

    \I__785\ : Odrv12
    port map (
            O => \N__5479\,
            I => \A_c_20\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__783\ : InMux
    port map (
            O => \N__5471\,
            I => \N__5468\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__781\ : Odrv4
    port map (
            O => \N__5465\,
            I => \U409_AUTOCONFIG.PR_OUTZ0Z_2\
        );

    \I__780\ : IoInMux
    port map (
            O => \N__5462\,
            I => \N__5459\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5459\,
            I => \N__5456\
        );

    \I__778\ : Span12Mux_s6_v
    port map (
            O => \N__5456\,
            I => \N__5453\
        );

    \I__777\ : Odrv12
    port map (
            O => \N__5453\,
            I => \D_OUT_2\
        );

    \I__776\ : InMux
    port map (
            O => \N__5450\,
            I => \N__5447\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5447\,
            I => \N__5444\
        );

    \I__774\ : Span4Mux_h
    port map (
            O => \N__5444\,
            I => \N__5441\
        );

    \I__773\ : Odrv4
    port map (
            O => \N__5441\,
            I => \U409_AUTOCONFIG.N_97\
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__5438\,
            I => \U409_AUTOCONFIG.STATE_d_2_cascade_\
        );

    \I__771\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5429\
        );

    \I__770\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5429\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5429\,
            I => \N__5426\
        );

    \I__768\ : Span12Mux_v
    port map (
            O => \N__5426\,
            I => \N__5423\
        );

    \I__767\ : Odrv12
    port map (
            O => \N__5423\,
            I => \D_in_6\
        );

    \I__766\ : InMux
    port map (
            O => \N__5420\,
            I => \N__5417\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__5417\,
            I => \U409_AUTOCONFIG.N_105\
        );

    \I__764\ : InMux
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5411\,
            I => \N__5404\
        );

    \I__762\ : InMux
    port map (
            O => \N__5410\,
            I => \N__5399\
        );

    \I__761\ : InMux
    port map (
            O => \N__5409\,
            I => \N__5399\
        );

    \I__760\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5396\
        );

    \I__759\ : InMux
    port map (
            O => \N__5407\,
            I => \N__5393\
        );

    \I__758\ : Odrv12
    port map (
            O => \N__5404\,
            I => \U409_AUTOCONFIG.N_49\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__5399\,
            I => \U409_AUTOCONFIG.N_49\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5396\,
            I => \U409_AUTOCONFIG.N_49\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__5393\,
            I => \U409_AUTOCONFIG.N_49\
        );

    \I__754\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5381\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5381\,
            I => \U409_AUTOCONFIG.PR_OUT_cnst_i_i_0_0_2\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__5378\,
            I => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1_cascade_\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__750\ : InMux
    port map (
            O => \N__5372\,
            I => \N__5365\
        );

    \I__749\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5360\
        );

    \I__748\ : InMux
    port map (
            O => \N__5370\,
            I => \N__5360\
        );

    \I__747\ : InMux
    port map (
            O => \N__5369\,
            I => \N__5356\
        );

    \I__746\ : InMux
    port map (
            O => \N__5368\,
            I => \N__5353\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__5365\,
            I => \N__5348\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5360\,
            I => \N__5348\
        );

    \I__743\ : CascadeMux
    port map (
            O => \N__5359\,
            I => \N__5345\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__5356\,
            I => \N__5340\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__5353\,
            I => \N__5340\
        );

    \I__740\ : Span4Mux_v
    port map (
            O => \N__5348\,
            I => \N__5337\
        );

    \I__739\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5334\
        );

    \I__738\ : Span4Mux_v
    port map (
            O => \N__5340\,
            I => \N__5331\
        );

    \I__737\ : Sp12to4
    port map (
            O => \N__5337\,
            I => \N__5324\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__5334\,
            I => \N__5324\
        );

    \I__735\ : Sp12to4
    port map (
            O => \N__5331\,
            I => \N__5324\
        );

    \I__734\ : Span12Mux_h
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__733\ : Span12Mux_v
    port map (
            O => \N__5321\,
            I => \N__5318\
        );

    \I__732\ : Odrv12
    port map (
            O => \N__5318\,
            I => \A_c_19\
        );

    \I__731\ : InMux
    port map (
            O => \N__5315\,
            I => \N__5309\
        );

    \I__730\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5309\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__5309\,
            I => \U409_AUTOCONFIG.N_84\
        );

    \I__728\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5303\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__5303\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\
        );

    \I__726\ : InMux
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5297\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\
        );

    \I__724\ : InMux
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__5291\,
            I => \N__5287\
        );

    \I__722\ : InMux
    port map (
            O => \N__5290\,
            I => \N__5284\
        );

    \I__721\ : Span4Mux_v
    port map (
            O => \N__5287\,
            I => \N__5281\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5284\,
            I => \N__5278\
        );

    \I__719\ : Span4Mux_h
    port map (
            O => \N__5281\,
            I => \N__5273\
        );

    \I__718\ : Span4Mux_h
    port map (
            O => \N__5278\,
            I => \N__5273\
        );

    \I__717\ : Span4Mux_v
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__716\ : Span4Mux_v
    port map (
            O => \N__5270\,
            I => \N__5267\
        );

    \I__715\ : Odrv4
    port map (
            O => \N__5267\,
            I => \D_in_7\
        );

    \I__714\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5261\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__5261\,
            I => \U409_ADDRESS_DECODE.PORTSIZEZ0Z_1\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__5258\,
            I => \U409_ADDRESS_DECODE.PORTSIZEZ0Z_0_cascade_\
        );

    \I__711\ : IoInMux
    port map (
            O => \N__5255\,
            I => \N__5252\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__709\ : IoSpan4Mux
    port map (
            O => \N__5249\,
            I => \N__5246\
        );

    \I__708\ : Span4Mux_s2_v
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__707\ : Sp12to4
    port map (
            O => \N__5243\,
            I => \N__5240\
        );

    \I__706\ : Span12Mux_s8_v
    port map (
            O => \N__5240\,
            I => \N__5237\
        );

    \I__705\ : Odrv12
    port map (
            O => \N__5237\,
            I => \PORTSIZE_0_i\
        );

    \I__704\ : IoInMux
    port map (
            O => \N__5234\,
            I => \N__5231\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5231\,
            I => \N__5228\
        );

    \I__702\ : Span4Mux_s3_v
    port map (
            O => \N__5228\,
            I => \N__5225\
        );

    \I__701\ : Span4Mux_v
    port map (
            O => \N__5225\,
            I => \N__5222\
        );

    \I__700\ : Sp12to4
    port map (
            O => \N__5222\,
            I => \N__5219\
        );

    \I__699\ : Span12Mux_h
    port map (
            O => \N__5219\,
            I => \N__5216\
        );

    \I__698\ : Odrv12
    port map (
            O => \N__5216\,
            I => \BUFENn_c\
        );

    \I__697\ : IoInMux
    port map (
            O => \N__5213\,
            I => \N__5210\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5210\,
            I => \N__5207\
        );

    \I__695\ : IoSpan4Mux
    port map (
            O => \N__5207\,
            I => \N__5204\
        );

    \I__694\ : Span4Mux_s2_h
    port map (
            O => \N__5204\,
            I => \N__5201\
        );

    \I__693\ : Sp12to4
    port map (
            O => \N__5201\,
            I => \N__5198\
        );

    \I__692\ : Span12Mux_s9_h
    port map (
            O => \N__5198\,
            I => \N__5195\
        );

    \I__691\ : Odrv12
    port map (
            O => \N__5195\,
            I => \U409_ADDRESS_DECODE_un1_ATA_ENn_i\
        );

    \I__690\ : CascadeMux
    port map (
            O => \N__5192\,
            I => \N__5188\
        );

    \I__689\ : InMux
    port map (
            O => \N__5191\,
            I => \N__5183\
        );

    \I__688\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5180\
        );

    \I__687\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5177\
        );

    \I__686\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5174\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__5183\,
            I => \N__5169\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__5180\,
            I => \N__5169\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__5177\,
            I => \N__5164\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5174\,
            I => \N__5164\
        );

    \I__681\ : Span4Mux_h
    port map (
            O => \N__5169\,
            I => \N__5161\
        );

    \I__680\ : Span12Mux_h
    port map (
            O => \N__5164\,
            I => \N__5156\
        );

    \I__679\ : Sp12to4
    port map (
            O => \N__5161\,
            I => \N__5156\
        );

    \I__678\ : Span12Mux_v
    port map (
            O => \N__5156\,
            I => \N__5153\
        );

    \I__677\ : Odrv12
    port map (
            O => \N__5153\,
            I => \A_c_18\
        );

    \I__676\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5146\
        );

    \I__675\ : InMux
    port map (
            O => \N__5149\,
            I => \N__5143\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__5146\,
            I => \LIDE_BASE_2\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__5143\,
            I => \LIDE_BASE_2\
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__5138\,
            I => \N__5134\
        );

    \I__671\ : CascadeMux
    port map (
            O => \N__5137\,
            I => \N__5131\
        );

    \I__670\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5128\
        );

    \I__669\ : InMux
    port map (
            O => \N__5131\,
            I => \N__5122\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5128\,
            I => \N__5119\
        );

    \I__667\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5116\
        );

    \I__666\ : InMux
    port map (
            O => \N__5126\,
            I => \N__5113\
        );

    \I__665\ : InMux
    port map (
            O => \N__5125\,
            I => \N__5110\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5122\,
            I => \N__5107\
        );

    \I__663\ : Span4Mux_h
    port map (
            O => \N__5119\,
            I => \N__5100\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__5116\,
            I => \N__5100\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5113\,
            I => \N__5100\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__5110\,
            I => \N__5093\
        );

    \I__659\ : Sp12to4
    port map (
            O => \N__5107\,
            I => \N__5093\
        );

    \I__658\ : Sp12to4
    port map (
            O => \N__5100\,
            I => \N__5093\
        );

    \I__657\ : Span12Mux_v
    port map (
            O => \N__5093\,
            I => \N__5090\
        );

    \I__656\ : Odrv12
    port map (
            O => \N__5090\,
            I => \A_c_17\
        );

    \I__655\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5083\
        );

    \I__654\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5080\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__5083\,
            I => \LIDE_BASE_1\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__5080\,
            I => \LIDE_BASE_1\
        );

    \I__651\ : InMux
    port map (
            O => \N__5075\,
            I => \N__5072\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__5072\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\
        );

    \I__649\ : CascadeMux
    port map (
            O => \N__5069\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_\
        );

    \I__648\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5063\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__5063\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2\
        );

    \I__646\ : InMux
    port map (
            O => \N__5060\,
            I => \N__5051\
        );

    \I__645\ : InMux
    port map (
            O => \N__5059\,
            I => \N__5051\
        );

    \I__644\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5051\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__5051\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__5048\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_\
        );

    \I__641\ : InMux
    port map (
            O => \N__5045\,
            I => \N__5036\
        );

    \I__640\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5036\
        );

    \I__639\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5036\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__5036\,
            I => \U409_ADDRESS_DECODE.ATA_ENZ0\
        );

    \I__637\ : CascadeMux
    port map (
            O => \N__5033\,
            I => \U409_AUTOCONFIG.N_121_cascade_\
        );

    \I__636\ : InMux
    port map (
            O => \N__5030\,
            I => \N__5025\
        );

    \I__635\ : InMux
    port map (
            O => \N__5029\,
            I => \N__5021\
        );

    \I__634\ : InMux
    port map (
            O => \N__5028\,
            I => \N__5018\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5025\,
            I => \N__5015\
        );

    \I__632\ : CascadeMux
    port map (
            O => \N__5024\,
            I => \N__5012\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__5021\,
            I => \N__5007\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__5018\,
            I => \N__5007\
        );

    \I__629\ : Span4Mux_v
    port map (
            O => \N__5015\,
            I => \N__5004\
        );

    \I__628\ : InMux
    port map (
            O => \N__5012\,
            I => \N__5001\
        );

    \I__627\ : Span12Mux_v
    port map (
            O => \N__5007\,
            I => \N__4994\
        );

    \I__626\ : Sp12to4
    port map (
            O => \N__5004\,
            I => \N__4994\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__5001\,
            I => \N__4994\
        );

    \I__624\ : Odrv12
    port map (
            O => \N__4994\,
            I => \A_c_7\
        );

    \I__623\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4987\
        );

    \I__622\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4984\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__4987\,
            I => \N__4981\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__4984\,
            I => \N__4978\
        );

    \I__619\ : Span4Mux_v
    port map (
            O => \N__4981\,
            I => \N__4968\
        );

    \I__618\ : Span4Mux_v
    port map (
            O => \N__4978\,
            I => \N__4968\
        );

    \I__617\ : InMux
    port map (
            O => \N__4977\,
            I => \N__4961\
        );

    \I__616\ : InMux
    port map (
            O => \N__4976\,
            I => \N__4961\
        );

    \I__615\ : InMux
    port map (
            O => \N__4975\,
            I => \N__4961\
        );

    \I__614\ : InMux
    port map (
            O => \N__4974\,
            I => \N__4956\
        );

    \I__613\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4956\
        );

    \I__612\ : Sp12to4
    port map (
            O => \N__4968\,
            I => \N__4949\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__4961\,
            I => \N__4949\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4956\,
            I => \N__4949\
        );

    \I__609\ : Odrv12
    port map (
            O => \N__4949\,
            I => \A_c_6\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__4946\,
            I => \N__4942\
        );

    \I__607\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4939\
        );

    \I__606\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4935\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4939\,
            I => \N__4932\
        );

    \I__604\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4929\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4935\,
            I => \N__4925\
        );

    \I__602\ : Span4Mux_v
    port map (
            O => \N__4932\,
            I => \N__4922\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__4929\,
            I => \N__4919\
        );

    \I__600\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4916\
        );

    \I__599\ : Span12Mux_v
    port map (
            O => \N__4925\,
            I => \N__4907\
        );

    \I__598\ : Sp12to4
    port map (
            O => \N__4922\,
            I => \N__4907\
        );

    \I__597\ : Sp12to4
    port map (
            O => \N__4919\,
            I => \N__4907\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__4916\,
            I => \N__4907\
        );

    \I__595\ : Odrv12
    port map (
            O => \N__4907\,
            I => \A_c_5\
        );

    \I__594\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4894\
        );

    \I__593\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4894\
        );

    \I__592\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4889\
        );

    \I__591\ : InMux
    port map (
            O => \N__4901\,
            I => \N__4889\
        );

    \I__590\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4884\
        );

    \I__589\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4884\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4894\,
            I => \N__4879\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4889\,
            I => \N__4879\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4884\,
            I => \N__4876\
        );

    \I__585\ : Sp12to4
    port map (
            O => \N__4879\,
            I => \N__4873\
        );

    \I__584\ : Span12Mux_h
    port map (
            O => \N__4876\,
            I => \N__4870\
        );

    \I__583\ : Span12Mux_v
    port map (
            O => \N__4873\,
            I => \N__4867\
        );

    \I__582\ : Span12Mux_v
    port map (
            O => \N__4870\,
            I => \N__4864\
        );

    \I__581\ : Odrv12
    port map (
            O => \N__4867\,
            I => \A_c_3\
        );

    \I__580\ : Odrv12
    port map (
            O => \N__4864\,
            I => \A_c_3\
        );

    \I__579\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4854\
        );

    \I__578\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4849\
        );

    \I__577\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4849\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__4854\,
            I => \U409_AUTOCONFIG.N_121\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__4849\,
            I => \U409_AUTOCONFIG.N_121\
        );

    \I__574\ : CascadeMux
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__573\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4838\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__571\ : Odrv12
    port map (
            O => \N__4835\,
            I => \U409_AUTOCONFIG.N_123\
        );

    \I__570\ : CascadeMux
    port map (
            O => \N__4832\,
            I => \N__4828\
        );

    \I__569\ : InMux
    port map (
            O => \N__4831\,
            I => \N__4825\
        );

    \I__568\ : InMux
    port map (
            O => \N__4828\,
            I => \N__4822\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4825\,
            I => \N__4819\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4822\,
            I => \N__4816\
        );

    \I__565\ : Span4Mux_v
    port map (
            O => \N__4819\,
            I => \N__4811\
        );

    \I__564\ : Span4Mux_v
    port map (
            O => \N__4816\,
            I => \N__4808\
        );

    \I__563\ : InMux
    port map (
            O => \N__4815\,
            I => \N__4805\
        );

    \I__562\ : InMux
    port map (
            O => \N__4814\,
            I => \N__4802\
        );

    \I__561\ : Span4Mux_v
    port map (
            O => \N__4811\,
            I => \N__4799\
        );

    \I__560\ : Span4Mux_v
    port map (
            O => \N__4808\,
            I => \N__4792\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4805\,
            I => \N__4792\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__4802\,
            I => \N__4792\
        );

    \I__557\ : Span4Mux_v
    port map (
            O => \N__4799\,
            I => \N__4789\
        );

    \I__556\ : Span4Mux_v
    port map (
            O => \N__4792\,
            I => \N__4786\
        );

    \I__555\ : Sp12to4
    port map (
            O => \N__4789\,
            I => \N__4781\
        );

    \I__554\ : Sp12to4
    port map (
            O => \N__4786\,
            I => \N__4781\
        );

    \I__553\ : Odrv12
    port map (
            O => \N__4781\,
            I => \A_c_16\
        );

    \I__552\ : InMux
    port map (
            O => \N__4778\,
            I => \N__4774\
        );

    \I__551\ : InMux
    port map (
            O => \N__4777\,
            I => \N__4771\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__4774\,
            I => \N__4766\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4771\,
            I => \N__4766\
        );

    \I__548\ : Span4Mux_v
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__547\ : Sp12to4
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__546\ : Odrv12
    port map (
            O => \N__4760\,
            I => \A_c_15\
        );

    \I__545\ : IoInMux
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4754\,
            I => \N__4749\
        );

    \I__543\ : IoInMux
    port map (
            O => \N__4753\,
            I => \N__4746\
        );

    \I__542\ : IoInMux
    port map (
            O => \N__4752\,
            I => \N__4743\
        );

    \I__541\ : IoSpan4Mux
    port map (
            O => \N__4749\,
            I => \N__4739\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4746\,
            I => \N__4734\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4743\,
            I => \N__4734\
        );

    \I__538\ : IoInMux
    port map (
            O => \N__4742\,
            I => \N__4731\
        );

    \I__537\ : Span4Mux_s3_v
    port map (
            O => \N__4739\,
            I => \N__4728\
        );

    \I__536\ : Span4Mux_s3_v
    port map (
            O => \N__4734\,
            I => \N__4725\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4731\,
            I => \N__4722\
        );

    \I__534\ : Span4Mux_v
    port map (
            O => \N__4728\,
            I => \N__4717\
        );

    \I__533\ : Span4Mux_v
    port map (
            O => \N__4725\,
            I => \N__4717\
        );

    \I__532\ : Span12Mux_s8_v
    port map (
            O => \N__4722\,
            I => \N__4714\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__4717\,
            I => \D_1_i\
        );

    \I__530\ : Odrv12
    port map (
            O => \N__4714\,
            I => \D_1_i\
        );

    \I__529\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4706\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__4706\,
            I => \N__4703\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__4703\,
            I => \U409_AUTOCONFIG.N_103\
        );

    \I__526\ : CascadeMux
    port map (
            O => \N__4700\,
            I => \N__4697\
        );

    \I__525\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4694\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4694\,
            I => \N__4690\
        );

    \I__523\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4687\
        );

    \I__522\ : Odrv4
    port map (
            O => \N__4690\,
            I => \LIDE_BASE_4\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4687\,
            I => \LIDE_BASE_4\
        );

    \I__520\ : InMux
    port map (
            O => \N__4682\,
            I => \N__4678\
        );

    \I__519\ : InMux
    port map (
            O => \N__4681\,
            I => \N__4675\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4678\,
            I => \LIDE_BASE_3\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4675\,
            I => \LIDE_BASE_3\
        );

    \I__516\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4667\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4667\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_5\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__4664\,
            I => \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0Z0Z_3_cascade_\
        );

    \I__513\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4658\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__4658\,
            I => \U409_ADDRESS_DECODE.HIROMZ0Z_0\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__4655\,
            I => \N__4652\
        );

    \I__510\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4649\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_0\
        );

    \I__508\ : CascadeMux
    port map (
            O => \N__4646\,
            I => \U409_AUTOCONFIG.N_99_cascade_\
        );

    \I__507\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4637\
        );

    \I__506\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4637\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4637\,
            I => \LIDE_BASE_5\
        );

    \I__504\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4631\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4631\,
            I => \N__4628\
        );

    \I__502\ : Sp12to4
    port map (
            O => \N__4628\,
            I => \N__4625\
        );

    \I__501\ : Span12Mux_v
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__500\ : Odrv12
    port map (
            O => \N__4622\,
            I => \D_in_4\
        );

    \I__499\ : InMux
    port map (
            O => \N__4619\,
            I => \N__4616\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4616\,
            I => \U409_AUTOCONFIG.N_101\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__4613\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2_cascade_\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__495\ : InMux
    port map (
            O => \N__4607\,
            I => \N__4604\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4604\,
            I => \N__4597\
        );

    \I__493\ : InMux
    port map (
            O => \N__4603\,
            I => \N__4594\
        );

    \I__492\ : InMux
    port map (
            O => \N__4602\,
            I => \N__4589\
        );

    \I__491\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4589\
        );

    \I__490\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4586\
        );

    \I__489\ : Odrv4
    port map (
            O => \N__4597\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4594\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4589\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__4586\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\
        );

    \I__485\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__4574\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2\
        );

    \I__483\ : IoInMux
    port map (
            O => \N__4571\,
            I => \N__4568\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4568\,
            I => \N__4565\
        );

    \I__481\ : Span4Mux_s3_v
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__480\ : Span4Mux_h
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__479\ : Sp12to4
    port map (
            O => \N__4559\,
            I => \N__4556\
        );

    \I__478\ : Span12Mux_v
    port map (
            O => \N__4556\,
            I => \N__4553\
        );

    \I__477\ : Span12Mux_h
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__476\ : Odrv12
    port map (
            O => \N__4550\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\
        );

    \I__475\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4544\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4544\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0Z0Z_0\
        );

    \I__473\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4538\,
            I => \N__4535\
        );

    \I__471\ : Span4Mux_h
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__470\ : Odrv4
    port map (
            O => \N__4532\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7\
        );

    \I__469\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4526\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4526\,
            I => \N__4523\
        );

    \I__467\ : Span4Mux_v
    port map (
            O => \N__4523\,
            I => \N__4520\
        );

    \I__466\ : IoSpan4Mux
    port map (
            O => \N__4520\,
            I => \N__4517\
        );

    \I__465\ : Odrv4
    port map (
            O => \N__4517\,
            I => \TT_c_1\
        );

    \I__464\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4511\,
            I => \N__4508\
        );

    \I__462\ : Span4Mux_h
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__461\ : Span4Mux_v
    port map (
            O => \N__4505\,
            I => \N__4502\
        );

    \I__460\ : Odrv4
    port map (
            O => \N__4502\,
            I => \TT_c_0\
        );

    \I__459\ : InMux
    port map (
            O => \N__4499\,
            I => \N__4495\
        );

    \I__458\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4492\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4495\,
            I => \LIDE_BASE_6\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4492\,
            I => \LIDE_BASE_6\
        );

    \I__455\ : CascadeMux
    port map (
            O => \N__4487\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_5_cascade_\
        );

    \I__454\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4480\
        );

    \I__453\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4477\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4480\,
            I => \N__4472\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__4477\,
            I => \N__4472\
        );

    \I__450\ : Span4Mux_v
    port map (
            O => \N__4472\,
            I => \N__4469\
        );

    \I__449\ : Span4Mux_h
    port map (
            O => \N__4469\,
            I => \N__4466\
        );

    \I__448\ : Odrv4
    port map (
            O => \N__4466\,
            I => \A_c_25\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__4463\,
            I => \N__4460\
        );

    \I__446\ : InMux
    port map (
            O => \N__4460\,
            I => \N__4457\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4457\,
            I => \N__4453\
        );

    \I__444\ : InMux
    port map (
            O => \N__4456\,
            I => \N__4450\
        );

    \I__443\ : Span4Mux_h
    port map (
            O => \N__4453\,
            I => \N__4445\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4450\,
            I => \N__4445\
        );

    \I__441\ : Span4Mux_v
    port map (
            O => \N__4445\,
            I => \N__4442\
        );

    \I__440\ : Span4Mux_h
    port map (
            O => \N__4442\,
            I => \N__4439\
        );

    \I__439\ : Odrv4
    port map (
            O => \N__4439\,
            I => \A_c_24\
        );

    \I__438\ : InMux
    port map (
            O => \N__4436\,
            I => \N__4433\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__4433\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4\
        );

    \I__436\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4424\
        );

    \I__435\ : InMux
    port map (
            O => \N__4429\,
            I => \N__4424\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__433\ : Span4Mux_v
    port map (
            O => \N__4421\,
            I => \N__4418\
        );

    \I__432\ : Span4Mux_h
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__431\ : Odrv4
    port map (
            O => \N__4415\,
            I => \A_c_29\
        );

    \I__430\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4406\
        );

    \I__429\ : InMux
    port map (
            O => \N__4411\,
            I => \N__4406\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__427\ : Span4Mux_v
    port map (
            O => \N__4403\,
            I => \N__4400\
        );

    \I__426\ : Span4Mux_h
    port map (
            O => \N__4400\,
            I => \N__4397\
        );

    \I__425\ : Odrv4
    port map (
            O => \N__4397\,
            I => \A_c_31\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__4394\,
            I => \N__4390\
        );

    \I__423\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4385\
        );

    \I__422\ : InMux
    port map (
            O => \N__4390\,
            I => \N__4385\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__4385\,
            I => \N__4382\
        );

    \I__420\ : Span4Mux_v
    port map (
            O => \N__4382\,
            I => \N__4379\
        );

    \I__419\ : Span4Mux_h
    port map (
            O => \N__4379\,
            I => \N__4376\
        );

    \I__418\ : Odrv4
    port map (
            O => \N__4376\,
            I => \A_c_30\
        );

    \I__417\ : InMux
    port map (
            O => \N__4373\,
            I => \N__4367\
        );

    \I__416\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4367\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__414\ : Span4Mux_v
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__413\ : Span4Mux_v
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__412\ : Sp12to4
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__411\ : Odrv12
    port map (
            O => \N__4355\,
            I => \A_c_28\
        );

    \I__410\ : IoInMux
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__408\ : IoSpan4Mux
    port map (
            O => \N__4346\,
            I => \N__4343\
        );

    \I__407\ : Span4Mux_s3_h
    port map (
            O => \N__4343\,
            I => \N__4340\
        );

    \I__406\ : Sp12to4
    port map (
            O => \N__4340\,
            I => \N__4337\
        );

    \I__405\ : Span12Mux_s11_h
    port map (
            O => \N__4337\,
            I => \N__4334\
        );

    \I__404\ : Span12Mux_h
    port map (
            O => \N__4334\,
            I => \N__4331\
        );

    \I__403\ : Odrv12
    port map (
            O => \N__4331\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn_i\
        );

    \I__402\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__4325\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0\
        );

    \I__400\ : CascadeMux
    port map (
            O => \N__4322\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_\
        );

    \I__399\ : CascadeMux
    port map (
            O => \N__4319\,
            I => \U409_ADDRESS_DECODE.HIROMZ0Z_0_cascade_\
        );

    \I__398\ : IoInMux
    port map (
            O => \N__4316\,
            I => \N__4313\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__396\ : Span12Mux_s2_h
    port map (
            O => \N__4310\,
            I => \N__4307\
        );

    \I__395\ : Span12Mux_v
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__394\ : Odrv12
    port map (
            O => \N__4304\,
            I => \SPIO_c\
        );

    \I__393\ : InMux
    port map (
            O => \N__4301\,
            I => \N__4298\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__4298\,
            I => \N__4294\
        );

    \I__391\ : InMux
    port map (
            O => \N__4297\,
            I => \N__4291\
        );

    \I__390\ : Span4Mux_v
    port map (
            O => \N__4294\,
            I => \N__4286\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__4291\,
            I => \N__4286\
        );

    \I__388\ : Span4Mux_h
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__387\ : Span4Mux_v
    port map (
            O => \N__4283\,
            I => \N__4280\
        );

    \I__386\ : Odrv4
    port map (
            O => \N__4280\,
            I => \A_c_26\
        );

    \I__385\ : CascadeMux
    port map (
            O => \N__4277\,
            I => \N__4274\
        );

    \I__384\ : InMux
    port map (
            O => \N__4274\,
            I => \N__4270\
        );

    \I__383\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4267\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__4270\,
            I => \N__4262\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__4267\,
            I => \N__4262\
        );

    \I__380\ : Span4Mux_v
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__379\ : Span4Mux_h
    port map (
            O => \N__4259\,
            I => \N__4256\
        );

    \I__378\ : Odrv4
    port map (
            O => \N__4256\,
            I => \A_c_27\
        );

    \I__377\ : IoInMux
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__4250\,
            I => \N__4247\
        );

    \I__375\ : IoSpan4Mux
    port map (
            O => \N__4247\,
            I => \N__4244\
        );

    \I__374\ : Sp12to4
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__373\ : Span12Mux_s1_h
    port map (
            O => \N__4241\,
            I => \N__4238\
        );

    \I__372\ : Span12Mux_v
    port map (
            O => \N__4238\,
            I => \N__4235\
        );

    \I__371\ : Odrv12
    port map (
            O => \N__4235\,
            I => \PPIO_c\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            I => \N__9161\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            I => \N__9160\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__9155\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            I => \N__9153\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            I => \N__9158\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            I => \N__9156\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            I => \N__9154\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            I => \N__9157\
        );

    \INVU409_AUTOCONFIG.AC_TACK_nesrC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.AC_TACK_nesrC_net\,
            I => \N__9821\
        );

    \INVU409_AUTOCONFIG.LIDE_OUT_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            I => \N__9820\
        );

    \INVU409_AUTOCONFIG.BRIDGE_OUT_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            I => \N__9824\
        );

    \INVU409_AUTOCONFIG.CONFIGUREDC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.CONFIGUREDC_net\,
            I => \N__9839\
        );

    \INVU409_AUTOCONFIG.LIDE_OUT_2C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_OUT_2C_net\,
            I => \N__9823\
        );

    \INVU409_AUTOCONFIG.STATE_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.STATE_0C_net\,
            I => \N__9833\
        );

    \INVU409_AUTOCONFIG.LIDE_BASE_7C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_BASE_7C_net\,
            I => \N__9838\
        );

    \INVU409_AUTOCONFIG.BRIDGE_OUT_3C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            I => \N__9830\
        );

    \INVU409_AUTOCONFIG.PR_OUT_2C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.PR_OUT_2C_net\,
            I => \N__9837\
        );

    \INVU409_AUTOCONFIG.LIDE_BASE_1C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            I => \N__9842\
        );

    \INVU409_AUTOCONFIG.LIDE_BASE_5C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_BASE_5C_net\,
            I => \N__9841\
        );

    \INVU409_AUTOCONFIG.LIDE_BASE_3C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_BASE_3C_net\,
            I => \N__9846\
        );

    \IN_MUX_bfv_17_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_5_0_\
        );

    \IN_MUX_bfv_17_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_17_6_0_\
        );

    \IN_MUX_bfv_15_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_6_0_\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_8_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8465\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_1_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4483\,
            in1 => \N__4273\,
            in2 => \N__4463\,
            in3 => \N__4301\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_5_LC_1_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4297\,
            in1 => \N__4412\,
            in2 => \N__4277\,
            in3 => \N__4373\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4436\,
            in1 => \N__4393\,
            in2 => \N__4487\,
            in3 => \N__4430\,
            lcout => \U409_ADDRESS_DECODE_Z2_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__4484\,
            in1 => \N__9062\,
            in2 => \_gnd_net_\,
            in3 => \N__4456\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4429\,
            in1 => \N__4411\,
            in2 => \N__4394\,
            in3 => \N__4372\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__5126\,
            in1 => \N__4328\,
            in2 => \N__4610\,
            in3 => \N__5619\,
            lcout => \U409_ADDRESS_DECODE_un1_RTC_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6267\,
            in1 => \N__5545\,
            in2 => \N__5192\,
            in3 => \N__5368\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0\,
            ltout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5127\,
            in1 => \N__4603\,
            in2 => \N__4322\,
            in3 => \N__5618\,
            lcout => \U409_ADDRESS_DECODE_un1_RTC_ENn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_0_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5536\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5617\,
            lcout => \U409_ADDRESS_DECODE.HIROMZ0Z_0\,
            ltout => \U409_ADDRESS_DECODE.HIROMZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6266\,
            in1 => \N__7946\,
            in2 => \N__4319\,
            in3 => \N__4600\,
            lcout => \CIA_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7710\,
            in2 => \_gnd_net_\,
            in3 => \N__6131\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6655\,
            in1 => \N__4547\,
            in2 => \N__5024\,
            in3 => \N__7314\,
            lcout => \U409_AUTOCONFIG.N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_5_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5186\,
            in1 => \N__5369\,
            in2 => \N__5137\,
            in3 => \N__4831\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_0_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4928\,
            in1 => \N__4973\,
            in2 => \N__6450\,
            in3 => \N__4901\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5030\,
            in1 => \N__4974\,
            in2 => \N__6451\,
            in3 => \N__4902\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_7_i_a3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100010"
        )
    port map (
            in0 => \N__7313\,
            in1 => \N__4945\,
            in2 => \_gnd_net_\,
            in3 => \N__6632\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_7_i_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4541\,
            in1 => \N__4529\,
            in2 => \_gnd_net_\,
            in3 => \N__4514\,
            lcout => \U409_ADDRESS_DECODE_AUTOVECTOR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_3_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111111000000"
        )
    port map (
            in0 => \N__5414\,
            in1 => \N__4709\,
            in2 => \N__5780\,
            in3 => \N__4682\,
            lcout => \LIDE_BASE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_3C_net\,
            ce => 'H',
            sr => \N__9751\
        );

    \U409_AUTOCONFIG.LIDE_BASE_6_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111111000000"
        )
    port map (
            in0 => \N__5719\,
            in1 => \N__5450\,
            in2 => \N__5781\,
            in3 => \N__4499\,
            lcout => \LIDE_BASE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_3C_net\,
            ce => 'H',
            sr => \N__9751\
        );

    \U409_AUTOCONFIG.LIDE_BASE_4_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011110000"
        )
    port map (
            in0 => \N__4619\,
            in1 => \N__5720\,
            in2 => \N__4700\,
            in3 => \N__5769\,
            lcout => \LIDE_BASE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_3C_net\,
            ce => 'H',
            sr => \N__9751\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__4498\,
            in1 => \N__6269\,
            in2 => \N__5633\,
            in3 => \N__4642\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_5_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5982\,
            in1 => \N__5718\,
            in2 => \N__5873\,
            in3 => \N__6902\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_5_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110110100000"
        )
    port map (
            in0 => \N__5749\,
            in1 => \N__5712\,
            in2 => \N__4646\,
            in3 => \N__4643\,
            lcout => \LIDE_BASE_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_5C_net\,
            ce => 'H',
            sr => \N__9749\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_4_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4634\,
            in1 => \N__5981\,
            in2 => \N__6924\,
            in3 => \N__5711\,
            lcout => \U409_AUTOCONFIG.N_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5541\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6268\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2\,
            ltout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7947\,
            in1 => \N__4601\,
            in2 => \N__4613\,
            in3 => \N__5624\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__4602\,
            in1 => \N__4577\,
            in2 => \N__5632\,
            in3 => \N__7948\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_1_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7876\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6879\,
            lcout => \U409_ADDRESS_DECODE.PORTSIZEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIU6QK1_1_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4991\,
            in1 => \N__6050\,
            in2 => \N__4844\,
            in3 => \N__7099\,
            lcout => \U409_AUTOCONFIG.un1_STATE_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5370\,
            in1 => \N__4670\,
            in2 => \N__4655\,
            in3 => \N__5603\,
            lcout => \AUTOCONFIG_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_5_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__7703\,
            in1 => \N__5187\,
            in2 => \N__4832\,
            in3 => \N__5125\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0_3_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__6513\,
            in1 => \N__6456\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0Z0Z_3\,
            ltout => \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110101"
        )
    port map (
            in0 => \N__9058\,
            in1 => \N__7320\,
            in2 => \N__4664\,
            in3 => \N__7477\,
            lcout => \U409_AUTOCONFIG.PR_OUT_cnst_i_i_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5371\,
            in1 => \N__4661\,
            in2 => \N__6135\,
            in3 => \N__6244\,
            lcout => \U409_ADDRESS_DECODE_HIROM\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_0_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5520\,
            in1 => \N__6238\,
            in2 => \_gnd_net_\,
            in3 => \N__6117\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_7_0_a3_3_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000001000"
        )
    port map (
            in0 => \N__7315\,
            in1 => \N__6495\,
            in2 => \N__6463\,
            in3 => \N__6656\,
            lcout => \U409_AUTOCONFIG.N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a3_2_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__4857\,
            in1 => \N__4976\,
            in2 => \_gnd_net_\,
            in3 => \N__7316\,
            lcout => \U409_AUTOCONFIG.N_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_13_0_a2_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4977\,
            in1 => \N__4858\,
            in2 => \N__7337\,
            in3 => \N__4904\,
            lcout => \U409_AUTOCONFIG.un1_A_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_2_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4938\,
            in1 => \N__5028\,
            in2 => \N__6673\,
            in3 => \N__6455\,
            lcout => \U409_AUTOCONFIG.N_121\,
            ltout => \U409_AUTOCONFIG.N_121_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__4975\,
            in1 => \_gnd_net_\,
            in2 => \N__5033\,
            in3 => \N__4903\,
            lcout => \U409_AUTOCONFIG.N_129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_3_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5029\,
            in1 => \N__4990\,
            in2 => \N__4946\,
            in3 => \N__4900\,
            lcout => \U409_AUTOCONFIG.N_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_0_3_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4899\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4859\,
            lcout => \U409_AUTOCONFIG.N_123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CS0_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__4814\,
            in1 => \N__4777\,
            in2 => \N__8383\,
            in3 => \N__8451\,
            lcout => \U409_ADDRESS_DECODE.CSZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CS1_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__4815\,
            in1 => \N__8379\,
            in2 => \N__8455\,
            in3 => \N__4778\,
            lcout => \U409_ADDRESS_DECODE.CSZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.D_1_i_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5985\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6936\,
            lcout => \D_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_3_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__6937\,
            in1 => \N__5290\,
            in2 => \N__5999\,
            in3 => \N__5408\,
            lcout => \U409_AUTOCONFIG.N_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__5546\,
            in1 => \N__4693\,
            in2 => \N__5359\,
            in3 => \N__4681\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_1_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111111000000"
        )
    port map (
            in0 => \N__5409\,
            in1 => \N__5840\,
            in2 => \N__5782\,
            in3 => \N__5087\,
            lcout => \LIDE_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            ce => 'H',
            sr => \N__9750\
        );

    \U409_AUTOCONFIG.LIDE_BASE_2_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111111000000"
        )
    port map (
            in0 => \N__5410\,
            in1 => \N__5420\,
            in2 => \N__5783\,
            in3 => \N__5150\,
            lcout => \LIDE_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            ce => 'H',
            sr => \N__9750\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_7_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5294\,
            in1 => \N__5984\,
            in2 => \N__6939\,
            in3 => \N__5709\,
            lcout => \U409_AUTOCONFIG.N_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8047\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7138\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.PORTSIZEZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNIOGLSO_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100111111"
        )
    port map (
            in0 => \N__5044\,
            in1 => \N__5264\,
            in2 => \N__5258\,
            in3 => \N__5058\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.LV_SPACE_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5060\,
            in1 => \N__7137\,
            in2 => \N__6935\,
            in3 => \N__7117\,
            lcout => \BUFENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5045\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5059\,
            lcout => \U409_ADDRESS_DECODE_un1_ATA_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__5191\,
            in1 => \N__5149\,
            in2 => \N__5138\,
            in3 => \N__5086\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5075\,
            in1 => \N__5789\,
            in2 => \N__5069\,
            in3 => \N__5066\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0\,
            ltout => \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010000"
        )
    port map (
            in0 => \N__5983\,
            in1 => \_gnd_net_\,
            in2 => \N__5048\,
            in3 => \N__5043\,
            lcout => \U409_ADDRESS_DECODE.ATA_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9840\,
            ce => 'H',
            sr => \N__9748\
        );

    \U409_AUTOCONFIG.PR_OUT_2_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__6712\,
            in1 => \N__6672\,
            in2 => \N__6464\,
            in3 => \N__5384\,
            lcout => \U409_AUTOCONFIG.PR_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.PR_OUT_2C_net\,
            ce => \N__7407\,
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_1_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5623\,
            in2 => \_gnd_net_\,
            in3 => \N__7704\,
            lcout => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1\,
            ltout => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6247\,
            in1 => \N__6184\,
            in2 => \N__5378\,
            in3 => \N__6138\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.LOWROM_3_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6137\,
            in1 => \N__6183\,
            in2 => \N__5375\,
            in3 => \N__6246\,
            lcout => \U409_ADDRESS_DECODE.LOWROMZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_4_0_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6245\,
            in1 => \N__6136\,
            in2 => \N__5631\,
            in3 => \N__5540\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTOR_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_1_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__6514\,
            in1 => \N__6457\,
            in2 => \_gnd_net_\,
            in3 => \N__6671\,
            lcout => \U409_AUTOCONFIG.N_131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__9045\,
            in1 => \N__7322\,
            in2 => \N__6553\,
            in3 => \N__5314\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            ce => \N__7412\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5315\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9046\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            ce => \N__7412\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5306\,
            in1 => \N__5300\,
            in2 => \_gnd_net_\,
            in3 => \N__6995\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_3_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6496\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7321\,
            lcout => \U409_AUTOCONFIG.N_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.LOWROM_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5642\,
            in1 => \N__5583\,
            in2 => \_gnd_net_\,
            in3 => \N__5519\,
            lcout => \U409_ADDRESS_DECODE_LOWROM\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__6566\,
            in1 => \N__7040\,
            in2 => \N__5474\,
            in3 => \N__6852\,
            lcout => \D_OUT_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_6_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5435\,
            in1 => \N__6011\,
            in2 => \N__6941\,
            in3 => \N__5697\,
            lcout => \U409_AUTOCONFIG.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIF4QU_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6049\,
            in2 => \_gnd_net_\,
            in3 => \N__7095\,
            lcout => \U409_AUTOCONFIG.STATE_d_2\,
            ltout => \U409_AUTOCONFIG.STATE_d_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5668\,
            in1 => \N__6984\,
            in2 => \N__5438\,
            in3 => \N__5825\,
            lcout => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_2_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5434\,
            in1 => \N__6010\,
            in2 => \N__6940\,
            in3 => \N__5407\,
            lcout => \U409_AUTOCONFIG.N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5672\,
            in3 => \N__6985\,
            lcout => \U409_AUTOCONFIG.N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__7339\,
            in1 => \N__5667\,
            in2 => \_gnd_net_\,
            in3 => \N__6983\,
            lcout => \U409_AUTOCONFIG.N_49\,
            ltout => \U409_AUTOCONFIG.N_49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_1_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6009\,
            in1 => \N__5860\,
            in2 => \N__5843\,
            in3 => \N__6928\,
            lcout => \U409_AUTOCONFIG.N_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__7338\,
            in1 => \N__5665\,
            in2 => \_gnd_net_\,
            in3 => \N__6981\,
            lcout => \U409_AUTOCONFIG.N_48\,
            ltout => \U409_AUTOCONFIG.N_48_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_7_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110110001000"
        )
    port map (
            in0 => \N__5779\,
            in1 => \N__5834\,
            in2 => \N__5828\,
            in3 => \N__5798\,
            lcout => \LIDE_BASE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_7C_net\,
            ce => 'H',
            sr => \N__9746\
        );

    \U409_AUTOCONFIG.BRIDGE_CONF_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__5821\,
            in1 => \N__5804\,
            in2 => \_gnd_net_\,
            in3 => \N__6982\,
            lcout => \U409_AUTOCONFIG.BRIDGE_CONFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_7C_net\,
            ce => 'H',
            sr => \N__9746\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000000000"
        )
    port map (
            in0 => \N__7690\,
            in1 => \N__5797\,
            in2 => \N__6143\,
            in3 => \N__6842\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100010"
        )
    port map (
            in0 => \N__6048\,
            in1 => \N__7094\,
            in2 => \N__5912\,
            in3 => \N__6809\,
            lcout => \U409_AUTOCONFIG.STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.STATE_0C_net\,
            ce => 'H',
            sr => \N__9743\
        );

    \U409_AUTOCONFIG.STATE_1_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111001100"
        )
    port map (
            in0 => \N__6001\,
            in1 => \N__6047\,
            in2 => \_gnd_net_\,
            in3 => \N__7093\,
            lcout => \U409_AUTOCONFIG.STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.STATE_0C_net\,
            ce => 'H',
            sr => \N__9743\
        );

    \U409_AUTOCONFIG.LIDE_CONF_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__5762\,
            in1 => \N__5666\,
            in2 => \_gnd_net_\,
            in3 => \N__5710\,
            lcout => \U409_AUTOCONFIG.LIDE_CONFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.STATE_0C_net\,
            ce => 'H',
            sr => \N__9743\
        );

    \U409_AUTOCONFIG.STATE_ns_1_0__m4_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100001010"
        )
    port map (
            in0 => \N__7088\,
            in1 => \_gnd_net_\,
            in2 => \N__6000\,
            in3 => \N__6042\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.STATE_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_TACK_nesr_RNO_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__9755\,
            in1 => \_gnd_net_\,
            in2 => \N__6272\,
            in3 => \_gnd_net_\,
            lcout => \U409_AUTOCONFIG.STATE_ns_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__6253\,
            in1 => \N__6194\,
            in2 => \N__6185\,
            in3 => \N__6139\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIBIND1_1_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6043\,
            in1 => \N__5989\,
            in2 => \_gnd_net_\,
            in3 => \N__7089\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_RNI10V92_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100110011"
        )
    port map (
            in0 => \N__5905\,
            in1 => \N__9035\,
            in2 => \N__5879\,
            in3 => \N__6808\,
            lcout => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNO_0_1_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6449\,
            in2 => \N__6524\,
            in3 => \N__7325\,
            lcout => \U409_AUTOCONFIG.N_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__6684\,
            in1 => \N__6520\,
            in2 => \N__6462\,
            in3 => \N__7324\,
            lcout => \U409_AUTOCONFIG.N_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6445\,
            in2 => \_gnd_net_\,
            in3 => \N__6670\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.N_227_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__6705\,
            in1 => \N__9041\,
            in2 => \N__5876\,
            in3 => \N__6533\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_2C_net\,
            ce => \N__7406\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000100"
        )
    port map (
            in0 => \N__6704\,
            in1 => \N__9040\,
            in2 => \N__6461\,
            in3 => \N__6532\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_2C_net\,
            ce => \N__7406\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6578\,
            in1 => \N__6994\,
            in2 => \_gnd_net_\,
            in3 => \N__6572\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6675\,
            in1 => \N__6512\,
            in2 => \_gnd_net_\,
            in3 => \N__6411\,
            lcout => \U409_AUTOCONFIG.N_133\,
            ltout => \U409_AUTOCONFIG.N_133_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_7_0_a2_2_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111010"
        )
    port map (
            in0 => \N__6557\,
            in1 => \_gnd_net_\,
            in2 => \N__6536\,
            in3 => \N__7323\,
            lcout => \U409_AUTOCONFIG.N_127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_1_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6674\,
            in1 => \N__6511\,
            in2 => \_gnd_net_\,
            in3 => \N__6410\,
            lcout => \U409_AUTOCONFIG.N_126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNISS912_1_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__7004\,
            in1 => \N__7044\,
            in2 => \N__6731\,
            in3 => \N__6848\,
            lcout => \D_OUT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001010"
        )
    port map (
            in0 => \N__6847\,
            in1 => \N__6341\,
            in2 => \N__7046\,
            in3 => \N__6761\,
            lcout => \D_OUT_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.CONFIGURED_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6308\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6846\,
            lcout => \CONFIGURED\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGUREDC_net\,
            ce => 'H',
            sr => \N__9747\
        );

    \U409_AUTOCONFIG.CONFIGENn_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6283\,
            in2 => \_gnd_net_\,
            in3 => \N__6307\,
            lcout => \CONFIGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGUREDC_net\,
            ce => 'H',
            sr => \N__9747\
        );

    \U409_AUTOCONFIG.PR_OUT_RNIPP912_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__6947\,
            in1 => \N__7045\,
            in2 => \N__6854\,
            in3 => \N__7454\,
            lcout => \D_OUT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNI7DMP_1_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6987\,
            in1 => \N__6782\,
            in2 => \_gnd_net_\,
            in3 => \N__6587\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_RNI7DMPZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNI5BMP_0_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7421\,
            in1 => \N__6797\,
            in2 => \_gnd_net_\,
            in3 => \N__6986\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_RNI5BMPZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__6938\,
            in1 => \N__7987\,
            in2 => \_gnd_net_\,
            in3 => \N__6853\,
            lcout => \U409_AUTOCONFIG.AC_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9831\,
            ce => 'H',
            sr => \N__9736\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000100"
        )
    port map (
            in0 => \N__7465\,
            in1 => \N__9025\,
            in2 => \N__6752\,
            in3 => \N__7333\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => \N__7390\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100010"
        )
    port map (
            in0 => \N__9027\,
            in1 => \N__7183\,
            in2 => \N__7340\,
            in3 => \N__6788\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => \N__7390\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_3_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__6719\,
            in1 => \N__9034\,
            in2 => \N__6773\,
            in3 => \N__6686\,
            lcout => \U409_AUTOCONFIG.PR_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => \N__7390\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7487\,
            in1 => \N__6751\,
            in2 => \N__9048\,
            in3 => \N__6737\,
            lcout => \U409_AUTOCONFIG.PR_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => \N__7390\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__6718\,
            in1 => \N__6685\,
            in2 => \N__7184\,
            in3 => \N__9026\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => \N__7390\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7486\,
            in1 => \N__7466\,
            in2 => \N__9047\,
            in3 => \N__7355\,
            lcout => \U409_AUTOCONFIG.PR_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => \N__7390\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__7445\,
            in1 => \N__7163\,
            in2 => \N__7436\,
            in3 => \N__9036\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            ce => \N__7411\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__7351\,
            in1 => \N__7332\,
            in2 => \N__7211\,
            in3 => \N__7174\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_7_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__7157\,
            in1 => \N__7142\,
            in2 => \N__7124\,
            in3 => \N__9007\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_TACK_nesr_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7100\,
            lcout => \AC_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.AC_TACK_nesrC_net\,
            ce => \N__7055\,
            sr => \N__9733\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8763\,
            in1 => \N__8832\,
            in2 => \N__8665\,
            in3 => \N__8734\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8802\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11149\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8602\,
            in1 => \N__8632\,
            in2 => \N__8701\,
            in3 => \N__8801\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_2_0\,
            ltout => \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__7786\,
            in1 => \N__8695\,
            in2 => \N__7508\,
            in3 => \N__7811\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11149\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__8314\,
            in1 => \N__7862\,
            in2 => \N__7850\,
            in3 => \N__8269\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__8086\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7860\,
            in1 => \N__8268\,
            in2 => \_gnd_net_\,
            in3 => \N__8313\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7843\,
            in2 => \N__7505\,
            in3 => \N__8230\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__8086\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__8229\,
            in1 => \N__8246\,
            in2 => \N__7502\,
            in3 => \N__7848\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__8086\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8124\,
            in1 => \N__8185\,
            in2 => \_gnd_net_\,
            in3 => \N__8207\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8291\,
            in2 => \N__7493\,
            in3 => \N__7847\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__8086\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_5_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__8008\,
            in1 => \N__9869\,
            in2 => \N__8156\,
            in3 => \N__8139\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__7861\,
            in1 => \_gnd_net_\,
            in2 => \N__7490\,
            in3 => \N__8315\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__8086\
        );

    \U409_TRANSFER_ACK.TACK_OUT_RNO_0_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10062\,
            in2 => \_gnd_net_\,
            in3 => \N__9185\,
            lcout => \U409_TRANSFER_ACK.TACK_EN8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_RNO_0_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111010"
        )
    port map (
            in0 => \N__10063\,
            in1 => \_gnd_net_\,
            in2 => \N__9193\,
            in3 => \N__7751\,
            lcout => \U409_TRANSFER_ACK.TACK_STATE_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUT_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110111001000"
        )
    port map (
            in0 => \N__7732\,
            in1 => \N__7586\,
            in2 => \N__7769\,
            in3 => \N__7752\,
            lcout => \TACK_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9818\,
            ce => 'H',
            sr => \N__9732\
        );

    \U409_TRANSFER_ACK.TACK_EN_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__9078\,
            in1 => \N__7731\,
            in2 => \_gnd_net_\,
            in3 => \N__7760\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9818\,
            ce => 'H',
            sr => \N__9732\
        );

    \U409_TRANSFER_ACK.TACK_STATE_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000100"
        )
    port map (
            in0 => \N__7754\,
            in1 => \N__10067\,
            in2 => \N__7733\,
            in3 => \N__9194\,
            lcout => \U409_TRANSFER_ACK.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9818\,
            ce => 'H',
            sr => \N__9732\
        );

    \U409_TRANSFER_ACK.TACK_STATE_1_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7753\,
            lcout => \U409_TRANSFER_ACK.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9818\,
            ce => 'H',
            sr => \N__9732\
        );

    \U409_TRANSFER_ACK.ROM_TACK_STATE5_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__7718\,
            in1 => \N__7565\,
            in2 => \N__7646\,
            in3 => \N__8007\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUT_RNIU3I06_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__7717\,
            in1 => \N__7645\,
            in2 => \N__7605\,
            in3 => \N__7561\,
            lcout => \U409_TRANSFER_ACK_un1_TACK_OUT_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9871\,
            lcout => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8730\,
            in2 => \N__8806\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8600\,
            in2 => \_gnd_net_\,
            in3 => \N__7820\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__11148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8629\,
            in2 => \_gnd_net_\,
            in3 => \N__7817\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8657\,
            in2 => \_gnd_net_\,
            in3 => \N__7814\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__11148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8696\,
            in2 => \_gnd_net_\,
            in3 => \N__7805\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_6_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8833\,
            in2 => \_gnd_net_\,
            in3 => \N__7802\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\,
            clk => \N__11148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_7_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8767\,
            in2 => \_gnd_net_\,
            in3 => \N__7799\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100101010"
        )
    port map (
            in0 => \N__8630\,
            in1 => \N__7796\,
            in2 => \N__7790\,
            in3 => \N__7775\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_1_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8762\,
            in2 => \_gnd_net_\,
            in3 => \N__8828\,
            lcout => \U409_CIA.CLK_CIA6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__8736\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8800\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_2_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8631\,
            in1 => \N__8601\,
            in2 => \N__8700\,
            in3 => \N__8799\,
            lcout => OPEN,
            ltout => \U409_CIA.un1_CIA_CLK_COUNT_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__8661\,
            in1 => \N__7895\,
            in2 => \N__7889\,
            in3 => \N__8735\,
            lcout => OPEN,
            ltout => \U409_CIA.VMA_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__8737\,
            in1 => \N__7886\,
            in2 => \N__7865\,
            in3 => \N__8544\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9311\,
            in2 => \_gnd_net_\,
            in3 => \N__9292\,
            lcout => \U409_TRANSFER_ACK.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8204\,
            in1 => \N__8118\,
            in2 => \N__8186\,
            in3 => \N__8290\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__8119\,
            in1 => \N__8184\,
            in2 => \_gnd_net_\,
            in3 => \N__8206\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__8090\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__8205\,
            in1 => \N__8120\,
            in2 => \_gnd_net_\,
            in3 => \N__7849\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__8090\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__8117\,
            in1 => \N__8289\,
            in2 => \N__8231\,
            in3 => \N__8244\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8312\,
            in1 => \N__8267\,
            in2 => \N__7823\,
            in3 => \N__8164\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8311\,
            in1 => \N__8288\,
            in2 => \N__8270\,
            in3 => \N__8245\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8126\,
            in1 => \N__8228\,
            in2 => \N__8210\,
            in3 => \N__8165\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8203\,
            in2 => \_gnd_net_\,
            in3 => \N__8180\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__8495\,
            in1 => \N__8140\,
            in2 => \_gnd_net_\,
            in3 => \N__8155\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            ce => 'H',
            sr => \N__8085\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000110011"
        )
    port map (
            in0 => \N__7997\,
            in1 => \N__8125\,
            in2 => \N__9872\,
            in3 => \N__8141\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            ce => 'H',
            sr => \N__8085\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_2_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__8054\,
            in1 => \N__7901\,
            in2 => \N__8033\,
            in3 => \N__8009\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_2\,
            ltout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERcZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__9864\,
            in1 => \_gnd_net_\,
            in2 => \N__7955\,
            in3 => \N__8476\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \N__9731\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_11_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7952\,
            in1 => \N__7928\,
            in2 => \N__9024\,
            in3 => \N__7919\,
            lcout => \U409_ADDRESS_DECODE_AUTOVECTOR_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8483\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8983\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__8477\,
            in1 => \N__9865\,
            in2 => \N__8468\,
            in3 => \N__9212\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \N__9731\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8969\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__8395\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8456\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNI692L_0_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8928\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8549\,
            lcout => \CIA_ENABLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8396\,
            in2 => \_gnd_net_\,
            in3 => \N__8384\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111101000101010"
        )
    port map (
            in0 => \N__9332\,
            in1 => \N__8321\,
            in2 => \N__8573\,
            in3 => \N__9338\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \N__9744\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__8568\,
            in1 => \N__9272\,
            in2 => \_gnd_net_\,
            in3 => \N__9344\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \N__9737\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111100001000"
        )
    port map (
            in0 => \N__9331\,
            in1 => \N__9353\,
            in2 => \N__8572\,
            in3 => \N__8507\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \N__9737\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8948\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8545\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \N__9737\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9293\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \N__9737\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9437\,
            in2 => \N__9958\,
            in3 => \N__9949\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_1_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9480\,
            in2 => \_gnd_net_\,
            in3 => \N__8528\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_0\,
            carryout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_2_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9244\,
            in2 => \_gnd_net_\,
            in3 => \N__8525\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_1\,
            carryout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_3_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9256\,
            in2 => \_gnd_net_\,
            in3 => \N__8522\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010001000"
        )
    port map (
            in0 => \N__8976\,
            in1 => \N__8519\,
            in2 => \N__9959\,
            in3 => \N__10036\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9825\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__10035\,
            in1 => \N__8513\,
            in2 => \N__9021\,
            in3 => \N__9957\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9825\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_START_RNO_1_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8506\,
            in2 => \_gnd_net_\,
            in3 => \N__8494\,
            lcout => \U409_TRANSFER_ACK.TACK_START_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__10037\,
            in1 => \N__9956\,
            in2 => \N__9022\,
            in3 => \N__9230\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9825\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_START_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__9224\,
            in1 => \N__9211\,
            in2 => \N__9192\,
            in3 => \N__9200\,
            lcout => \U409_TRANSFER_ACK.TACK_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9159\,
            ce => 'H',
            sr => \N__8849\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__10034\,
            in1 => \N__9131\,
            in2 => \N__9023\,
            in3 => \N__9936\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9819\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_START_RNO_0_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9096\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8984\,
            lcout => \U409_TRANSFER_ACK.TACK_RST_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_0_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8834\,
            in1 => \N__8807\,
            in2 => \N__8771\,
            in3 => \N__8741\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001101010"
        )
    port map (
            in0 => \N__9620\,
            in1 => \N__8579\,
            in2 => \N__8705\,
            in3 => \N__8702\,
            lcout => \CLK_CIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9583\,
            in1 => \N__9656\,
            in2 => \N__9527\,
            in3 => \N__9566\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_1_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011000"
        )
    port map (
            in0 => \N__8666\,
            in1 => \N__8636\,
            in2 => \N__9627\,
            in3 => \N__8606\,
            lcout => \U409_CIA.CLK_CIA_r_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9870\,
            in1 => \N__9597\,
            in2 => \_gnd_net_\,
            in3 => \N__9265\,
            lcout => \U409_TRANSFER_ACK.N_17_mux\,
            ltout => \U409_TRANSFER_ACK.N_17_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101011111"
        )
    port map (
            in0 => \N__9329\,
            in1 => \N__9309\,
            in2 => \N__9347\,
            in3 => \N__9290\,
            lcout => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9598\,
            in2 => \_gnd_net_\,
            in3 => \N__9266\,
            lcout => \U409_TRANSFER_ACK.N_3_0\,
            ltout => \U409_TRANSFER_ACK.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__9330\,
            in1 => \N__9310\,
            in2 => \N__9296\,
            in3 => \N__9291\,
            lcout => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10169\,
            in2 => \_gnd_net_\,
            in3 => \N__9584\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10869\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9599\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \N__9738\
        );

    \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m6_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100000000001"
        )
    port map (
            in0 => \N__9463\,
            in1 => \N__9481\,
            in2 => \N__9509\,
            in3 => \N__9435\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.N_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m10_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__9257\,
            in1 => \N__9245\,
            in2 => \N__9233\,
            in3 => \N__9419\,
            lcout => \U409_TRANSFER_ACK.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_STATE_ns_1_0__m8_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9508\,
            in1 => \N__9482\,
            in2 => \N__9467\,
            in3 => \N__9436\,
            lcout => \U409_TRANSFER_ACK.N_19_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_STATE_0_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111111010"
        )
    port map (
            in0 => \N__10015\,
            in1 => \N__10082\,
            in2 => \N__9982\,
            in3 => \N__9934\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9822\,
            ce => 'H',
            sr => \N__9734\
        );

    \U409_TICK.TICK60_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__10320\,
            in1 => \N__9397\,
            in2 => \N__10262\,
            in3 => \N__10284\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10619\,
            in1 => \N__10640\,
            in2 => \N__10685\,
            in3 => \N__11090\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10319\,
            in1 => \N__10283\,
            in2 => \N__9386\,
            in3 => \N__10667\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__10987\,
            in1 => \N__11032\,
            in2 => \N__10946\,
            in3 => \N__9370\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10340\,
            in1 => \N__10366\,
            in2 => \_gnd_net_\,
            in3 => \N__10424\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__9686\,
            in1 => \N__10580\,
            in2 => \N__9359\,
            in3 => \N__10388\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10318\,
            in1 => \N__10258\,
            in2 => \N__9356\,
            in3 => \N__10352\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__10945\,
            in1 => \N__11031\,
            in2 => \N__9542\,
            in3 => \N__10993\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10868\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9582\,
            in2 => \N__10164\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_6_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9565\,
            in2 => \_gnd_net_\,
            in3 => \N__9554\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__10870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10225\,
            in2 => \_gnd_net_\,
            in3 => \N__9551\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__10870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10492\,
            in2 => \_gnd_net_\,
            in3 => \N__9548\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__10870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10519\,
            in2 => \_gnd_net_\,
            in3 => \N__9545\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10102\,
            in2 => \_gnd_net_\,
            in3 => \N__9533\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10507\,
            in2 => \_gnd_net_\,
            in3 => \N__9530\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__10870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9523\,
            in2 => \_gnd_net_\,
            in3 => \N__9512\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__10870\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10117\,
            in2 => \_gnd_net_\,
            in3 => \N__9680\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10189\,
            in2 => \_gnd_net_\,
            in3 => \N__9677\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__10872\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10129\,
            in2 => \_gnd_net_\,
            in3 => \N__9674\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10204\,
            in2 => \_gnd_net_\,
            in3 => \N__9671\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__10872\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10892\,
            in2 => \_gnd_net_\,
            in3 => \N__9668\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10480\,
            in2 => \_gnd_net_\,
            in3 => \N__9665\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10459\,
            in2 => \_gnd_net_\,
            in3 => \N__9662\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9655\,
            in2 => \_gnd_net_\,
            in3 => \N__9659\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10872\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9628\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__9745\
        );

    \U409_TRANSFER_ACK.ROM_TACK_STATE_1_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__10011\,
            in1 => \N__10080\,
            in2 => \_gnd_net_\,
            in3 => \N__9932\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9832\,
            ce => 'H',
            sr => \N__9739\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000001010"
        )
    port map (
            in0 => \N__10058\,
            in1 => \N__10081\,
            in2 => \N__10023\,
            in3 => \N__9933\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9832\,
            ce => 'H',
            sr => \N__9739\
        );

    \U409_TRANSFER_ACK.ROMENn_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111010001100"
        )
    port map (
            in0 => \N__10016\,
            in1 => \N__9883\,
            in2 => \N__9986\,
            in3 => \N__9935\,
            lcout => \ROMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9826\,
            ce => 'H',
            sr => \N__9735\
        );

    \U409_TICK.COUNTER60_0_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__10253\,
            in1 => \N__10285\,
            in2 => \N__10430\,
            in3 => \N__10310\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10287\,
            in1 => \N__10256\,
            in2 => \N__10321\,
            in3 => \N__11057\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10559\,
            in1 => \N__10403\,
            in2 => \N__10448\,
            in3 => \N__11044\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10288\,
            in1 => \N__10257\,
            in2 => \N__10322\,
            in3 => \N__10628\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__10254\,
            in1 => \N__10289\,
            in2 => \N__10607\,
            in3 => \N__10317\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10425\,
            in2 => \_gnd_net_\,
            in3 => \N__10447\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__10595\,
            in1 => \N__11069\,
            in2 => \N__10544\,
            in3 => \N__10655\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10286\,
            in1 => \N__10255\,
            in2 => \N__10229\,
            in3 => \N__11078\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__10520\,
            in1 => \N__10226\,
            in2 => \_gnd_net_\,
            in3 => \N__10157\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__10214\,
            in1 => \N__10205\,
            in2 => \N__10193\,
            in3 => \N__10190\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11023\,
            in1 => \N__10932\,
            in2 => \N__10178\,
            in3 => \N__10175\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__10928\,
            in1 => \N__11024\,
            in2 => \N__10165\,
            in3 => \N__10983\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10981\,
            in1 => \N__10930\,
            in2 => \N__11033\,
            in3 => \N__10136\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10130\,
            in1 => \N__10118\,
            in2 => \N__10106\,
            in3 => \N__10891\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10982\,
            in1 => \N__10931\,
            in2 => \N__10091\,
            in3 => \N__10088\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__10929\,
            in1 => \N__10526\,
            in2 => \N__10994\,
            in3 => \N__11028\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10873\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__10460\,
            in1 => \N__10508\,
            in2 => \N__10496\,
            in3 => \N__10481\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11029\,
            in1 => \N__10988\,
            in2 => \N__10469\,
            in3 => \N__10466\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10875\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10443\,
            in2 => \N__10429\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_5_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10402\,
            in2 => \_gnd_net_\,
            in3 => \N__10391\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__10874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10384\,
            in2 => \_gnd_net_\,
            in3 => \N__10373\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__10874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10370\,
            in3 => \N__10343\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10336\,
            in2 => \_gnd_net_\,
            in3 => \N__10325\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__10874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_17_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10681\,
            in2 => \_gnd_net_\,
            in3 => \N__10658\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_17_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10654\,
            in2 => \_gnd_net_\,
            in3 => \N__10643\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__10874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_17_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10639\,
            in2 => \_gnd_net_\,
            in3 => \N__10622\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10618\,
            in2 => \_gnd_net_\,
            in3 => \N__10598\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_6_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10594\,
            in2 => \_gnd_net_\,
            in3 => \N__10583\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__10876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10573\,
            in2 => \_gnd_net_\,
            in3 => \N__10562\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__10876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10558\,
            in2 => \_gnd_net_\,
            in3 => \N__10547\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__10876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10540\,
            in2 => \_gnd_net_\,
            in3 => \N__10529\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__10876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11089\,
            in2 => \_gnd_net_\,
            in3 => \N__11072\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11068\,
            in2 => \_gnd_net_\,
            in3 => \N__11051\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11045\,
            in2 => \_gnd_net_\,
            in3 => \N__11048\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11030\,
            in1 => \N__10989\,
            in2 => \N__10941\,
            in3 => \N__10901\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10877\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PCS1_LC_20_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10804\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10766\,
            lcout => \PCS1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.SCS0_LC_20_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10767\,
            in2 => \_gnd_net_\,
            in3 => \N__10720\,
            lcout => \SCS0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PCS0_LC_22_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__10768\,
            in1 => \N__10805\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCS0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.SCS1_LC_22_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10769\,
            in2 => \_gnd_net_\,
            in3 => \N__10721\,
            lcout => \SCS1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_22_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \AGNUS_CLK_obuf_RNO_LC_24_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11153\,
            in1 => \N__11126\,
            in2 => \_gnd_net_\,
            in3 => \N__11114\,
            lcout => \AGNUS_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Sep 13 2025 21:18:13

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    ROM_DELAY,
    TM,
    TT,
    A,
    D,
    RESETn,
    OVL,
    CONFIGENn,
    PPIO,
    PORTSIZE,
    TICK60,
    PCS1,
    CIACS0n,
    SCS0,
    CPUCONFn,
    CLK6,
    AGNUS_CLK,
    CLK_CIA,
    BUFENn,
    AUTOBOOT,
    RnW,
    XCLK,
    CIACS1n,
    PPIO_J,
    TICK50,
    TCIn,
    TBIn,
    RAMSPACEn,
    PCS0,
    CLK40_IN,
    CLK28_IN,
    XCLK_ENn,
    SCS1,
    REGSPACEn,
    F_ENn,
    TSn,
    SPIO_J,
    SPIO,
    RTC_ENn,
    ATA_ENn,
    TACKn,
    ROMENn);

    input [1:0] ROM_DELAY;
    input [2:0] TM;
    input [1:0] TT;
    input [31:1] A;
    inout [7:4] D;
    input RESETn;
    input OVL;
    output CONFIGENn;
    output PPIO;
    output PORTSIZE;
    output TICK60;
    output PCS1;
    output CIACS0n;
    output SCS0;
    input CPUCONFn;
    input CLK6;
    output AGNUS_CLK;
    output CLK_CIA;
    output BUFENn;
    input AUTOBOOT;
    input RnW;
    input XCLK;
    output CIACS1n;
    input PPIO_J;
    output TICK50;
    output TCIn;
    output TBIn;
    output RAMSPACEn;
    output PCS0;
    input CLK40_IN;
    input CLK28_IN;
    input XCLK_ENn;
    output SCS1;
    output REGSPACEn;
    output F_ENn;
    input TSn;
    input SPIO_J;
    output SPIO;
    output RTC_ENn;
    output ATA_ENn;
    inout TACKn;
    output ROMENn;

    wire N__11620;
    wire N__11619;
    wire N__11618;
    wire N__11610;
    wire N__11609;
    wire N__11608;
    wire N__11600;
    wire N__11599;
    wire N__11598;
    wire N__11589;
    wire N__11588;
    wire N__11587;
    wire N__11580;
    wire N__11579;
    wire N__11578;
    wire N__11571;
    wire N__11570;
    wire N__11569;
    wire N__11562;
    wire N__11561;
    wire N__11560;
    wire N__11553;
    wire N__11552;
    wire N__11551;
    wire N__11544;
    wire N__11543;
    wire N__11542;
    wire N__11535;
    wire N__11534;
    wire N__11533;
    wire N__11526;
    wire N__11525;
    wire N__11524;
    wire N__11517;
    wire N__11516;
    wire N__11515;
    wire N__11508;
    wire N__11507;
    wire N__11506;
    wire N__11499;
    wire N__11498;
    wire N__11497;
    wire N__11490;
    wire N__11489;
    wire N__11488;
    wire N__11481;
    wire N__11480;
    wire N__11479;
    wire N__11472;
    wire N__11471;
    wire N__11470;
    wire N__11463;
    wire N__11462;
    wire N__11461;
    wire N__11454;
    wire N__11453;
    wire N__11452;
    wire N__11445;
    wire N__11444;
    wire N__11443;
    wire N__11436;
    wire N__11435;
    wire N__11434;
    wire N__11427;
    wire N__11426;
    wire N__11425;
    wire N__11418;
    wire N__11417;
    wire N__11416;
    wire N__11409;
    wire N__11408;
    wire N__11407;
    wire N__11400;
    wire N__11399;
    wire N__11398;
    wire N__11391;
    wire N__11390;
    wire N__11389;
    wire N__11382;
    wire N__11381;
    wire N__11380;
    wire N__11373;
    wire N__11372;
    wire N__11371;
    wire N__11364;
    wire N__11363;
    wire N__11362;
    wire N__11355;
    wire N__11354;
    wire N__11353;
    wire N__11346;
    wire N__11345;
    wire N__11344;
    wire N__11337;
    wire N__11336;
    wire N__11335;
    wire N__11328;
    wire N__11327;
    wire N__11326;
    wire N__11319;
    wire N__11318;
    wire N__11317;
    wire N__11310;
    wire N__11309;
    wire N__11308;
    wire N__11301;
    wire N__11300;
    wire N__11299;
    wire N__11292;
    wire N__11291;
    wire N__11290;
    wire N__11283;
    wire N__11282;
    wire N__11281;
    wire N__11274;
    wire N__11273;
    wire N__11272;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11256;
    wire N__11255;
    wire N__11254;
    wire N__11247;
    wire N__11246;
    wire N__11245;
    wire N__11238;
    wire N__11237;
    wire N__11236;
    wire N__11229;
    wire N__11228;
    wire N__11227;
    wire N__11220;
    wire N__11219;
    wire N__11218;
    wire N__11211;
    wire N__11210;
    wire N__11209;
    wire N__11202;
    wire N__11201;
    wire N__11200;
    wire N__11193;
    wire N__11192;
    wire N__11191;
    wire N__11184;
    wire N__11183;
    wire N__11182;
    wire N__11175;
    wire N__11174;
    wire N__11173;
    wire N__11166;
    wire N__11165;
    wire N__11164;
    wire N__11157;
    wire N__11156;
    wire N__11155;
    wire N__11148;
    wire N__11147;
    wire N__11146;
    wire N__11139;
    wire N__11138;
    wire N__11137;
    wire N__11130;
    wire N__11129;
    wire N__11128;
    wire N__11121;
    wire N__11120;
    wire N__11119;
    wire N__11112;
    wire N__11111;
    wire N__11110;
    wire N__11103;
    wire N__11102;
    wire N__11101;
    wire N__11094;
    wire N__11093;
    wire N__11092;
    wire N__11085;
    wire N__11084;
    wire N__11083;
    wire N__11076;
    wire N__11075;
    wire N__11074;
    wire N__11067;
    wire N__11066;
    wire N__11065;
    wire N__11058;
    wire N__11057;
    wire N__11056;
    wire N__11049;
    wire N__11048;
    wire N__11047;
    wire N__11040;
    wire N__11039;
    wire N__11038;
    wire N__11031;
    wire N__11030;
    wire N__11029;
    wire N__11022;
    wire N__11021;
    wire N__11020;
    wire N__11013;
    wire N__11012;
    wire N__11011;
    wire N__11004;
    wire N__11003;
    wire N__11002;
    wire N__10995;
    wire N__10994;
    wire N__10993;
    wire N__10976;
    wire N__10975;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10957;
    wire N__10956;
    wire N__10955;
    wire N__10948;
    wire N__10945;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10912;
    wire N__10911;
    wire N__10910;
    wire N__10909;
    wire N__10906;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10841;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10828;
    wire N__10825;
    wire N__10822;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10804;
    wire N__10801;
    wire N__10798;
    wire N__10793;
    wire N__10792;
    wire N__10791;
    wire N__10790;
    wire N__10789;
    wire N__10788;
    wire N__10787;
    wire N__10786;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10747;
    wire N__10744;
    wire N__10741;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10672;
    wire N__10669;
    wire N__10666;
    wire N__10663;
    wire N__10660;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10615;
    wire N__10612;
    wire N__10609;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10577;
    wire N__10574;
    wire N__10571;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10559;
    wire N__10556;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10534;
    wire N__10531;
    wire N__10528;
    wire N__10523;
    wire N__10520;
    wire N__10519;
    wire N__10516;
    wire N__10513;
    wire N__10508;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10487;
    wire N__10484;
    wire N__10483;
    wire N__10480;
    wire N__10477;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10462;
    wire N__10461;
    wire N__10458;
    wire N__10453;
    wire N__10448;
    wire N__10447;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10435;
    wire N__10434;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10420;
    wire N__10419;
    wire N__10414;
    wire N__10413;
    wire N__10412;
    wire N__10409;
    wire N__10408;
    wire N__10407;
    wire N__10406;
    wire N__10405;
    wire N__10404;
    wire N__10403;
    wire N__10402;
    wire N__10399;
    wire N__10398;
    wire N__10395;
    wire N__10394;
    wire N__10393;
    wire N__10390;
    wire N__10387;
    wire N__10384;
    wire N__10381;
    wire N__10378;
    wire N__10377;
    wire N__10376;
    wire N__10375;
    wire N__10374;
    wire N__10371;
    wire N__10368;
    wire N__10365;
    wire N__10364;
    wire N__10363;
    wire N__10362;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10318;
    wire N__10315;
    wire N__10306;
    wire N__10305;
    wire N__10302;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10281;
    wire N__10272;
    wire N__10271;
    wire N__10260;
    wire N__10255;
    wire N__10252;
    wire N__10247;
    wire N__10244;
    wire N__10239;
    wire N__10234;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10218;
    wire N__10215;
    wire N__10212;
    wire N__10209;
    wire N__10204;
    wire N__10201;
    wire N__10196;
    wire N__10189;
    wire N__10186;
    wire N__10183;
    wire N__10178;
    wire N__10175;
    wire N__10172;
    wire N__10171;
    wire N__10168;
    wire N__10165;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10148;
    wire N__10147;
    wire N__10146;
    wire N__10145;
    wire N__10142;
    wire N__10135;
    wire N__10130;
    wire N__10129;
    wire N__10128;
    wire N__10127;
    wire N__10126;
    wire N__10125;
    wire N__10124;
    wire N__10123;
    wire N__10122;
    wire N__10121;
    wire N__10120;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10090;
    wire N__10087;
    wire N__10084;
    wire N__10083;
    wire N__10078;
    wire N__10075;
    wire N__10070;
    wire N__10069;
    wire N__10066;
    wire N__10065;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10053;
    wire N__10050;
    wire N__10043;
    wire N__10042;
    wire N__10039;
    wire N__10036;
    wire N__10031;
    wire N__10028;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10016;
    wire N__10013;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10001;
    wire N__9998;
    wire N__9997;
    wire N__9994;
    wire N__9991;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9964;
    wire N__9961;
    wire N__9958;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9935;
    wire N__9934;
    wire N__9933;
    wire N__9932;
    wire N__9931;
    wire N__9928;
    wire N__9927;
    wire N__9924;
    wire N__9921;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9909;
    wire N__9906;
    wire N__9905;
    wire N__9904;
    wire N__9903;
    wire N__9900;
    wire N__9899;
    wire N__9898;
    wire N__9897;
    wire N__9896;
    wire N__9895;
    wire N__9892;
    wire N__9891;
    wire N__9890;
    wire N__9889;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9794;
    wire N__9793;
    wire N__9792;
    wire N__9791;
    wire N__9790;
    wire N__9789;
    wire N__9788;
    wire N__9781;
    wire N__9772;
    wire N__9767;
    wire N__9766;
    wire N__9765;
    wire N__9764;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9753;
    wire N__9750;
    wire N__9749;
    wire N__9748;
    wire N__9737;
    wire N__9730;
    wire N__9725;
    wire N__9724;
    wire N__9721;
    wire N__9720;
    wire N__9717;
    wire N__9716;
    wire N__9715;
    wire N__9714;
    wire N__9713;
    wire N__9712;
    wire N__9705;
    wire N__9694;
    wire N__9691;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9661;
    wire N__9660;
    wire N__9659;
    wire N__9658;
    wire N__9655;
    wire N__9652;
    wire N__9645;
    wire N__9638;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9625;
    wire N__9624;
    wire N__9623;
    wire N__9620;
    wire N__9619;
    wire N__9618;
    wire N__9617;
    wire N__9616;
    wire N__9607;
    wire N__9598;
    wire N__9593;
    wire N__9592;
    wire N__9591;
    wire N__9590;
    wire N__9589;
    wire N__9588;
    wire N__9587;
    wire N__9586;
    wire N__9585;
    wire N__9574;
    wire N__9565;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9533;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9521;
    wire N__9518;
    wire N__9517;
    wire N__9514;
    wire N__9511;
    wire N__9506;
    wire N__9503;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9491;
    wire N__9488;
    wire N__9487;
    wire N__9484;
    wire N__9483;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9445;
    wire N__9442;
    wire N__9439;
    wire N__9434;
    wire N__9433;
    wire N__9430;
    wire N__9427;
    wire N__9422;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9410;
    wire N__9409;
    wire N__9406;
    wire N__9405;
    wire N__9402;
    wire N__9399;
    wire N__9396;
    wire N__9389;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9341;
    wire N__9340;
    wire N__9339;
    wire N__9338;
    wire N__9337;
    wire N__9336;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9328;
    wire N__9319;
    wire N__9310;
    wire N__9305;
    wire N__9304;
    wire N__9303;
    wire N__9302;
    wire N__9299;
    wire N__9298;
    wire N__9297;
    wire N__9290;
    wire N__9287;
    wire N__9282;
    wire N__9275;
    wire N__9274;
    wire N__9273;
    wire N__9272;
    wire N__9269;
    wire N__9268;
    wire N__9267;
    wire N__9266;
    wire N__9263;
    wire N__9256;
    wire N__9253;
    wire N__9248;
    wire N__9239;
    wire N__9238;
    wire N__9237;
    wire N__9236;
    wire N__9235;
    wire N__9234;
    wire N__9227;
    wire N__9220;
    wire N__9215;
    wire N__9214;
    wire N__9213;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9205;
    wire N__9202;
    wire N__9199;
    wire N__9198;
    wire N__9191;
    wire N__9188;
    wire N__9183;
    wire N__9176;
    wire N__9175;
    wire N__9172;
    wire N__9171;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9101;
    wire N__9100;
    wire N__9097;
    wire N__9094;
    wire N__9091;
    wire N__9088;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9017;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8987;
    wire N__8986;
    wire N__8985;
    wire N__8982;
    wire N__8979;
    wire N__8976;
    wire N__8973;
    wire N__8966;
    wire N__8965;
    wire N__8962;
    wire N__8959;
    wire N__8956;
    wire N__8951;
    wire N__8948;
    wire N__8947;
    wire N__8944;
    wire N__8941;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8895;
    wire N__8890;
    wire N__8887;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8795;
    wire N__8794;
    wire N__8793;
    wire N__8792;
    wire N__8791;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8773;
    wire N__8762;
    wire N__8761;
    wire N__8760;
    wire N__8757;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8735;
    wire N__8734;
    wire N__8733;
    wire N__8730;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8705;
    wire N__8704;
    wire N__8703;
    wire N__8702;
    wire N__8701;
    wire N__8700;
    wire N__8697;
    wire N__8692;
    wire N__8687;
    wire N__8682;
    wire N__8675;
    wire N__8674;
    wire N__8673;
    wire N__8672;
    wire N__8671;
    wire N__8668;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8638;
    wire N__8637;
    wire N__8636;
    wire N__8635;
    wire N__8634;
    wire N__8629;
    wire N__8626;
    wire N__8623;
    wire N__8618;
    wire N__8609;
    wire N__8606;
    wire N__8605;
    wire N__8602;
    wire N__8599;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8578;
    wire N__8577;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8569;
    wire N__8566;
    wire N__8563;
    wire N__8558;
    wire N__8555;
    wire N__8550;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8518;
    wire N__8517;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8503;
    wire N__8500;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8461;
    wire N__8460;
    wire N__8457;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8443;
    wire N__8440;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8413;
    wire N__8412;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8390;
    wire N__8387;
    wire N__8386;
    wire N__8385;
    wire N__8384;
    wire N__8383;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8363;
    wire N__8360;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8327;
    wire N__8324;
    wire N__8323;
    wire N__8318;
    wire N__8315;
    wire N__8312;
    wire N__8309;
    wire N__8306;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8279;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8267;
    wire N__8266;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8233;
    wire N__8228;
    wire N__8227;
    wire N__8224;
    wire N__8221;
    wire N__8216;
    wire N__8215;
    wire N__8214;
    wire N__8213;
    wire N__8208;
    wire N__8203;
    wire N__8198;
    wire N__8197;
    wire N__8194;
    wire N__8193;
    wire N__8192;
    wire N__8189;
    wire N__8184;
    wire N__8181;
    wire N__8174;
    wire N__8173;
    wire N__8172;
    wire N__8167;
    wire N__8164;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8132;
    wire N__8131;
    wire N__8130;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8118;
    wire N__8111;
    wire N__8110;
    wire N__8109;
    wire N__8106;
    wire N__8101;
    wire N__8096;
    wire N__8093;
    wire N__8092;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8064;
    wire N__8061;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8044;
    wire N__8043;
    wire N__8042;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8034;
    wire N__8033;
    wire N__8028;
    wire N__8025;
    wire N__8020;
    wire N__8015;
    wire N__8006;
    wire N__8005;
    wire N__8002;
    wire N__8001;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7987;
    wire N__7980;
    wire N__7975;
    wire N__7970;
    wire N__7969;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7933;
    wire N__7930;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7900;
    wire N__7899;
    wire N__7898;
    wire N__7891;
    wire N__7888;
    wire N__7883;
    wire N__7882;
    wire N__7881;
    wire N__7878;
    wire N__7877;
    wire N__7876;
    wire N__7875;
    wire N__7872;
    wire N__7869;
    wire N__7866;
    wire N__7861;
    wire N__7858;
    wire N__7847;
    wire N__7846;
    wire N__7845;
    wire N__7844;
    wire N__7843;
    wire N__7840;
    wire N__7837;
    wire N__7832;
    wire N__7829;
    wire N__7820;
    wire N__7819;
    wire N__7818;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7806;
    wire N__7803;
    wire N__7800;
    wire N__7793;
    wire N__7792;
    wire N__7791;
    wire N__7790;
    wire N__7789;
    wire N__7782;
    wire N__7777;
    wire N__7772;
    wire N__7769;
    wire N__7768;
    wire N__7767;
    wire N__7762;
    wire N__7759;
    wire N__7754;
    wire N__7751;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7739;
    wire N__7736;
    wire N__7735;
    wire N__7732;
    wire N__7729;
    wire N__7724;
    wire N__7721;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7654;
    wire N__7653;
    wire N__7652;
    wire N__7651;
    wire N__7650;
    wire N__7647;
    wire N__7642;
    wire N__7639;
    wire N__7634;
    wire N__7625;
    wire N__7624;
    wire N__7623;
    wire N__7622;
    wire N__7621;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7613;
    wire N__7612;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7604;
    wire N__7601;
    wire N__7598;
    wire N__7595;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7579;
    wire N__7576;
    wire N__7575;
    wire N__7574;
    wire N__7569;
    wire N__7566;
    wire N__7561;
    wire N__7558;
    wire N__7555;
    wire N__7550;
    wire N__7547;
    wire N__7542;
    wire N__7539;
    wire N__7532;
    wire N__7525;
    wire N__7522;
    wire N__7519;
    wire N__7516;
    wire N__7513;
    wire N__7508;
    wire N__7505;
    wire N__7504;
    wire N__7503;
    wire N__7502;
    wire N__7501;
    wire N__7500;
    wire N__7497;
    wire N__7492;
    wire N__7489;
    wire N__7486;
    wire N__7483;
    wire N__7472;
    wire N__7469;
    wire N__7468;
    wire N__7465;
    wire N__7462;
    wire N__7461;
    wire N__7458;
    wire N__7455;
    wire N__7452;
    wire N__7445;
    wire N__7444;
    wire N__7441;
    wire N__7438;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7424;
    wire N__7421;
    wire N__7418;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7382;
    wire N__7379;
    wire N__7376;
    wire N__7373;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7360;
    wire N__7359;
    wire N__7358;
    wire N__7357;
    wire N__7356;
    wire N__7353;
    wire N__7348;
    wire N__7345;
    wire N__7342;
    wire N__7339;
    wire N__7328;
    wire N__7325;
    wire N__7322;
    wire N__7319;
    wire N__7316;
    wire N__7313;
    wire N__7312;
    wire N__7309;
    wire N__7306;
    wire N__7301;
    wire N__7298;
    wire N__7297;
    wire N__7296;
    wire N__7295;
    wire N__7294;
    wire N__7293;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7277;
    wire N__7268;
    wire N__7265;
    wire N__7264;
    wire N__7263;
    wire N__7260;
    wire N__7257;
    wire N__7256;
    wire N__7255;
    wire N__7254;
    wire N__7251;
    wire N__7250;
    wire N__7249;
    wire N__7248;
    wire N__7245;
    wire N__7242;
    wire N__7237;
    wire N__7234;
    wire N__7225;
    wire N__7214;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7199;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7187;
    wire N__7184;
    wire N__7181;
    wire N__7178;
    wire N__7175;
    wire N__7174;
    wire N__7173;
    wire N__7170;
    wire N__7167;
    wire N__7164;
    wire N__7157;
    wire N__7156;
    wire N__7153;
    wire N__7152;
    wire N__7149;
    wire N__7146;
    wire N__7143;
    wire N__7142;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7125;
    wire N__7124;
    wire N__7121;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7105;
    wire N__7104;
    wire N__7103;
    wire N__7102;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7084;
    wire N__7081;
    wire N__7070;
    wire N__7067;
    wire N__7066;
    wire N__7065;
    wire N__7064;
    wire N__7063;
    wire N__7062;
    wire N__7059;
    wire N__7058;
    wire N__7055;
    wire N__7050;
    wire N__7047;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7025;
    wire N__7024;
    wire N__7023;
    wire N__7020;
    wire N__7013;
    wire N__7012;
    wire N__7009;
    wire N__7006;
    wire N__7003;
    wire N__7000;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6985;
    wire N__6982;
    wire N__6979;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6953;
    wire N__6950;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6940;
    wire N__6935;
    wire N__6932;
    wire N__6931;
    wire N__6926;
    wire N__6923;
    wire N__6922;
    wire N__6919;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6909;
    wire N__6902;
    wire N__6901;
    wire N__6896;
    wire N__6895;
    wire N__6892;
    wire N__6889;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6874;
    wire N__6873;
    wire N__6870;
    wire N__6867;
    wire N__6864;
    wire N__6859;
    wire N__6858;
    wire N__6857;
    wire N__6856;
    wire N__6853;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6841;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6829;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6804;
    wire N__6801;
    wire N__6796;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6781;
    wire N__6780;
    wire N__6779;
    wire N__6778;
    wire N__6777;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6769;
    wire N__6768;
    wire N__6765;
    wire N__6764;
    wire N__6763;
    wire N__6762;
    wire N__6761;
    wire N__6760;
    wire N__6755;
    wire N__6750;
    wire N__6745;
    wire N__6740;
    wire N__6737;
    wire N__6732;
    wire N__6729;
    wire N__6724;
    wire N__6715;
    wire N__6712;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6694;
    wire N__6689;
    wire N__6686;
    wire N__6685;
    wire N__6680;
    wire N__6679;
    wire N__6678;
    wire N__6677;
    wire N__6676;
    wire N__6675;
    wire N__6674;
    wire N__6673;
    wire N__6672;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6657;
    wire N__6652;
    wire N__6647;
    wire N__6644;
    wire N__6643;
    wire N__6642;
    wire N__6631;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6614;
    wire N__6609;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6587;
    wire N__6586;
    wire N__6585;
    wire N__6584;
    wire N__6583;
    wire N__6582;
    wire N__6579;
    wire N__6578;
    wire N__6577;
    wire N__6576;
    wire N__6571;
    wire N__6566;
    wire N__6563;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6551;
    wire N__6546;
    wire N__6543;
    wire N__6540;
    wire N__6533;
    wire N__6532;
    wire N__6531;
    wire N__6530;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6512;
    wire N__6507;
    wire N__6494;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6484;
    wire N__6483;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6469;
    wire N__6468;
    wire N__6465;
    wire N__6462;
    wire N__6457;
    wire N__6456;
    wire N__6455;
    wire N__6452;
    wire N__6449;
    wire N__6442;
    wire N__6439;
    wire N__6434;
    wire N__6425;
    wire N__6424;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6377;
    wire N__6374;
    wire N__6373;
    wire N__6372;
    wire N__6365;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6296;
    wire N__6295;
    wire N__6290;
    wire N__6287;
    wire N__6286;
    wire N__6285;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6259;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6238;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6221;
    wire N__6218;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6185;
    wire N__6182;
    wire N__6181;
    wire N__6180;
    wire N__6179;
    wire N__6174;
    wire N__6171;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6119;
    wire N__6116;
    wire N__6113;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6103;
    wire N__6100;
    wire N__6099;
    wire N__6098;
    wire N__6097;
    wire N__6096;
    wire N__6095;
    wire N__6094;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6075;
    wire N__6072;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6041;
    wire N__6038;
    wire N__6037;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6016;
    wire N__6015;
    wire N__6014;
    wire N__6013;
    wire N__6010;
    wire N__6003;
    wire N__6002;
    wire N__6001;
    wire N__5998;
    wire N__5993;
    wire N__5990;
    wire N__5985;
    wire N__5980;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5965;
    wire N__5964;
    wire N__5961;
    wire N__5956;
    wire N__5955;
    wire N__5950;
    wire N__5949;
    wire N__5946;
    wire N__5945;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5931;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5894;
    wire N__5893;
    wire N__5890;
    wire N__5887;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5875;
    wire N__5872;
    wire N__5871;
    wire N__5868;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5854;
    wire N__5853;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5836;
    wire N__5835;
    wire N__5830;
    wire N__5827;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5808;
    wire N__5805;
    wire N__5800;
    wire N__5795;
    wire N__5794;
    wire N__5793;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5782;
    wire N__5781;
    wire N__5778;
    wire N__5777;
    wire N__5774;
    wire N__5773;
    wire N__5772;
    wire N__5771;
    wire N__5770;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5741;
    wire N__5740;
    wire N__5737;
    wire N__5732;
    wire N__5729;
    wire N__5726;
    wire N__5721;
    wire N__5714;
    wire N__5711;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5648;
    wire N__5647;
    wire N__5646;
    wire N__5645;
    wire N__5642;
    wire N__5641;
    wire N__5638;
    wire N__5635;
    wire N__5634;
    wire N__5633;
    wire N__5630;
    wire N__5623;
    wire N__5616;
    wire N__5613;
    wire N__5610;
    wire N__5603;
    wire N__5602;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5557;
    wire N__5556;
    wire N__5551;
    wire N__5548;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5522;
    wire N__5519;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5506;
    wire N__5505;
    wire N__5502;
    wire N__5499;
    wire N__5496;
    wire N__5493;
    wire N__5488;
    wire N__5487;
    wire N__5482;
    wire N__5479;
    wire N__5476;
    wire N__5473;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5459;
    wire N__5456;
    wire N__5453;
    wire N__5452;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5434;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5387;
    wire N__5384;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5372;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5319;
    wire N__5314;
    wire N__5311;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5272;
    wire N__5271;
    wire N__5270;
    wire N__5269;
    wire N__5266;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5233;
    wire N__5228;
    wire N__5225;
    wire N__5224;
    wire N__5221;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5210;
    wire N__5209;
    wire N__5206;
    wire N__5205;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5191;
    wire N__5188;
    wire N__5187;
    wire N__5186;
    wire N__5179;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5157;
    wire N__5154;
    wire N__5149;
    wire N__5146;
    wire N__5141;
    wire N__5138;
    wire N__5137;
    wire N__5136;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5128;
    wire N__5127;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5115;
    wire N__5110;
    wire N__5107;
    wire N__5106;
    wire N__5103;
    wire N__5094;
    wire N__5091;
    wire N__5088;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5072;
    wire N__5069;
    wire N__5068;
    wire N__5063;
    wire N__5062;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5052;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5033;
    wire N__5030;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4975;
    wire N__4972;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4942;
    wire N__4939;
    wire N__4936;
    wire N__4931;
    wire N__4928;
    wire N__4927;
    wire N__4924;
    wire N__4921;
    wire N__4916;
    wire N__4913;
    wire N__4912;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4902;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4879;
    wire N__4874;
    wire N__4873;
    wire N__4872;
    wire N__4869;
    wire N__4864;
    wire N__4863;
    wire N__4858;
    wire N__4855;
    wire N__4852;
    wire N__4849;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4828;
    wire N__4827;
    wire N__4824;
    wire N__4821;
    wire N__4818;
    wire N__4817;
    wire N__4816;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4791;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4777;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4750;
    wire N__4749;
    wire N__4744;
    wire N__4741;
    wire N__4740;
    wire N__4739;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4709;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4695;
    wire N__4692;
    wire N__4689;
    wire N__4682;
    wire N__4679;
    wire N__4678;
    wire N__4677;
    wire N__4672;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4662;
    wire N__4659;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4645;
    wire N__4642;
    wire N__4639;
    wire N__4634;
    wire N__4633;
    wire N__4628;
    wire N__4625;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4613;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4525;
    wire N__4522;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4504;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4483;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4450;
    wire N__4447;
    wire N__4444;
    wire N__4439;
    wire N__4436;
    wire N__4435;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4414;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4393;
    wire N__4390;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4366;
    wire N__4363;
    wire N__4360;
    wire N__4357;
    wire N__4354;
    wire N__4351;
    wire N__4348;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4291;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4249;
    wire N__4248;
    wire N__4247;
    wire N__4246;
    wire N__4245;
    wire N__4244;
    wire N__4243;
    wire N__4242;
    wire N__4241;
    wire N__4240;
    wire N__4239;
    wire N__4238;
    wire N__4211;
    wire CLK80_OUT;
    wire PPIO_c;
    wire GNDG0;
    wire SPIO_c;
    wire VCCG0;
    wire A_c_26;
    wire A_c_25;
    wire \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_3_cascade_ ;
    wire A_c_24;
    wire \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4 ;
    wire A_c_27;
    wire A_c_30;
    wire A_c_28;
    wire A_c_29;
    wire A_c_31;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_9 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_11_cascade_ ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_10 ;
    wire N_61_i;
    wire N_89_cascade_;
    wire N_94_cascade_;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3Z0Z_1 ;
    wire TT_c_0;
    wire TT_c_1;
    wire N_89;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_8 ;
    wire A_c_15;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_1_cascade_ ;
    wire A_c_16;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn_i;
    wire A_c_18;
    wire A_c_17;
    wire LIDE_BASE_1;
    wire \INVU409_AUTOCONFIG.LIDE_BASE_1C_net ;
    wire LIDE_BASE_4;
    wire LIDE_BASE_3;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4 ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2_cascade_ ;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1 ;
    wire ATA_SPACE_cascade_;
    wire \U409_ADDRESS_DECODE.ATA_ENZ0 ;
    wire \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1 ;
    wire OVL_c;
    wire A_c_19;
    wire \U409_ADDRESS_DECODE.Z2_SPACE ;
    wire \U409_ADDRESS_DECODE.N_34 ;
    wire \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_3 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACE_cascade_ ;
    wire \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_2 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_0Z0Z_2_cascade_ ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_4 ;
    wire \U409_AUTOCONFIG.N_227_3 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_4_cascade_ ;
    wire \U409_ADDRESS_DECODE.N_34_1 ;
    wire \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0Z0Z_0 ;
    wire N_100;
    wire N_94;
    wire \U409_AUTOCONFIG.PORTSIZEZ0Z_1_cascade_ ;
    wire PORTSIZE_0_i;
    wire \U409_AUTOCONFIG.un1_STATE_6_0_0 ;
    wire A_c_5;
    wire A_c_20;
    wire \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_1_cascade_ ;
    wire A_c_23;
    wire \U409_ADDRESS_DECODE.N_92 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACE_4 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACE_5 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACE_4_cascade_ ;
    wire \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_1 ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn_i;
    wire D_1_i;
    wire D_in_4;
    wire \U409_AUTOCONFIG.N_76 ;
    wire D_in_6;
    wire D_in_5;
    wire \U409_AUTOCONFIG.N_82 ;
    wire D_OUT_3;
    wire \U409_AUTOCONFIG.N_80 ;
    wire LIDE_BASE_2;
    wire LIDE_BASE_7;
    wire \U409_AUTOCONFIG.N_74 ;
    wire \INVU409_AUTOCONFIG.LIDE_BASE_2C_net ;
    wire A_c_22;
    wire A_c_21;
    wire LIDE_BASE_5;
    wire \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ;
    wire \U409_AUTOCONFIG.N_72 ;
    wire \U409_AUTOCONFIG.un1_STATE_6Z0Z_0 ;
    wire LIDE_BASE_6;
    wire \INVU409_AUTOCONFIG.LIDE_BASE_6C_net ;
    wire \U409_AUTOCONFIG.PR_OUTZ0Z_3 ;
    wire \U409_AUTOCONFIG.PR_OUT_cnst_i_0_2 ;
    wire \INVU409_AUTOCONFIG.PR_OUT_3C_net ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ;
    wire \INVU409_AUTOCONFIG.LIDE_OUT_3C_net ;
    wire \U409_AUTOCONFIG.N_225 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_3_cascade_ ;
    wire \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_3 ;
    wire A_c_6;
    wire A_c_7;
    wire \U409_AUTOCONFIG.un1_A_13Z0Z_3 ;
    wire \U409_AUTOCONFIG.un1_A_13Z0Z_0_cascade_ ;
    wire \U409_AUTOCONFIG.N_70 ;
    wire \U409_AUTOCONFIG.PR_OUTZ0Z_2 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2_cascade_ ;
    wire D_OUT_2;
    wire \U409_AUTOCONFIG.LIDE_BASE_10 ;
    wire D_in_7;
    wire \U409_AUTOCONFIG.LIDE_BASE_10_cascade_ ;
    wire \U409_AUTOCONFIG.N_78 ;
    wire \U409_AUTOCONFIG.LIDE_BASE_10_2 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNIOO061Z0Z_1_cascade_ ;
    wire D_OUT_1;
    wire \U409_AUTOCONFIG.LIDE_OUT_RNIMM061Z0Z_0_cascade_ ;
    wire D_OUT_0;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxaZ0Z_1 ;
    wire AUTOBOOT_c;
    wire \U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ;
    wire \U409_AUTOCONFIG.PR_OUTZ0Z_0 ;
    wire \U409_AUTOCONFIG.N_214_0 ;
    wire \U409_AUTOCONFIG.N_193_1 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ;
    wire \U409_AUTOCONFIG.N_159 ;
    wire \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_2 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ;
    wire \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ;
    wire \U409_AUTOCONFIG.N_192 ;
    wire \U409_AUTOCONFIG.PR_OUTZ0Z_1 ;
    wire \INVU409_AUTOCONFIG.LIDE_OUT_1C_net ;
    wire \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ;
    wire \U409_AUTOCONFIG.N_184_0 ;
    wire \U409_AUTOCONFIG.N_167 ;
    wire \U409_AUTOCONFIG.N_213_i ;
    wire \U409_AUTOCONFIG.N_182_0 ;
    wire \U409_AUTOCONFIG.N_223 ;
    wire \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_0_0 ;
    wire A_c_3;
    wire \U409_AUTOCONFIG.N_190 ;
    wire A_c_4;
    wire A_c_1;
    wire A_c_2;
    wire \U409_AUTOCONFIG.N_198 ;
    wire \U409_AUTOCONFIG.N_222 ;
    wire ATA_SPACE;
    wire BUFENn_c;
    wire \U409_AUTOCONFIG.D_OUT_sm0_0 ;
    wire CONFIGENn_c;
    wire \U409_AUTOCONFIG.LIDE_CONFZ0 ;
    wire \U409_AUTOCONFIG.BRIDGE_CONFZ0 ;
    wire \INVU409_AUTOCONFIG.CONFIGENnC_net ;
    wire \U409_AUTOCONFIG.STATE_d_2 ;
    wire \U409_AUTOCONFIG.un1_AZ0Z_13 ;
    wire \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1 ;
    wire \INVU409_AUTOCONFIG.STATE_0C_net ;
    wire AUTOCONFIG_SPACE;
    wire CONFIGURED;
    wire CPUCONFn_c;
    wire \U409_AUTOCONFIG.AC_STARTZ0 ;
    wire \U409_AUTOCONFIG.STATE4 ;
    wire \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_0 ;
    wire \U409_AUTOCONFIG.STATEZ0Z_0 ;
    wire RnW_c;
    wire \U409_AUTOCONFIG.STATEZ0Z_1 ;
    wire \INVU409_AUTOCONFIG.AC_TACKC_net ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn;
    wire TACKn_in;
    wire \U409_TRANSFER_ACK.N_53 ;
    wire \U409_TRANSFER_ACK.N_53_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ;
    wire \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire AC_TACK;
    wire \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a3_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ;
    wire GB_BUFFER_CLK40_IN_c_g_THRU_CO;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6 ;
    wire TACK_OUT;
    wire \INVU409_TRANSFER_ACK.TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.N_62 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire RESETn_c_i;
    wire \U409_CIA.CLK_CIA6_3_cascade_ ;
    wire \U409_CIA.un1_CIA_CLK_COUNT_2_1 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_0 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNT11_3 ;
    wire \U409_CIA.CLK_CIA6_0_cascade_ ;
    wire \U409_CIA.CLK_CIA6_3 ;
    wire \U409_CIA.CLK_CIA6_cascade_ ;
    wire \U409_CIA.CLK_CIA_RNOZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ;
    wire TSn_c;
    wire CIA_ENABLE_cascade_;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire CIA_ENABLE;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire bfn_14_9_0_;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_6 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_6 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_7 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.CLK_CIA6_0 ;
    wire \U409_CIA.un1_CIA_CLK_COUNT_3_1_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire CIA_SPACE;
    wire \U409_CIA.VMA_RNOZ0Z_0_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_5_0_0 ;
    wire \U409_TRANSFER_ACK.N_19_cascade_ ;
    wire \U409_TRANSFER_ACK.N_23 ;
    wire \U409_TRANSFER_ACK.N_22 ;
    wire ROMENn_c;
    wire \INVU409_TRANSFER_ACK.ROMENnC_net ;
    wire bfn_15_7_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire bfn_15_8_0_;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_0C_net ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.N_101 ;
    wire \U409_TRANSFER_ACK.N_19 ;
    wire CLK_CIA_c;
    wire \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ;
    wire ROMEN;
    wire TACK_EN;
    wire TCIn_1_i;
    wire TICK50_c;
    wire \U409_TICK.TICK503_11 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire TICK60_c;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.TICK603_8_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.TICK603_11 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire CLK40_IN_c_g;
    wire \U409_TRANSFER_ACK.N_17_mux ;
    wire \U409_TRANSFER_ACK.N_17_mux_cascade_ ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0 ;
    wire \U409_TRANSFER_ACK.N_3_0_cascade_ ;
    wire \U409_TRANSFER_ACK.N_6_0 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_10 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_3_0 ;
    wire \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire RESETn_c;
    wire \U409_CIA.VMAZ0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.LASTCLK_1C_net ;
    wire RESETn_c_i_g;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire bfn_17_6_0_;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire bfn_17_7_0_;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire CLK6_c_g;
    wire CONSTANT_ONE_NET;
    wire U409_ADDRESS_DECODE_un1_ATA_ENn;
    wire U409_ADDRESS_DECODE_un1_ATA_ENn_i;
    wire PCS1_c;
    wire \U409_ADDRESS_DECODE.CSZ0Z0 ;
    wire PCS0_c;
    wire SCS0_c;
    wire \U409_ADDRESS_DECODE.CSZ0Z1 ;
    wire A_c_14;
    wire SCS1_c;
    wire CLK28_IN_c_g;
    wire XCLK_c;
    wire XCLK_ENn_c;
    wire AGNUS_CLK_c;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__7754),
            .RESETB(N__10763),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11618),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__11620),
            .DIN(N__11619),
            .DOUT(N__11618),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__11620),
            .PADOUT(N__11619),
            .PADIN(N__11618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK40_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11608),
            .GLOBALBUFFEROUTPUT(CLK40_IN_c_g));
    IO_PAD CLK40_IN_ibuf_gb_io_iopad (
            .OE(N__11610),
            .DIN(N__11609),
            .DOUT(N__11608),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_gb_io_preio (
            .PADOEN(N__11610),
            .PADOUT(N__11609),
            .PADIN(N__11608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__11598),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__11600),
            .DIN(N__11599),
            .DOUT(N__11598),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__11600),
            .PADOUT(N__11599),
            .PADIN(N__11598),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11589),
            .DIN(N__11588),
            .DOUT(N__11587),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11589),
            .PADOUT(N__11588),
            .PADIN(N__11587),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__11580),
            .DIN(N__11579),
            .DOUT(N__11578),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__11580),
            .PADOUT(N__11579),
            .PADIN(N__11578),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_7_iopad (
            .OE(N__11571),
            .DIN(N__11570),
            .DOUT(N__11569),
            .PACKAGEPIN(D[7]));
    defparam D_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_7_preio (
            .PADOEN(N__11571),
            .PADOUT(N__11570),
            .PADIN(N__11569),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5510),
            .DIN0(D_in_7),
            .DOUT0(N__5411),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11562),
            .DIN(N__11561),
            .DOUT(N__11560),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11562),
            .PADOUT(N__11561),
            .PADIN(N__11560),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CPUCONFn_ibuf_iopad (
            .OE(N__11553),
            .DIN(N__11552),
            .DOUT(N__11551),
            .PACKAGEPIN(CPUCONFn));
    defparam CPUCONFn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CPUCONFn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CPUCONFn_ibuf_preio (
            .PADOEN(N__11553),
            .PADOUT(N__11552),
            .PADIN(N__11551),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CPUCONFn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RTC_ENn_obuf_iopad (
            .OE(N__11544),
            .DIN(N__11543),
            .DOUT(N__11542),
            .PACKAGEPIN(RTC_ENn));
    defparam RTC_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RTC_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RTC_ENn_obuf_preio (
            .PADOEN(N__11544),
            .PADOUT(N__11543),
            .PADIN(N__11542),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4322),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__11535),
            .DIN(N__11534),
            .DOUT(N__11533),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__11535),
            .PADOUT(N__11534),
            .PADIN(N__11533),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SPIO_J_ibuf_iopad.PULLUP=1'b1;
    IO_PAD SPIO_J_ibuf_iopad (
            .OE(N__11526),
            .DIN(N__11525),
            .DOUT(N__11524),
            .PACKAGEPIN(SPIO_J));
    defparam SPIO_J_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SPIO_J_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SPIO_J_ibuf_preio (
            .PADOEN(N__11526),
            .PADOUT(N__11525),
            .PADIN(N__11524),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SPIO_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_4_iopad (
            .OE(N__11517),
            .DIN(N__11516),
            .DOUT(N__11515),
            .PACKAGEPIN(D[4]));
    defparam D_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_4_preio (
            .PADOEN(N__11517),
            .PADOUT(N__11516),
            .PADIN(N__11515),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5487),
            .DIN0(D_in_4),
            .DOUT0(N__6410),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PPIO_obuf_iopad (
            .OE(N__11508),
            .DIN(N__11507),
            .DOUT(N__11506),
            .PACKAGEPIN(PPIO));
    defparam PPIO_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PPIO_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PPIO_obuf_preio (
            .PADOEN(N__11508),
            .PADOUT(N__11507),
            .PADIN(N__11506),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4271),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11499),
            .DIN(N__11498),
            .DOUT(N__11497),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11499),
            .PADOUT(N__11498),
            .PADIN(N__11497),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__11490),
            .DIN(N__11489),
            .DOUT(N__11488),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__11490),
            .PADOUT(N__11489),
            .PADIN(N__11488),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam PPIO_J_ibuf_iopad.PULLUP=1'b1;
    IO_PAD PPIO_J_ibuf_iopad (
            .OE(N__11481),
            .DIN(N__11480),
            .DOUT(N__11479),
            .PACKAGEPIN(PPIO_J));
    defparam PPIO_J_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam PPIO_J_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO PPIO_J_ibuf_preio (
            .PADOEN(N__11481),
            .PADOUT(N__11480),
            .PADIN(N__11479),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(PPIO_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__11472),
            .DIN(N__11471),
            .DOUT(N__11470),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__11472),
            .PADOUT(N__11471),
            .PADIN(N__11470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4772),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11463),
            .DIN(N__11462),
            .DOUT(N__11461),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11463),
            .PADOUT(N__11462),
            .PADIN(N__11461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__11454),
            .DIN(N__11453),
            .DOUT(N__11452),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__11454),
            .PADOUT(N__11453),
            .PADIN(N__11452),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8840),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__11445),
            .DIN(N__11444),
            .DOUT(N__11443),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__11445),
            .PADOUT(N__11444),
            .PADIN(N__11443),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9137),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam AUTOBOOT_ibuf_iopad.PULLUP=1'b1;
    IO_PAD AUTOBOOT_ibuf_iopad (
            .OE(N__11436),
            .DIN(N__11435),
            .DOUT(N__11434),
            .PACKAGEPIN(AUTOBOOT));
    defparam AUTOBOOT_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AUTOBOOT_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AUTOBOOT_ibuf_preio (
            .PADOEN(N__11436),
            .PADOUT(N__11435),
            .PADIN(N__11434),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AUTOBOOT_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11427),
            .DIN(N__11426),
            .DOUT(N__11425),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11427),
            .PADOUT(N__11426),
            .PADIN(N__11425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__11418),
            .DIN(N__11417),
            .DOUT(N__11416),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__11418),
            .PADOUT(N__11417),
            .PADIN(N__11416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5303),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD F_ENn_obuf_iopad (
            .OE(N__11409),
            .DIN(N__11408),
            .DOUT(N__11407),
            .PACKAGEPIN(F_ENn));
    defparam F_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam F_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO F_ENn_obuf_preio (
            .PADOEN(N__11409),
            .PADOUT(N__11408),
            .PADIN(N__11407),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10762),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11400),
            .DIN(N__11399),
            .DOUT(N__11398),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11400),
            .PADOUT(N__11399),
            .PADIN(N__11398),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__11391),
            .DIN(N__11390),
            .DOUT(N__11389),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__11391),
            .PADOUT(N__11390),
            .PADIN(N__11389),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11382),
            .DIN(N__11381),
            .DOUT(N__11380),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11382),
            .PADOUT(N__11381),
            .PADIN(N__11380),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11373),
            .DIN(N__11372),
            .DOUT(N__11371),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11373),
            .PADOUT(N__11372),
            .PADIN(N__11371),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11364),
            .DIN(N__11363),
            .DOUT(N__11362),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11364),
            .PADOUT(N__11363),
            .PADIN(N__11362),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SCS1_obuf_iopad (
            .OE(N__11355),
            .DIN(N__11354),
            .DOUT(N__11353),
            .PACKAGEPIN(SCS1));
    defparam SCS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SCS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SCS1_obuf_preio (
            .PADOEN(N__11355),
            .PADOUT(N__11354),
            .PADIN(N__11353),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10928),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_CLK_obuf_iopad (
            .OE(N__11346),
            .DIN(N__11345),
            .DOUT(N__11344),
            .PACKAGEPIN(AGNUS_CLK));
    defparam AGNUS_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO AGNUS_CLK_obuf_preio (
            .PADOEN(N__11346),
            .PADOUT(N__11345),
            .PADIN(N__11344),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10865),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__11337),
            .DIN(N__11336),
            .DOUT(N__11335),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__11337),
            .PADOUT(N__11336),
            .PADIN(N__11335),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__11328),
            .DIN(N__11327),
            .DOUT(N__11326),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__11328),
            .PADOUT(N__11327),
            .PADIN(N__11326),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8492),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__11319),
            .DIN(N__11318),
            .DOUT(N__11317),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__11319),
            .PADOUT(N__11318),
            .PADIN(N__11317),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9062),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11310),
            .DIN(N__11309),
            .DOUT(N__11308),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11310),
            .PADOUT(N__11309),
            .PADIN(N__11308),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__11301),
            .DIN(N__11300),
            .DOUT(N__11299),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__11301),
            .PADOUT(N__11300),
            .PADIN(N__11299),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__11292),
            .DIN(N__11291),
            .DOUT(N__11290),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__11292),
            .PADOUT(N__11291),
            .PADIN(N__11290),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__11283),
            .DIN(N__11282),
            .DOUT(N__11281),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__11283),
            .PADOUT(N__11282),
            .PADIN(N__11281),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__11274),
            .DIN(N__11273),
            .DOUT(N__11272),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__11274),
            .PADOUT(N__11273),
            .PADIN(N__11272),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9083),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_5_iopad (
            .OE(N__11265),
            .DIN(N__11264),
            .DOUT(N__11263),
            .PACKAGEPIN(D[5]));
    defparam D_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_5_preio (
            .PADOEN(N__11265),
            .PADOUT(N__11264),
            .PADIN(N__11263),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5505),
            .DIN0(D_in_5),
            .DOUT0(N__6056),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD XCLK_ENn_ibuf_iopad (
            .OE(N__11256),
            .DIN(N__11255),
            .DOUT(N__11254),
            .PACKAGEPIN(XCLK_ENn));
    defparam XCLK_ENn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam XCLK_ENn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO XCLK_ENn_ibuf_preio (
            .PADOEN(N__11256),
            .PADOUT(N__11255),
            .PADIN(N__11254),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(XCLK_ENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11247),
            .DIN(N__11246),
            .DOUT(N__11245),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11247),
            .PADOUT(N__11246),
            .PADIN(N__11245),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11238),
            .DIN(N__11237),
            .DOUT(N__11236),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11238),
            .PADOUT(N__11237),
            .PADIN(N__11236),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11229),
            .DIN(N__11228),
            .DOUT(N__11227),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11229),
            .PADOUT(N__11228),
            .PADIN(N__11227),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CONFIGENn_obuf_iopad (
            .OE(N__11220),
            .DIN(N__11219),
            .DOUT(N__11218),
            .PACKAGEPIN(CONFIGENn));
    defparam CONFIGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CONFIGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CONFIGENn_obuf_preio (
            .PADOEN(N__11220),
            .PADOUT(N__11219),
            .PADIN(N__11218),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7328),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SPIO_obuf_iopad (
            .OE(N__11211),
            .DIN(N__11210),
            .DOUT(N__11209),
            .PACKAGEPIN(SPIO));
    defparam SPIO_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SPIO_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SPIO_obuf_preio (
            .PADOEN(N__11211),
            .PADOUT(N__11210),
            .PADIN(N__11209),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4307),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__11202),
            .DIN(N__11201),
            .DOUT(N__11200),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__11202),
            .PADOUT(N__11201),
            .PADIN(N__11200),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9557),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__11193),
            .DIN(N__11192),
            .DOUT(N__11191),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__11193),
            .PADOUT(N__11192),
            .PADIN(N__11191),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__11184),
            .DIN(N__11183),
            .DOUT(N__11182),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__11184),
            .PADOUT(N__11183),
            .PADIN(N__11182),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11175),
            .DIN(N__11174),
            .DOUT(N__11173),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11175),
            .PADOUT(N__11174),
            .PADIN(N__11173),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ATA_ENn_obuf_iopad (
            .OE(N__11166),
            .DIN(N__11165),
            .DOUT(N__11164),
            .PACKAGEPIN(ATA_ENn));
    defparam ATA_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ATA_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ATA_ENn_obuf_preio (
            .PADOEN(N__11166),
            .PADOUT(N__11165),
            .PADIN(N__11164),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10700),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__11157),
            .DIN(N__11156),
            .DOUT(N__11155),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__11157),
            .PADOUT(N__11156),
            .PADIN(N__11155),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__11148),
            .DIN(N__11147),
            .DOUT(N__11146),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__11148),
            .PADOUT(N__11147),
            .PADIN(N__11146),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8435),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__11139),
            .DIN(N__11138),
            .DOUT(N__11137),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__11139),
            .PADOUT(N__11138),
            .PADIN(N__11137),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5534),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCS0_obuf_iopad (
            .OE(N__11130),
            .DIN(N__11129),
            .DOUT(N__11128),
            .PACKAGEPIN(PCS0));
    defparam PCS0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PCS0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PCS0_obuf_preio (
            .PADOEN(N__11130),
            .PADOUT(N__11129),
            .PADIN(N__11128),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10649),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11121),
            .DIN(N__11120),
            .DOUT(N__11119),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11121),
            .PADOUT(N__11120),
            .PADIN(N__11119),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_CIA_obuf_iopad (
            .OE(N__11112),
            .DIN(N__11111),
            .DOUT(N__11110),
            .PACKAGEPIN(CLK_CIA));
    defparam CLK_CIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_CIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_CIA_obuf_preio (
            .PADOEN(N__11112),
            .PADOUT(N__11111),
            .PADIN(N__11110),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8918),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11103),
            .DIN(N__11102),
            .DOUT(N__11101),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11103),
            .PADOUT(N__11102),
            .PADIN(N__11101),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCS1_obuf_iopad (
            .OE(N__11094),
            .DIN(N__11093),
            .DOUT(N__11092),
            .PACKAGEPIN(PCS1));
    defparam PCS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PCS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PCS1_obuf_preio (
            .PADOEN(N__11094),
            .PADOUT(N__11093),
            .PADIN(N__11092),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10691),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__11085),
            .DIN(N__11084),
            .DOUT(N__11083),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__11085),
            .PADOUT(N__11084),
            .PADIN(N__11083),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__9133),
            .DIN0(TACKn_in),
            .DOUT0(N__8159),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__11076),
            .DIN(N__11075),
            .DOUT(N__11074),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__11076),
            .PADOUT(N__11075),
            .PADIN(N__11074),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__11067),
            .DIN(N__11066),
            .DOUT(N__11065),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__11067),
            .PADOUT(N__11066),
            .PADIN(N__11065),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7382),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__11058),
            .DIN(N__11057),
            .DOUT(N__11056),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__11058),
            .PADOUT(N__11057),
            .PADIN(N__11056),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_iobuf_6_iopad (
            .OE(N__11049),
            .DIN(N__11048),
            .DOUT(N__11047),
            .PACKAGEPIN(D[6]));
    defparam D_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam D_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_iobuf_6_preio (
            .PADOEN(N__11049),
            .PADOUT(N__11048),
            .PADIN(N__11047),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5506),
            .DIN0(D_in_6),
            .DOUT0(N__6194),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11040),
            .DIN(N__11039),
            .DOUT(N__11038),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11040),
            .PADOUT(N__11039),
            .PADIN(N__11038),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__11031),
            .DIN(N__11030),
            .DOUT(N__11029),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__11031),
            .PADOUT(N__11030),
            .PADIN(N__11029),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SCS0_obuf_iopad (
            .OE(N__11022),
            .DIN(N__11021),
            .DOUT(N__11020),
            .PACKAGEPIN(SCS0));
    defparam SCS0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SCS0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SCS0_obuf_preio (
            .PADOEN(N__11022),
            .PADOUT(N__11021),
            .PADIN(N__11020),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10634),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD XCLK_ibuf_iopad (
            .OE(N__11013),
            .DIN(N__11012),
            .DOUT(N__11011),
            .PACKAGEPIN(XCLK));
    defparam XCLK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam XCLK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO XCLK_ibuf_preio (
            .PADOEN(N__11013),
            .PADOUT(N__11012),
            .PADIN(N__11011),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(XCLK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11004),
            .DIN(N__11003),
            .DOUT(N__11002),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11004),
            .PADOUT(N__11003),
            .PADIN(N__11002),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__10995),
            .DIN(N__10994),
            .DOUT(N__10993),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__10995),
            .PADOUT(N__10994),
            .PADIN(N__10993),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2625 (
            .O(N__10976),
            .I(N__10970));
    InMux I__2624 (
            .O(N__10975),
            .I(N__10970));
    LocalMux I__2623 (
            .O(N__10970),
            .I(N__10967));
    Sp12to4 I__2622 (
            .O(N__10967),
            .I(N__10964));
    Span12Mux_h I__2621 (
            .O(N__10964),
            .I(N__10961));
    Odrv12 I__2620 (
            .O(N__10961),
            .I(\U409_ADDRESS_DECODE.CSZ0Z1 ));
    InMux I__2619 (
            .O(N__10958),
            .I(N__10948));
    InMux I__2618 (
            .O(N__10957),
            .I(N__10948));
    InMux I__2617 (
            .O(N__10956),
            .I(N__10948));
    InMux I__2616 (
            .O(N__10955),
            .I(N__10945));
    LocalMux I__2615 (
            .O(N__10948),
            .I(N__10940));
    LocalMux I__2614 (
            .O(N__10945),
            .I(N__10940));
    Span12Mux_v I__2613 (
            .O(N__10940),
            .I(N__10937));
    Span12Mux_h I__2612 (
            .O(N__10937),
            .I(N__10934));
    Span12Mux_h I__2611 (
            .O(N__10934),
            .I(N__10931));
    Odrv12 I__2610 (
            .O(N__10931),
            .I(A_c_14));
    IoInMux I__2609 (
            .O(N__10928),
            .I(N__10925));
    LocalMux I__2608 (
            .O(N__10925),
            .I(N__10922));
    Span12Mux_s4_h I__2607 (
            .O(N__10922),
            .I(N__10919));
    Odrv12 I__2606 (
            .O(N__10919),
            .I(SCS1_c));
    InMux I__2605 (
            .O(N__10916),
            .I(N__10913));
    LocalMux I__2604 (
            .O(N__10913),
            .I(N__10906));
    ClkMux I__2603 (
            .O(N__10912),
            .I(N__10895));
    ClkMux I__2602 (
            .O(N__10911),
            .I(N__10895));
    ClkMux I__2601 (
            .O(N__10910),
            .I(N__10895));
    ClkMux I__2600 (
            .O(N__10909),
            .I(N__10895));
    Glb2LocalMux I__2599 (
            .O(N__10906),
            .I(N__10895));
    GlobalMux I__2598 (
            .O(N__10895),
            .I(N__10892));
    gio2CtrlBuf I__2597 (
            .O(N__10892),
            .I(CLK28_IN_c_g));
    InMux I__2596 (
            .O(N__10889),
            .I(N__10886));
    LocalMux I__2595 (
            .O(N__10886),
            .I(N__10883));
    Span4Mux_v I__2594 (
            .O(N__10883),
            .I(N__10880));
    Odrv4 I__2593 (
            .O(N__10880),
            .I(XCLK_c));
    InMux I__2592 (
            .O(N__10877),
            .I(N__10874));
    LocalMux I__2591 (
            .O(N__10874),
            .I(N__10871));
    Span12Mux_v I__2590 (
            .O(N__10871),
            .I(N__10868));
    Odrv12 I__2589 (
            .O(N__10868),
            .I(XCLK_ENn_c));
    IoInMux I__2588 (
            .O(N__10865),
            .I(N__10862));
    LocalMux I__2587 (
            .O(N__10862),
            .I(N__10859));
    Span4Mux_s3_h I__2586 (
            .O(N__10859),
            .I(N__10856));
    Odrv4 I__2585 (
            .O(N__10856),
            .I(AGNUS_CLK_c));
    InMux I__2584 (
            .O(N__10853),
            .I(N__10849));
    InMux I__2583 (
            .O(N__10852),
            .I(N__10846));
    LocalMux I__2582 (
            .O(N__10849),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__2581 (
            .O(N__10846),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    CascadeMux I__2580 (
            .O(N__10841),
            .I(N__10838));
    InMux I__2579 (
            .O(N__10838),
            .I(N__10835));
    LocalMux I__2578 (
            .O(N__10835),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    InMux I__2577 (
            .O(N__10832),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__2576 (
            .O(N__10829),
            .I(N__10825));
    InMux I__2575 (
            .O(N__10828),
            .I(N__10822));
    LocalMux I__2574 (
            .O(N__10825),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__2573 (
            .O(N__10822),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    InMux I__2572 (
            .O(N__10817),
            .I(N__10814));
    LocalMux I__2571 (
            .O(N__10814),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__2570 (
            .O(N__10811),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__2569 (
            .O(N__10808),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    InMux I__2568 (
            .O(N__10805),
            .I(N__10801));
    InMux I__2567 (
            .O(N__10804),
            .I(N__10798));
    LocalMux I__2566 (
            .O(N__10801),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__2565 (
            .O(N__10798),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    ClkMux I__2564 (
            .O(N__10793),
            .I(N__10769));
    ClkMux I__2563 (
            .O(N__10792),
            .I(N__10769));
    ClkMux I__2562 (
            .O(N__10791),
            .I(N__10769));
    ClkMux I__2561 (
            .O(N__10790),
            .I(N__10769));
    ClkMux I__2560 (
            .O(N__10789),
            .I(N__10769));
    ClkMux I__2559 (
            .O(N__10788),
            .I(N__10769));
    ClkMux I__2558 (
            .O(N__10787),
            .I(N__10769));
    ClkMux I__2557 (
            .O(N__10786),
            .I(N__10769));
    GlobalMux I__2556 (
            .O(N__10769),
            .I(N__10766));
    gio2CtrlBuf I__2555 (
            .O(N__10766),
            .I(CLK6_c_g));
    IoInMux I__2554 (
            .O(N__10763),
            .I(N__10759));
    IoInMux I__2553 (
            .O(N__10762),
            .I(N__10756));
    LocalMux I__2552 (
            .O(N__10759),
            .I(N__10753));
    LocalMux I__2551 (
            .O(N__10756),
            .I(N__10750));
    IoSpan4Mux I__2550 (
            .O(N__10753),
            .I(N__10747));
    IoSpan4Mux I__2549 (
            .O(N__10750),
            .I(N__10744));
    Sp12to4 I__2548 (
            .O(N__10747),
            .I(N__10741));
    Span4Mux_s2_h I__2547 (
            .O(N__10744),
            .I(N__10738));
    Span12Mux_s9_v I__2546 (
            .O(N__10741),
            .I(N__10735));
    Span4Mux_h I__2545 (
            .O(N__10738),
            .I(N__10732));
    Odrv12 I__2544 (
            .O(N__10735),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2543 (
            .O(N__10732),
            .I(CONSTANT_ONE_NET));
    InMux I__2542 (
            .O(N__10727),
            .I(N__10724));
    LocalMux I__2541 (
            .O(N__10724),
            .I(N__10721));
    Span4Mux_v I__2540 (
            .O(N__10721),
            .I(N__10718));
    Span4Mux_h I__2539 (
            .O(N__10718),
            .I(N__10714));
    InMux I__2538 (
            .O(N__10717),
            .I(N__10711));
    Sp12to4 I__2537 (
            .O(N__10714),
            .I(N__10708));
    LocalMux I__2536 (
            .O(N__10711),
            .I(N__10705));
    Odrv12 I__2535 (
            .O(N__10708),
            .I(U409_ADDRESS_DECODE_un1_ATA_ENn));
    Odrv4 I__2534 (
            .O(N__10705),
            .I(U409_ADDRESS_DECODE_un1_ATA_ENn));
    IoInMux I__2533 (
            .O(N__10700),
            .I(N__10697));
    LocalMux I__2532 (
            .O(N__10697),
            .I(N__10694));
    Odrv12 I__2531 (
            .O(N__10694),
            .I(U409_ADDRESS_DECODE_un1_ATA_ENn_i));
    IoInMux I__2530 (
            .O(N__10691),
            .I(N__10688));
    LocalMux I__2529 (
            .O(N__10688),
            .I(N__10685));
    IoSpan4Mux I__2528 (
            .O(N__10685),
            .I(N__10682));
    Span4Mux_s3_h I__2527 (
            .O(N__10682),
            .I(N__10679));
    Odrv4 I__2526 (
            .O(N__10679),
            .I(PCS1_c));
    InMux I__2525 (
            .O(N__10676),
            .I(N__10673));
    LocalMux I__2524 (
            .O(N__10673),
            .I(N__10669));
    InMux I__2523 (
            .O(N__10672),
            .I(N__10666));
    Sp12to4 I__2522 (
            .O(N__10669),
            .I(N__10663));
    LocalMux I__2521 (
            .O(N__10666),
            .I(N__10660));
    Span12Mux_v I__2520 (
            .O(N__10663),
            .I(N__10655));
    Sp12to4 I__2519 (
            .O(N__10660),
            .I(N__10655));
    Span12Mux_h I__2518 (
            .O(N__10655),
            .I(N__10652));
    Odrv12 I__2517 (
            .O(N__10652),
            .I(\U409_ADDRESS_DECODE.CSZ0Z0 ));
    IoInMux I__2516 (
            .O(N__10649),
            .I(N__10646));
    LocalMux I__2515 (
            .O(N__10646),
            .I(N__10643));
    Span4Mux_s3_h I__2514 (
            .O(N__10643),
            .I(N__10640));
    Span4Mux_v I__2513 (
            .O(N__10640),
            .I(N__10637));
    Odrv4 I__2512 (
            .O(N__10637),
            .I(PCS0_c));
    IoInMux I__2511 (
            .O(N__10634),
            .I(N__10631));
    LocalMux I__2510 (
            .O(N__10631),
            .I(N__10628));
    Span4Mux_s3_h I__2509 (
            .O(N__10628),
            .I(N__10625));
    Span4Mux_v I__2508 (
            .O(N__10625),
            .I(N__10622));
    Odrv4 I__2507 (
            .O(N__10622),
            .I(SCS0_c));
    CascadeMux I__2506 (
            .O(N__10619),
            .I(N__10616));
    InMux I__2505 (
            .O(N__10616),
            .I(N__10612));
    InMux I__2504 (
            .O(N__10615),
            .I(N__10609));
    LocalMux I__2503 (
            .O(N__10612),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__2502 (
            .O(N__10609),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    CascadeMux I__2501 (
            .O(N__10604),
            .I(N__10601));
    InMux I__2500 (
            .O(N__10601),
            .I(N__10598));
    LocalMux I__2499 (
            .O(N__10598),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__2498 (
            .O(N__10595),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    CascadeMux I__2497 (
            .O(N__10592),
            .I(N__10589));
    InMux I__2496 (
            .O(N__10589),
            .I(N__10585));
    InMux I__2495 (
            .O(N__10588),
            .I(N__10582));
    LocalMux I__2494 (
            .O(N__10585),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__2493 (
            .O(N__10582),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    InMux I__2492 (
            .O(N__10577),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__2491 (
            .O(N__10574),
            .I(N__10571));
    LocalMux I__2490 (
            .O(N__10571),
            .I(N__10567));
    InMux I__2489 (
            .O(N__10570),
            .I(N__10564));
    Odrv4 I__2488 (
            .O(N__10567),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__2487 (
            .O(N__10564),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__2486 (
            .O(N__10559),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__2485 (
            .O(N__10556),
            .I(N__10552));
    InMux I__2484 (
            .O(N__10555),
            .I(N__10549));
    LocalMux I__2483 (
            .O(N__10552),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__2482 (
            .O(N__10549),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    InMux I__2481 (
            .O(N__10544),
            .I(N__10541));
    LocalMux I__2480 (
            .O(N__10541),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__2479 (
            .O(N__10538),
            .I(bfn_17_7_0_));
    InMux I__2478 (
            .O(N__10535),
            .I(N__10531));
    InMux I__2477 (
            .O(N__10534),
            .I(N__10528));
    LocalMux I__2476 (
            .O(N__10531),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__2475 (
            .O(N__10528),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__2474 (
            .O(N__10523),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__2473 (
            .O(N__10520),
            .I(N__10516));
    InMux I__2472 (
            .O(N__10519),
            .I(N__10513));
    LocalMux I__2471 (
            .O(N__10516),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__2470 (
            .O(N__10513),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__2469 (
            .O(N__10508),
            .I(N__10505));
    LocalMux I__2468 (
            .O(N__10505),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__2467 (
            .O(N__10502),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    InMux I__2466 (
            .O(N__10499),
            .I(N__10495));
    InMux I__2465 (
            .O(N__10498),
            .I(N__10492));
    LocalMux I__2464 (
            .O(N__10495),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__2463 (
            .O(N__10492),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    InMux I__2462 (
            .O(N__10487),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__2461 (
            .O(N__10484),
            .I(N__10480));
    InMux I__2460 (
            .O(N__10483),
            .I(N__10477));
    LocalMux I__2459 (
            .O(N__10480),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__2458 (
            .O(N__10477),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__2457 (
            .O(N__10472),
            .I(N__10469));
    LocalMux I__2456 (
            .O(N__10469),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__2455 (
            .O(N__10466),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__2454 (
            .O(N__10463),
            .I(N__10458));
    InMux I__2453 (
            .O(N__10462),
            .I(N__10453));
    InMux I__2452 (
            .O(N__10461),
            .I(N__10453));
    LocalMux I__2451 (
            .O(N__10458),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__2450 (
            .O(N__10453),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__2449 (
            .O(N__10448),
            .I(N__10442));
    InMux I__2448 (
            .O(N__10447),
            .I(N__10442));
    LocalMux I__2447 (
            .O(N__10442),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    CascadeMux I__2446 (
            .O(N__10439),
            .I(N__10436));
    InMux I__2445 (
            .O(N__10436),
            .I(N__10427));
    InMux I__2444 (
            .O(N__10435),
            .I(N__10427));
    InMux I__2443 (
            .O(N__10434),
            .I(N__10427));
    LocalMux I__2442 (
            .O(N__10427),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    CascadeMux I__2441 (
            .O(N__10424),
            .I(N__10421));
    InMux I__2440 (
            .O(N__10421),
            .I(N__10414));
    InMux I__2439 (
            .O(N__10420),
            .I(N__10414));
    CascadeMux I__2438 (
            .O(N__10419),
            .I(N__10409));
    LocalMux I__2437 (
            .O(N__10414),
            .I(N__10399));
    InMux I__2436 (
            .O(N__10413),
            .I(N__10395));
    InMux I__2435 (
            .O(N__10412),
            .I(N__10390));
    InMux I__2434 (
            .O(N__10409),
            .I(N__10387));
    CascadeMux I__2433 (
            .O(N__10408),
            .I(N__10384));
    CascadeMux I__2432 (
            .O(N__10407),
            .I(N__10381));
    CascadeMux I__2431 (
            .O(N__10406),
            .I(N__10378));
    CascadeMux I__2430 (
            .O(N__10405),
            .I(N__10371));
    CascadeMux I__2429 (
            .O(N__10404),
            .I(N__10368));
    CascadeMux I__2428 (
            .O(N__10403),
            .I(N__10365));
    CascadeMux I__2427 (
            .O(N__10402),
            .I(N__10358));
    Span4Mux_h I__2426 (
            .O(N__10399),
            .I(N__10355));
    InMux I__2425 (
            .O(N__10398),
            .I(N__10352));
    LocalMux I__2424 (
            .O(N__10395),
            .I(N__10349));
    InMux I__2423 (
            .O(N__10394),
            .I(N__10346));
    InMux I__2422 (
            .O(N__10393),
            .I(N__10343));
    LocalMux I__2421 (
            .O(N__10390),
            .I(N__10340));
    LocalMux I__2420 (
            .O(N__10387),
            .I(N__10337));
    InMux I__2419 (
            .O(N__10384),
            .I(N__10334));
    InMux I__2418 (
            .O(N__10381),
            .I(N__10329));
    InMux I__2417 (
            .O(N__10378),
            .I(N__10329));
    InMux I__2416 (
            .O(N__10377),
            .I(N__10326));
    InMux I__2415 (
            .O(N__10376),
            .I(N__10323));
    InMux I__2414 (
            .O(N__10375),
            .I(N__10318));
    InMux I__2413 (
            .O(N__10374),
            .I(N__10318));
    InMux I__2412 (
            .O(N__10371),
            .I(N__10315));
    InMux I__2411 (
            .O(N__10368),
            .I(N__10306));
    InMux I__2410 (
            .O(N__10365),
            .I(N__10306));
    InMux I__2409 (
            .O(N__10364),
            .I(N__10306));
    InMux I__2408 (
            .O(N__10363),
            .I(N__10306));
    CascadeMux I__2407 (
            .O(N__10362),
            .I(N__10302));
    InMux I__2406 (
            .O(N__10361),
            .I(N__10297));
    InMux I__2405 (
            .O(N__10358),
            .I(N__10297));
    Span4Mux_h I__2404 (
            .O(N__10355),
            .I(N__10294));
    LocalMux I__2403 (
            .O(N__10352),
            .I(N__10291));
    Span4Mux_v I__2402 (
            .O(N__10349),
            .I(N__10287));
    LocalMux I__2401 (
            .O(N__10346),
            .I(N__10284));
    LocalMux I__2400 (
            .O(N__10343),
            .I(N__10281));
    Span4Mux_h I__2399 (
            .O(N__10340),
            .I(N__10272));
    Span4Mux_v I__2398 (
            .O(N__10337),
            .I(N__10272));
    LocalMux I__2397 (
            .O(N__10334),
            .I(N__10272));
    LocalMux I__2396 (
            .O(N__10329),
            .I(N__10272));
    LocalMux I__2395 (
            .O(N__10326),
            .I(N__10260));
    LocalMux I__2394 (
            .O(N__10323),
            .I(N__10260));
    LocalMux I__2393 (
            .O(N__10318),
            .I(N__10260));
    LocalMux I__2392 (
            .O(N__10315),
            .I(N__10260));
    LocalMux I__2391 (
            .O(N__10306),
            .I(N__10260));
    InMux I__2390 (
            .O(N__10305),
            .I(N__10255));
    InMux I__2389 (
            .O(N__10302),
            .I(N__10255));
    LocalMux I__2388 (
            .O(N__10297),
            .I(N__10252));
    Span4Mux_h I__2387 (
            .O(N__10294),
            .I(N__10247));
    Span4Mux_v I__2386 (
            .O(N__10291),
            .I(N__10247));
    InMux I__2385 (
            .O(N__10290),
            .I(N__10244));
    Span4Mux_v I__2384 (
            .O(N__10287),
            .I(N__10239));
    Span4Mux_v I__2383 (
            .O(N__10284),
            .I(N__10239));
    Span4Mux_h I__2382 (
            .O(N__10281),
            .I(N__10234));
    Span4Mux_v I__2381 (
            .O(N__10272),
            .I(N__10234));
    InMux I__2380 (
            .O(N__10271),
            .I(N__10231));
    Span4Mux_v I__2379 (
            .O(N__10260),
            .I(N__10228));
    LocalMux I__2378 (
            .O(N__10255),
            .I(N__10225));
    Span4Mux_v I__2377 (
            .O(N__10252),
            .I(N__10218));
    Span4Mux_v I__2376 (
            .O(N__10247),
            .I(N__10218));
    LocalMux I__2375 (
            .O(N__10244),
            .I(N__10218));
    Span4Mux_h I__2374 (
            .O(N__10239),
            .I(N__10215));
    Span4Mux_h I__2373 (
            .O(N__10234),
            .I(N__10212));
    LocalMux I__2372 (
            .O(N__10231),
            .I(N__10209));
    Span4Mux_h I__2371 (
            .O(N__10228),
            .I(N__10204));
    Span4Mux_v I__2370 (
            .O(N__10225),
            .I(N__10204));
    Span4Mux_h I__2369 (
            .O(N__10218),
            .I(N__10201));
    Sp12to4 I__2368 (
            .O(N__10215),
            .I(N__10196));
    Sp12to4 I__2367 (
            .O(N__10212),
            .I(N__10196));
    Span12Mux_v I__2366 (
            .O(N__10209),
            .I(N__10189));
    Sp12to4 I__2365 (
            .O(N__10204),
            .I(N__10189));
    Sp12to4 I__2364 (
            .O(N__10201),
            .I(N__10189));
    Span12Mux_h I__2363 (
            .O(N__10196),
            .I(N__10186));
    Span12Mux_v I__2362 (
            .O(N__10189),
            .I(N__10183));
    Span12Mux_v I__2361 (
            .O(N__10186),
            .I(N__10178));
    Span12Mux_h I__2360 (
            .O(N__10183),
            .I(N__10178));
    Odrv12 I__2359 (
            .O(N__10178),
            .I(RESETn_c));
    InMux I__2358 (
            .O(N__10175),
            .I(N__10172));
    LocalMux I__2357 (
            .O(N__10172),
            .I(N__10168));
    InMux I__2356 (
            .O(N__10171),
            .I(N__10165));
    Span4Mux_v I__2355 (
            .O(N__10168),
            .I(N__10161));
    LocalMux I__2354 (
            .O(N__10165),
            .I(N__10158));
    InMux I__2353 (
            .O(N__10164),
            .I(N__10155));
    Odrv4 I__2352 (
            .O(N__10161),
            .I(\U409_CIA.VMAZ0 ));
    Odrv4 I__2351 (
            .O(N__10158),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__2350 (
            .O(N__10155),
            .I(\U409_CIA.VMAZ0 ));
    InMux I__2349 (
            .O(N__10148),
            .I(N__10142));
    InMux I__2348 (
            .O(N__10147),
            .I(N__10135));
    InMux I__2347 (
            .O(N__10146),
            .I(N__10135));
    InMux I__2346 (
            .O(N__10145),
            .I(N__10135));
    LocalMux I__2345 (
            .O(N__10142),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__2344 (
            .O(N__10135),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    SRMux I__2343 (
            .O(N__10130),
            .I(N__10097));
    SRMux I__2342 (
            .O(N__10129),
            .I(N__10097));
    SRMux I__2341 (
            .O(N__10128),
            .I(N__10097));
    SRMux I__2340 (
            .O(N__10127),
            .I(N__10097));
    SRMux I__2339 (
            .O(N__10126),
            .I(N__10097));
    SRMux I__2338 (
            .O(N__10125),
            .I(N__10097));
    SRMux I__2337 (
            .O(N__10124),
            .I(N__10097));
    SRMux I__2336 (
            .O(N__10123),
            .I(N__10097));
    SRMux I__2335 (
            .O(N__10122),
            .I(N__10097));
    SRMux I__2334 (
            .O(N__10121),
            .I(N__10097));
    SRMux I__2333 (
            .O(N__10120),
            .I(N__10097));
    GlobalMux I__2332 (
            .O(N__10097),
            .I(N__10094));
    gio2CtrlBuf I__2331 (
            .O(N__10094),
            .I(RESETn_c_i_g));
    CascadeMux I__2330 (
            .O(N__10091),
            .I(N__10087));
    CascadeMux I__2329 (
            .O(N__10090),
            .I(N__10084));
    InMux I__2328 (
            .O(N__10087),
            .I(N__10078));
    InMux I__2327 (
            .O(N__10084),
            .I(N__10078));
    InMux I__2326 (
            .O(N__10083),
            .I(N__10075));
    LocalMux I__2325 (
            .O(N__10078),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__2324 (
            .O(N__10075),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    CascadeMux I__2323 (
            .O(N__10070),
            .I(N__10066));
    CascadeMux I__2322 (
            .O(N__10069),
            .I(N__10061));
    InMux I__2321 (
            .O(N__10066),
            .I(N__10058));
    InMux I__2320 (
            .O(N__10065),
            .I(N__10053));
    InMux I__2319 (
            .O(N__10064),
            .I(N__10053));
    InMux I__2318 (
            .O(N__10061),
            .I(N__10050));
    LocalMux I__2317 (
            .O(N__10058),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2316 (
            .O(N__10053),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__2315 (
            .O(N__10050),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__2314 (
            .O(N__10043),
            .I(N__10039));
    InMux I__2313 (
            .O(N__10042),
            .I(N__10036));
    LocalMux I__2312 (
            .O(N__10039),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__2311 (
            .O(N__10036),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    InMux I__2310 (
            .O(N__10031),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    InMux I__2309 (
            .O(N__10028),
            .I(N__10024));
    InMux I__2308 (
            .O(N__10027),
            .I(N__10021));
    LocalMux I__2307 (
            .O(N__10024),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__2306 (
            .O(N__10021),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    InMux I__2305 (
            .O(N__10016),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__2304 (
            .O(N__10013),
            .I(N__10009));
    InMux I__2303 (
            .O(N__10012),
            .I(N__10006));
    LocalMux I__2302 (
            .O(N__10009),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__2301 (
            .O(N__10006),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    InMux I__2300 (
            .O(N__10001),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__2299 (
            .O(N__9998),
            .I(N__9994));
    InMux I__2298 (
            .O(N__9997),
            .I(N__9991));
    LocalMux I__2297 (
            .O(N__9994),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__2296 (
            .O(N__9991),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    CascadeMux I__2295 (
            .O(N__9986),
            .I(N__9983));
    InMux I__2294 (
            .O(N__9983),
            .I(N__9980));
    LocalMux I__2293 (
            .O(N__9980),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__2292 (
            .O(N__9977),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    CascadeMux I__2291 (
            .O(N__9974),
            .I(N__9971));
    InMux I__2290 (
            .O(N__9971),
            .I(N__9968));
    LocalMux I__2289 (
            .O(N__9968),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__2288 (
            .O(N__9965),
            .I(N__9961));
    InMux I__2287 (
            .O(N__9964),
            .I(N__9958));
    LocalMux I__2286 (
            .O(N__9961),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__2285 (
            .O(N__9958),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    InMux I__2284 (
            .O(N__9953),
            .I(N__9950));
    LocalMux I__2283 (
            .O(N__9950),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__2282 (
            .O(N__9947),
            .I(N__9943));
    InMux I__2281 (
            .O(N__9946),
            .I(N__9940));
    LocalMux I__2280 (
            .O(N__9943),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__2279 (
            .O(N__9940),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    CascadeMux I__2278 (
            .O(N__9935),
            .I(N__9928));
    CascadeMux I__2277 (
            .O(N__9934),
            .I(N__9924));
    InMux I__2276 (
            .O(N__9933),
            .I(N__9921));
    InMux I__2275 (
            .O(N__9932),
            .I(N__9918));
    InMux I__2274 (
            .O(N__9931),
            .I(N__9915));
    InMux I__2273 (
            .O(N__9928),
            .I(N__9912));
    InMux I__2272 (
            .O(N__9927),
            .I(N__9909));
    InMux I__2271 (
            .O(N__9924),
            .I(N__9906));
    LocalMux I__2270 (
            .O(N__9921),
            .I(N__9900));
    LocalMux I__2269 (
            .O(N__9918),
            .I(N__9892));
    LocalMux I__2268 (
            .O(N__9915),
            .I(N__9886));
    LocalMux I__2267 (
            .O(N__9912),
            .I(N__9883));
    LocalMux I__2266 (
            .O(N__9909),
            .I(N__9880));
    LocalMux I__2265 (
            .O(N__9906),
            .I(N__9877));
    ClkMux I__2264 (
            .O(N__9905),
            .I(N__9842));
    ClkMux I__2263 (
            .O(N__9904),
            .I(N__9842));
    ClkMux I__2262 (
            .O(N__9903),
            .I(N__9842));
    Glb2LocalMux I__2261 (
            .O(N__9900),
            .I(N__9842));
    ClkMux I__2260 (
            .O(N__9899),
            .I(N__9842));
    ClkMux I__2259 (
            .O(N__9898),
            .I(N__9842));
    ClkMux I__2258 (
            .O(N__9897),
            .I(N__9842));
    ClkMux I__2257 (
            .O(N__9896),
            .I(N__9842));
    ClkMux I__2256 (
            .O(N__9895),
            .I(N__9842));
    Glb2LocalMux I__2255 (
            .O(N__9892),
            .I(N__9842));
    ClkMux I__2254 (
            .O(N__9891),
            .I(N__9842));
    ClkMux I__2253 (
            .O(N__9890),
            .I(N__9842));
    ClkMux I__2252 (
            .O(N__9889),
            .I(N__9842));
    Glb2LocalMux I__2251 (
            .O(N__9886),
            .I(N__9842));
    Glb2LocalMux I__2250 (
            .O(N__9883),
            .I(N__9842));
    Glb2LocalMux I__2249 (
            .O(N__9880),
            .I(N__9842));
    Glb2LocalMux I__2248 (
            .O(N__9877),
            .I(N__9842));
    GlobalMux I__2247 (
            .O(N__9842),
            .I(N__9839));
    gio2CtrlBuf I__2246 (
            .O(N__9839),
            .I(CLK40_IN_c_g));
    InMux I__2245 (
            .O(N__9836),
            .I(N__9833));
    LocalMux I__2244 (
            .O(N__9833),
            .I(\U409_TRANSFER_ACK.N_17_mux ));
    CascadeMux I__2243 (
            .O(N__9830),
            .I(\U409_TRANSFER_ACK.N_17_mux_cascade_ ));
    InMux I__2242 (
            .O(N__9827),
            .I(N__9824));
    LocalMux I__2241 (
            .O(N__9824),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0 ));
    CascadeMux I__2240 (
            .O(N__9821),
            .I(\U409_TRANSFER_ACK.N_3_0_cascade_ ));
    InMux I__2239 (
            .O(N__9818),
            .I(N__9815));
    LocalMux I__2238 (
            .O(N__9815),
            .I(\U409_TRANSFER_ACK.N_6_0 ));
    InMux I__2237 (
            .O(N__9812),
            .I(N__9809));
    LocalMux I__2236 (
            .O(N__9809),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__2235 (
            .O(N__9806),
            .I(N__9802));
    InMux I__2234 (
            .O(N__9805),
            .I(N__9799));
    LocalMux I__2233 (
            .O(N__9802),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__2232 (
            .O(N__9799),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__2231 (
            .O(N__9794),
            .I(N__9781));
    InMux I__2230 (
            .O(N__9793),
            .I(N__9781));
    InMux I__2229 (
            .O(N__9792),
            .I(N__9781));
    InMux I__2228 (
            .O(N__9791),
            .I(N__9772));
    InMux I__2227 (
            .O(N__9790),
            .I(N__9772));
    InMux I__2226 (
            .O(N__9789),
            .I(N__9772));
    InMux I__2225 (
            .O(N__9788),
            .I(N__9772));
    LocalMux I__2224 (
            .O(N__9781),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__2223 (
            .O(N__9772),
            .I(\U409_TICK.TICK603_14 ));
    CascadeMux I__2222 (
            .O(N__9767),
            .I(N__9760));
    CascadeMux I__2221 (
            .O(N__9766),
            .I(N__9757));
    CascadeMux I__2220 (
            .O(N__9765),
            .I(N__9754));
    CascadeMux I__2219 (
            .O(N__9764),
            .I(N__9750));
    InMux I__2218 (
            .O(N__9763),
            .I(N__9737));
    InMux I__2217 (
            .O(N__9760),
            .I(N__9737));
    InMux I__2216 (
            .O(N__9757),
            .I(N__9737));
    InMux I__2215 (
            .O(N__9754),
            .I(N__9737));
    InMux I__2214 (
            .O(N__9753),
            .I(N__9737));
    InMux I__2213 (
            .O(N__9750),
            .I(N__9730));
    InMux I__2212 (
            .O(N__9749),
            .I(N__9730));
    InMux I__2211 (
            .O(N__9748),
            .I(N__9730));
    LocalMux I__2210 (
            .O(N__9737),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__2209 (
            .O(N__9730),
            .I(\U409_TICK.TICK603_9 ));
    CascadeMux I__2208 (
            .O(N__9725),
            .I(N__9721));
    CascadeMux I__2207 (
            .O(N__9724),
            .I(N__9717));
    InMux I__2206 (
            .O(N__9721),
            .I(N__9705));
    InMux I__2205 (
            .O(N__9720),
            .I(N__9705));
    InMux I__2204 (
            .O(N__9717),
            .I(N__9705));
    InMux I__2203 (
            .O(N__9716),
            .I(N__9694));
    InMux I__2202 (
            .O(N__9715),
            .I(N__9694));
    InMux I__2201 (
            .O(N__9714),
            .I(N__9694));
    InMux I__2200 (
            .O(N__9713),
            .I(N__9694));
    InMux I__2199 (
            .O(N__9712),
            .I(N__9694));
    LocalMux I__2198 (
            .O(N__9705),
            .I(N__9691));
    LocalMux I__2197 (
            .O(N__9694),
            .I(\U409_TICK.TICK603_10 ));
    Odrv4 I__2196 (
            .O(N__9691),
            .I(\U409_TICK.TICK603_10 ));
    InMux I__2195 (
            .O(N__9686),
            .I(N__9683));
    LocalMux I__2194 (
            .O(N__9683),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__2193 (
            .O(N__9680),
            .I(N__9676));
    InMux I__2192 (
            .O(N__9679),
            .I(N__9673));
    LocalMux I__2191 (
            .O(N__9676),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__2190 (
            .O(N__9673),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    CascadeMux I__2189 (
            .O(N__9668),
            .I(N__9665));
    InMux I__2188 (
            .O(N__9665),
            .I(N__9662));
    LocalMux I__2187 (
            .O(N__9662),
            .I(N__9655));
    InMux I__2186 (
            .O(N__9661),
            .I(N__9652));
    InMux I__2185 (
            .O(N__9660),
            .I(N__9645));
    InMux I__2184 (
            .O(N__9659),
            .I(N__9645));
    InMux I__2183 (
            .O(N__9658),
            .I(N__9645));
    Odrv4 I__2182 (
            .O(N__9655),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__2181 (
            .O(N__9652),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__2180 (
            .O(N__9645),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    InMux I__2179 (
            .O(N__9638),
            .I(N__9635));
    LocalMux I__2178 (
            .O(N__9635),
            .I(\U409_TRANSFER_ACK.N_3_0 ));
    InMux I__2177 (
            .O(N__9632),
            .I(N__9629));
    LocalMux I__2176 (
            .O(N__9629),
            .I(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ));
    CascadeMux I__2175 (
            .O(N__9626),
            .I(N__9620));
    InMux I__2174 (
            .O(N__9625),
            .I(N__9607));
    InMux I__2173 (
            .O(N__9624),
            .I(N__9607));
    InMux I__2172 (
            .O(N__9623),
            .I(N__9607));
    InMux I__2171 (
            .O(N__9620),
            .I(N__9607));
    InMux I__2170 (
            .O(N__9619),
            .I(N__9598));
    InMux I__2169 (
            .O(N__9618),
            .I(N__9598));
    InMux I__2168 (
            .O(N__9617),
            .I(N__9598));
    InMux I__2167 (
            .O(N__9616),
            .I(N__9598));
    LocalMux I__2166 (
            .O(N__9607),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__2165 (
            .O(N__9598),
            .I(\U409_TICK.TICK503_10 ));
    InMux I__2164 (
            .O(N__9593),
            .I(N__9574));
    InMux I__2163 (
            .O(N__9592),
            .I(N__9574));
    InMux I__2162 (
            .O(N__9591),
            .I(N__9574));
    InMux I__2161 (
            .O(N__9590),
            .I(N__9574));
    InMux I__2160 (
            .O(N__9589),
            .I(N__9574));
    InMux I__2159 (
            .O(N__9588),
            .I(N__9565));
    InMux I__2158 (
            .O(N__9587),
            .I(N__9565));
    InMux I__2157 (
            .O(N__9586),
            .I(N__9565));
    InMux I__2156 (
            .O(N__9585),
            .I(N__9565));
    LocalMux I__2155 (
            .O(N__9574),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__2154 (
            .O(N__9565),
            .I(\U409_TICK.TICK503_14 ));
    CascadeMux I__2153 (
            .O(N__9560),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    IoInMux I__2152 (
            .O(N__9557),
            .I(N__9554));
    LocalMux I__2151 (
            .O(N__9554),
            .I(N__9551));
    Span4Mux_s1_v I__2150 (
            .O(N__9551),
            .I(N__9548));
    Sp12to4 I__2149 (
            .O(N__9548),
            .I(N__9545));
    Span12Mux_h I__2148 (
            .O(N__9545),
            .I(N__9541));
    InMux I__2147 (
            .O(N__9544),
            .I(N__9538));
    Odrv12 I__2146 (
            .O(N__9541),
            .I(TICK60_c));
    LocalMux I__2145 (
            .O(N__9538),
            .I(TICK60_c));
    InMux I__2144 (
            .O(N__9533),
            .I(N__9529));
    InMux I__2143 (
            .O(N__9532),
            .I(N__9526));
    LocalMux I__2142 (
            .O(N__9529),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__2141 (
            .O(N__9526),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__2140 (
            .O(N__9521),
            .I(N__9518));
    LocalMux I__2139 (
            .O(N__9518),
            .I(N__9514));
    InMux I__2138 (
            .O(N__9517),
            .I(N__9511));
    Odrv4 I__2137 (
            .O(N__9514),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__2136 (
            .O(N__9511),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    CascadeMux I__2135 (
            .O(N__9506),
            .I(\U409_TICK.TICK603_8_cascade_ ));
    InMux I__2134 (
            .O(N__9503),
            .I(N__9499));
    InMux I__2133 (
            .O(N__9502),
            .I(N__9496));
    LocalMux I__2132 (
            .O(N__9499),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__2131 (
            .O(N__9496),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    CascadeMux I__2130 (
            .O(N__9491),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    InMux I__2129 (
            .O(N__9488),
            .I(N__9484));
    CascadeMux I__2128 (
            .O(N__9487),
            .I(N__9479));
    LocalMux I__2127 (
            .O(N__9484),
            .I(N__9476));
    InMux I__2126 (
            .O(N__9483),
            .I(N__9473));
    InMux I__2125 (
            .O(N__9482),
            .I(N__9470));
    InMux I__2124 (
            .O(N__9479),
            .I(N__9467));
    Odrv4 I__2123 (
            .O(N__9476),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2122 (
            .O(N__9473),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2121 (
            .O(N__9470),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__2120 (
            .O(N__9467),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__2119 (
            .O(N__9458),
            .I(N__9455));
    LocalMux I__2118 (
            .O(N__9455),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    CascadeMux I__2117 (
            .O(N__9452),
            .I(N__9449));
    InMux I__2116 (
            .O(N__9449),
            .I(N__9446));
    LocalMux I__2115 (
            .O(N__9446),
            .I(N__9442));
    InMux I__2114 (
            .O(N__9445),
            .I(N__9439));
    Odrv4 I__2113 (
            .O(N__9442),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__2112 (
            .O(N__9439),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    InMux I__2111 (
            .O(N__9434),
            .I(N__9430));
    InMux I__2110 (
            .O(N__9433),
            .I(N__9427));
    LocalMux I__2109 (
            .O(N__9430),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__2108 (
            .O(N__9427),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__2107 (
            .O(N__9422),
            .I(N__9418));
    InMux I__2106 (
            .O(N__9421),
            .I(N__9415));
    LocalMux I__2105 (
            .O(N__9418),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__2104 (
            .O(N__9415),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    CascadeMux I__2103 (
            .O(N__9410),
            .I(N__9406));
    InMux I__2102 (
            .O(N__9409),
            .I(N__9402));
    InMux I__2101 (
            .O(N__9406),
            .I(N__9399));
    InMux I__2100 (
            .O(N__9405),
            .I(N__9396));
    LocalMux I__2099 (
            .O(N__9402),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__2098 (
            .O(N__9399),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__2097 (
            .O(N__9396),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    InMux I__2096 (
            .O(N__9389),
            .I(N__9385));
    InMux I__2095 (
            .O(N__9388),
            .I(N__9382));
    LocalMux I__2094 (
            .O(N__9385),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__2093 (
            .O(N__9382),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    InMux I__2092 (
            .O(N__9377),
            .I(N__9374));
    LocalMux I__2091 (
            .O(N__9374),
            .I(\U409_TICK.TICK603_11 ));
    InMux I__2090 (
            .O(N__9371),
            .I(N__9368));
    LocalMux I__2089 (
            .O(N__9368),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__2088 (
            .O(N__9365),
            .I(N__9361));
    InMux I__2087 (
            .O(N__9364),
            .I(N__9358));
    LocalMux I__2086 (
            .O(N__9361),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__2085 (
            .O(N__9358),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    InMux I__2084 (
            .O(N__9353),
            .I(N__9350));
    LocalMux I__2083 (
            .O(N__9350),
            .I(\U409_TICK.TICK503_11 ));
    CascadeMux I__2082 (
            .O(N__9347),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    CascadeMux I__2081 (
            .O(N__9344),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    CascadeMux I__2080 (
            .O(N__9341),
            .I(N__9332));
    CascadeMux I__2079 (
            .O(N__9340),
            .I(N__9329));
    InMux I__2078 (
            .O(N__9339),
            .I(N__9319));
    InMux I__2077 (
            .O(N__9338),
            .I(N__9319));
    InMux I__2076 (
            .O(N__9337),
            .I(N__9319));
    InMux I__2075 (
            .O(N__9336),
            .I(N__9319));
    InMux I__2074 (
            .O(N__9335),
            .I(N__9310));
    InMux I__2073 (
            .O(N__9332),
            .I(N__9310));
    InMux I__2072 (
            .O(N__9329),
            .I(N__9310));
    InMux I__2071 (
            .O(N__9328),
            .I(N__9310));
    LocalMux I__2070 (
            .O(N__9319),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__2069 (
            .O(N__9310),
            .I(\U409_TICK.TICK503_9 ));
    InMux I__2068 (
            .O(N__9305),
            .I(N__9299));
    InMux I__2067 (
            .O(N__9304),
            .I(N__9290));
    InMux I__2066 (
            .O(N__9303),
            .I(N__9290));
    InMux I__2065 (
            .O(N__9302),
            .I(N__9290));
    LocalMux I__2064 (
            .O(N__9299),
            .I(N__9287));
    InMux I__2063 (
            .O(N__9298),
            .I(N__9282));
    InMux I__2062 (
            .O(N__9297),
            .I(N__9282));
    LocalMux I__2061 (
            .O(N__9290),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    Odrv4 I__2060 (
            .O(N__9287),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__2059 (
            .O(N__9282),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    CascadeMux I__2058 (
            .O(N__9275),
            .I(N__9269));
    InMux I__2057 (
            .O(N__9274),
            .I(N__9263));
    InMux I__2056 (
            .O(N__9273),
            .I(N__9256));
    InMux I__2055 (
            .O(N__9272),
            .I(N__9256));
    InMux I__2054 (
            .O(N__9269),
            .I(N__9256));
    InMux I__2053 (
            .O(N__9268),
            .I(N__9253));
    InMux I__2052 (
            .O(N__9267),
            .I(N__9248));
    InMux I__2051 (
            .O(N__9266),
            .I(N__9248));
    LocalMux I__2050 (
            .O(N__9263),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__2049 (
            .O(N__9256),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__2048 (
            .O(N__9253),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__2047 (
            .O(N__9248),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    InMux I__2046 (
            .O(N__9239),
            .I(N__9227));
    InMux I__2045 (
            .O(N__9238),
            .I(N__9227));
    InMux I__2044 (
            .O(N__9237),
            .I(N__9227));
    InMux I__2043 (
            .O(N__9236),
            .I(N__9220));
    InMux I__2042 (
            .O(N__9235),
            .I(N__9220));
    InMux I__2041 (
            .O(N__9234),
            .I(N__9220));
    LocalMux I__2040 (
            .O(N__9227),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__2039 (
            .O(N__9220),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__2038 (
            .O(N__9215),
            .I(N__9209));
    CascadeMux I__2037 (
            .O(N__9214),
            .I(N__9206));
    InMux I__2036 (
            .O(N__9213),
            .I(N__9202));
    CascadeMux I__2035 (
            .O(N__9212),
            .I(N__9199));
    InMux I__2034 (
            .O(N__9209),
            .I(N__9191));
    InMux I__2033 (
            .O(N__9206),
            .I(N__9191));
    InMux I__2032 (
            .O(N__9205),
            .I(N__9191));
    LocalMux I__2031 (
            .O(N__9202),
            .I(N__9188));
    InMux I__2030 (
            .O(N__9199),
            .I(N__9183));
    InMux I__2029 (
            .O(N__9198),
            .I(N__9183));
    LocalMux I__2028 (
            .O(N__9191),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    Odrv4 I__2027 (
            .O(N__9188),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__2026 (
            .O(N__9183),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    InMux I__2025 (
            .O(N__9176),
            .I(N__9172));
    CascadeMux I__2024 (
            .O(N__9175),
            .I(N__9168));
    LocalMux I__2023 (
            .O(N__9172),
            .I(N__9165));
    InMux I__2022 (
            .O(N__9171),
            .I(N__9162));
    InMux I__2021 (
            .O(N__9168),
            .I(N__9159));
    Span4Mux_v I__2020 (
            .O(N__9165),
            .I(N__9154));
    LocalMux I__2019 (
            .O(N__9162),
            .I(N__9154));
    LocalMux I__2018 (
            .O(N__9159),
            .I(N__9151));
    Span4Mux_v I__2017 (
            .O(N__9154),
            .I(N__9148));
    Span4Mux_v I__2016 (
            .O(N__9151),
            .I(N__9143));
    Span4Mux_h I__2015 (
            .O(N__9148),
            .I(N__9143));
    Sp12to4 I__2014 (
            .O(N__9143),
            .I(N__9140));
    Odrv12 I__2013 (
            .O(N__9140),
            .I(ROMEN));
    IoInMux I__2012 (
            .O(N__9137),
            .I(N__9134));
    LocalMux I__2011 (
            .O(N__9134),
            .I(N__9130));
    IoInMux I__2010 (
            .O(N__9133),
            .I(N__9127));
    IoSpan4Mux I__2009 (
            .O(N__9130),
            .I(N__9122));
    LocalMux I__2008 (
            .O(N__9127),
            .I(N__9122));
    IoSpan4Mux I__2007 (
            .O(N__9122),
            .I(N__9119));
    IoSpan4Mux I__2006 (
            .O(N__9119),
            .I(N__9116));
    Span4Mux_s0_v I__2005 (
            .O(N__9116),
            .I(N__9113));
    Span4Mux_v I__2004 (
            .O(N__9113),
            .I(N__9109));
    InMux I__2003 (
            .O(N__9112),
            .I(N__9106));
    Span4Mux_v I__2002 (
            .O(N__9109),
            .I(N__9101));
    LocalMux I__2001 (
            .O(N__9106),
            .I(N__9101));
    Span4Mux_v I__2000 (
            .O(N__9101),
            .I(N__9097));
    CascadeMux I__1999 (
            .O(N__9100),
            .I(N__9094));
    Span4Mux_v I__1998 (
            .O(N__9097),
            .I(N__9091));
    InMux I__1997 (
            .O(N__9094),
            .I(N__9088));
    Odrv4 I__1996 (
            .O(N__9091),
            .I(TACK_EN));
    LocalMux I__1995 (
            .O(N__9088),
            .I(TACK_EN));
    IoInMux I__1994 (
            .O(N__9083),
            .I(N__9080));
    LocalMux I__1993 (
            .O(N__9080),
            .I(N__9077));
    Span4Mux_s2_v I__1992 (
            .O(N__9077),
            .I(N__9074));
    Span4Mux_v I__1991 (
            .O(N__9074),
            .I(N__9071));
    Span4Mux_v I__1990 (
            .O(N__9071),
            .I(N__9068));
    Sp12to4 I__1989 (
            .O(N__9068),
            .I(N__9065));
    Odrv12 I__1988 (
            .O(N__9065),
            .I(TCIn_1_i));
    IoInMux I__1987 (
            .O(N__9062),
            .I(N__9059));
    LocalMux I__1986 (
            .O(N__9059),
            .I(N__9056));
    Span4Mux_s3_v I__1985 (
            .O(N__9056),
            .I(N__9053));
    Span4Mux_v I__1984 (
            .O(N__9053),
            .I(N__9050));
    Span4Mux_h I__1983 (
            .O(N__9050),
            .I(N__9047));
    Span4Mux_h I__1982 (
            .O(N__9047),
            .I(N__9043));
    InMux I__1981 (
            .O(N__9046),
            .I(N__9040));
    Odrv4 I__1980 (
            .O(N__9043),
            .I(TICK50_c));
    LocalMux I__1979 (
            .O(N__9040),
            .I(TICK50_c));
    InMux I__1978 (
            .O(N__9035),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__1977 (
            .O(N__9032),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__1976 (
            .O(N__9029),
            .I(N__9025));
    InMux I__1975 (
            .O(N__9028),
            .I(N__9022));
    LocalMux I__1974 (
            .O(N__9025),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__1973 (
            .O(N__9022),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__1972 (
            .O(N__9017),
            .I(N__9013));
    InMux I__1971 (
            .O(N__9016),
            .I(N__9010));
    LocalMux I__1970 (
            .O(N__9013),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__1969 (
            .O(N__9010),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    CascadeMux I__1968 (
            .O(N__9005),
            .I(N__9002));
    InMux I__1967 (
            .O(N__9002),
            .I(N__8999));
    LocalMux I__1966 (
            .O(N__8999),
            .I(N__8995));
    InMux I__1965 (
            .O(N__8998),
            .I(N__8992));
    Odrv4 I__1964 (
            .O(N__8995),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__1963 (
            .O(N__8992),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    CascadeMux I__1962 (
            .O(N__8987),
            .I(N__8982));
    InMux I__1961 (
            .O(N__8986),
            .I(N__8979));
    InMux I__1960 (
            .O(N__8985),
            .I(N__8976));
    InMux I__1959 (
            .O(N__8982),
            .I(N__8973));
    LocalMux I__1958 (
            .O(N__8979),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1957 (
            .O(N__8976),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__1956 (
            .O(N__8973),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    InMux I__1955 (
            .O(N__8966),
            .I(N__8962));
    InMux I__1954 (
            .O(N__8965),
            .I(N__8959));
    LocalMux I__1953 (
            .O(N__8962),
            .I(N__8956));
    LocalMux I__1952 (
            .O(N__8959),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    Odrv12 I__1951 (
            .O(N__8956),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    InMux I__1950 (
            .O(N__8951),
            .I(N__8948));
    LocalMux I__1949 (
            .O(N__8948),
            .I(N__8944));
    InMux I__1948 (
            .O(N__8947),
            .I(N__8941));
    Span4Mux_v I__1947 (
            .O(N__8944),
            .I(N__8937));
    LocalMux I__1946 (
            .O(N__8941),
            .I(N__8934));
    InMux I__1945 (
            .O(N__8940),
            .I(N__8931));
    Odrv4 I__1944 (
            .O(N__8937),
            .I(\U409_TRANSFER_ACK.N_101 ));
    Odrv4 I__1943 (
            .O(N__8934),
            .I(\U409_TRANSFER_ACK.N_101 ));
    LocalMux I__1942 (
            .O(N__8931),
            .I(\U409_TRANSFER_ACK.N_101 ));
    InMux I__1941 (
            .O(N__8924),
            .I(N__8921));
    LocalMux I__1940 (
            .O(N__8921),
            .I(\U409_TRANSFER_ACK.N_19 ));
    IoInMux I__1939 (
            .O(N__8918),
            .I(N__8915));
    LocalMux I__1938 (
            .O(N__8915),
            .I(N__8912));
    Span4Mux_s0_v I__1937 (
            .O(N__8912),
            .I(N__8909));
    Span4Mux_v I__1936 (
            .O(N__8909),
            .I(N__8906));
    Span4Mux_v I__1935 (
            .O(N__8906),
            .I(N__8903));
    Span4Mux_v I__1934 (
            .O(N__8903),
            .I(N__8899));
    InMux I__1933 (
            .O(N__8902),
            .I(N__8896));
    Span4Mux_v I__1932 (
            .O(N__8899),
            .I(N__8890));
    LocalMux I__1931 (
            .O(N__8896),
            .I(N__8890));
    InMux I__1930 (
            .O(N__8895),
            .I(N__8887));
    Odrv4 I__1929 (
            .O(N__8890),
            .I(CLK_CIA_c));
    LocalMux I__1928 (
            .O(N__8887),
            .I(CLK_CIA_c));
    InMux I__1927 (
            .O(N__8882),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    InMux I__1926 (
            .O(N__8879),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    InMux I__1925 (
            .O(N__8876),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__1924 (
            .O(N__8873),
            .I(bfn_15_8_0_));
    InMux I__1923 (
            .O(N__8870),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__1922 (
            .O(N__8867),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__1921 (
            .O(N__8864),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__1920 (
            .O(N__8861),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__1919 (
            .O(N__8858),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    CascadeMux I__1918 (
            .O(N__8855),
            .I(\U409_TRANSFER_ACK.N_19_cascade_ ));
    InMux I__1917 (
            .O(N__8852),
            .I(N__8849));
    LocalMux I__1916 (
            .O(N__8849),
            .I(\U409_TRANSFER_ACK.N_23 ));
    InMux I__1915 (
            .O(N__8846),
            .I(N__8843));
    LocalMux I__1914 (
            .O(N__8843),
            .I(\U409_TRANSFER_ACK.N_22 ));
    IoInMux I__1913 (
            .O(N__8840),
            .I(N__8837));
    LocalMux I__1912 (
            .O(N__8837),
            .I(N__8834));
    Span4Mux_s3_v I__1911 (
            .O(N__8834),
            .I(N__8831));
    Sp12to4 I__1910 (
            .O(N__8831),
            .I(N__8828));
    Span12Mux_h I__1909 (
            .O(N__8828),
            .I(N__8824));
    InMux I__1908 (
            .O(N__8827),
            .I(N__8821));
    Odrv12 I__1907 (
            .O(N__8824),
            .I(ROMENn_c));
    LocalMux I__1906 (
            .O(N__8821),
            .I(ROMENn_c));
    InMux I__1905 (
            .O(N__8816),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__1904 (
            .O(N__8813),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__1903 (
            .O(N__8810),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__1902 (
            .O(N__8807),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    InMux I__1901 (
            .O(N__8804),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    InMux I__1900 (
            .O(N__8801),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ));
    InMux I__1899 (
            .O(N__8798),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ));
    InMux I__1898 (
            .O(N__8795),
            .I(N__8787));
    InMux I__1897 (
            .O(N__8794),
            .I(N__8784));
    InMux I__1896 (
            .O(N__8793),
            .I(N__8781));
    InMux I__1895 (
            .O(N__8792),
            .I(N__8778));
    InMux I__1894 (
            .O(N__8791),
            .I(N__8773));
    InMux I__1893 (
            .O(N__8790),
            .I(N__8773));
    LocalMux I__1892 (
            .O(N__8787),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1891 (
            .O(N__8784),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1890 (
            .O(N__8781),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1889 (
            .O(N__8778),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__1888 (
            .O(N__8773),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    CascadeMux I__1887 (
            .O(N__8762),
            .I(N__8757));
    InMux I__1886 (
            .O(N__8761),
            .I(N__8753));
    InMux I__1885 (
            .O(N__8760),
            .I(N__8750));
    InMux I__1884 (
            .O(N__8757),
            .I(N__8747));
    InMux I__1883 (
            .O(N__8756),
            .I(N__8744));
    LocalMux I__1882 (
            .O(N__8753),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__1881 (
            .O(N__8750),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__1880 (
            .O(N__8747),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__1879 (
            .O(N__8744),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    CascadeMux I__1878 (
            .O(N__8735),
            .I(N__8730));
    CascadeMux I__1877 (
            .O(N__8734),
            .I(N__8726));
    InMux I__1876 (
            .O(N__8733),
            .I(N__8723));
    InMux I__1875 (
            .O(N__8730),
            .I(N__8720));
    InMux I__1874 (
            .O(N__8729),
            .I(N__8717));
    InMux I__1873 (
            .O(N__8726),
            .I(N__8714));
    LocalMux I__1872 (
            .O(N__8723),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__1871 (
            .O(N__8720),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__1870 (
            .O(N__8717),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__1869 (
            .O(N__8714),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    CascadeMux I__1868 (
            .O(N__8705),
            .I(N__8697));
    InMux I__1867 (
            .O(N__8704),
            .I(N__8692));
    InMux I__1866 (
            .O(N__8703),
            .I(N__8692));
    InMux I__1865 (
            .O(N__8702),
            .I(N__8687));
    InMux I__1864 (
            .O(N__8701),
            .I(N__8687));
    InMux I__1863 (
            .O(N__8700),
            .I(N__8682));
    InMux I__1862 (
            .O(N__8697),
            .I(N__8682));
    LocalMux I__1861 (
            .O(N__8692),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1860 (
            .O(N__8687),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__1859 (
            .O(N__8682),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    InMux I__1858 (
            .O(N__8675),
            .I(N__8668));
    InMux I__1857 (
            .O(N__8674),
            .I(N__8663));
    InMux I__1856 (
            .O(N__8673),
            .I(N__8663));
    InMux I__1855 (
            .O(N__8672),
            .I(N__8660));
    InMux I__1854 (
            .O(N__8671),
            .I(N__8657));
    LocalMux I__1853 (
            .O(N__8668),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1852 (
            .O(N__8663),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1851 (
            .O(N__8660),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__1850 (
            .O(N__8657),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__1849 (
            .O(N__8648),
            .I(N__8645));
    LocalMux I__1848 (
            .O(N__8645),
            .I(\U409_CIA.CLK_CIA6_0 ));
    CascadeMux I__1847 (
            .O(N__8642),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_3_1_cascade_ ));
    InMux I__1846 (
            .O(N__8639),
            .I(N__8629));
    InMux I__1845 (
            .O(N__8638),
            .I(N__8629));
    InMux I__1844 (
            .O(N__8637),
            .I(N__8626));
    InMux I__1843 (
            .O(N__8636),
            .I(N__8623));
    InMux I__1842 (
            .O(N__8635),
            .I(N__8618));
    InMux I__1841 (
            .O(N__8634),
            .I(N__8618));
    LocalMux I__1840 (
            .O(N__8629),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1839 (
            .O(N__8626),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1838 (
            .O(N__8623),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__1837 (
            .O(N__8618),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    InMux I__1836 (
            .O(N__8609),
            .I(N__8606));
    LocalMux I__1835 (
            .O(N__8606),
            .I(N__8602));
    InMux I__1834 (
            .O(N__8605),
            .I(N__8599));
    Odrv12 I__1833 (
            .O(N__8602),
            .I(CIA_SPACE));
    LocalMux I__1832 (
            .O(N__8599),
            .I(CIA_SPACE));
    CascadeMux I__1831 (
            .O(N__8594),
            .I(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ));
    CascadeMux I__1830 (
            .O(N__8591),
            .I(N__8588));
    InMux I__1829 (
            .O(N__8588),
            .I(N__8585));
    LocalMux I__1828 (
            .O(N__8585),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_5_0_0 ));
    InMux I__1827 (
            .O(N__8582),
            .I(N__8579));
    LocalMux I__1826 (
            .O(N__8579),
            .I(N__8573));
    InMux I__1825 (
            .O(N__8578),
            .I(N__8570));
    InMux I__1824 (
            .O(N__8577),
            .I(N__8566));
    InMux I__1823 (
            .O(N__8576),
            .I(N__8563));
    Span4Mux_h I__1822 (
            .O(N__8573),
            .I(N__8558));
    LocalMux I__1821 (
            .O(N__8570),
            .I(N__8558));
    InMux I__1820 (
            .O(N__8569),
            .I(N__8555));
    LocalMux I__1819 (
            .O(N__8566),
            .I(N__8550));
    LocalMux I__1818 (
            .O(N__8563),
            .I(N__8550));
    Span4Mux_h I__1817 (
            .O(N__8558),
            .I(N__8545));
    LocalMux I__1816 (
            .O(N__8555),
            .I(N__8545));
    Span4Mux_v I__1815 (
            .O(N__8550),
            .I(N__8542));
    Span4Mux_v I__1814 (
            .O(N__8545),
            .I(N__8539));
    Sp12to4 I__1813 (
            .O(N__8542),
            .I(N__8534));
    Sp12to4 I__1812 (
            .O(N__8539),
            .I(N__8534));
    Span12Mux_h I__1811 (
            .O(N__8534),
            .I(N__8531));
    Span12Mux_v I__1810 (
            .O(N__8531),
            .I(N__8528));
    Odrv12 I__1809 (
            .O(N__8528),
            .I(TSn_c));
    CascadeMux I__1808 (
            .O(N__8525),
            .I(CIA_ENABLE_cascade_));
    CascadeMux I__1807 (
            .O(N__8522),
            .I(N__8519));
    InMux I__1806 (
            .O(N__8519),
            .I(N__8512));
    InMux I__1805 (
            .O(N__8518),
            .I(N__8512));
    InMux I__1804 (
            .O(N__8517),
            .I(N__8509));
    LocalMux I__1803 (
            .O(N__8512),
            .I(N__8506));
    LocalMux I__1802 (
            .O(N__8509),
            .I(N__8503));
    Span4Mux_v I__1801 (
            .O(N__8506),
            .I(N__8500));
    Span12Mux_h I__1800 (
            .O(N__8503),
            .I(N__8495));
    Sp12to4 I__1799 (
            .O(N__8500),
            .I(N__8495));
    Odrv12 I__1798 (
            .O(N__8495),
            .I(A_c_12));
    IoInMux I__1797 (
            .O(N__8492),
            .I(N__8489));
    LocalMux I__1796 (
            .O(N__8489),
            .I(N__8486));
    IoSpan4Mux I__1795 (
            .O(N__8486),
            .I(N__8483));
    Span4Mux_s3_h I__1794 (
            .O(N__8483),
            .I(N__8480));
    Sp12to4 I__1793 (
            .O(N__8480),
            .I(N__8477));
    Span12Mux_h I__1792 (
            .O(N__8477),
            .I(N__8474));
    Odrv12 I__1791 (
            .O(N__8474),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    InMux I__1790 (
            .O(N__8471),
            .I(N__8468));
    LocalMux I__1789 (
            .O(N__8468),
            .I(CIA_ENABLE));
    InMux I__1788 (
            .O(N__8465),
            .I(N__8462));
    LocalMux I__1787 (
            .O(N__8462),
            .I(N__8457));
    InMux I__1786 (
            .O(N__8461),
            .I(N__8452));
    InMux I__1785 (
            .O(N__8460),
            .I(N__8452));
    Span12Mux_v I__1784 (
            .O(N__8457),
            .I(N__8449));
    LocalMux I__1783 (
            .O(N__8452),
            .I(N__8446));
    Span12Mux_h I__1782 (
            .O(N__8449),
            .I(N__8443));
    Span12Mux_v I__1781 (
            .O(N__8446),
            .I(N__8440));
    Odrv12 I__1780 (
            .O(N__8443),
            .I(A_c_13));
    Odrv12 I__1779 (
            .O(N__8440),
            .I(A_c_13));
    IoInMux I__1778 (
            .O(N__8435),
            .I(N__8432));
    LocalMux I__1777 (
            .O(N__8432),
            .I(N__8429));
    Span4Mux_s2_h I__1776 (
            .O(N__8429),
            .I(N__8426));
    Sp12to4 I__1775 (
            .O(N__8426),
            .I(N__8423));
    Span12Mux_s10_v I__1774 (
            .O(N__8423),
            .I(N__8420));
    Odrv12 I__1773 (
            .O(N__8420),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    CascadeMux I__1772 (
            .O(N__8417),
            .I(N__8414));
    InMux I__1771 (
            .O(N__8414),
            .I(N__8408));
    InMux I__1770 (
            .O(N__8413),
            .I(N__8405));
    InMux I__1769 (
            .O(N__8412),
            .I(N__8402));
    InMux I__1768 (
            .O(N__8411),
            .I(N__8399));
    LocalMux I__1767 (
            .O(N__8408),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1766 (
            .O(N__8405),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1765 (
            .O(N__8402),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__1764 (
            .O(N__8399),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    InMux I__1763 (
            .O(N__8390),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__1762 (
            .O(N__8387),
            .I(N__8376));
    InMux I__1761 (
            .O(N__8386),
            .I(N__8376));
    InMux I__1760 (
            .O(N__8385),
            .I(N__8376));
    InMux I__1759 (
            .O(N__8384),
            .I(N__8373));
    InMux I__1758 (
            .O(N__8383),
            .I(N__8370));
    LocalMux I__1757 (
            .O(N__8376),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1756 (
            .O(N__8373),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__1755 (
            .O(N__8370),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    CascadeMux I__1754 (
            .O(N__8363),
            .I(N__8360));
    InMux I__1753 (
            .O(N__8360),
            .I(N__8357));
    LocalMux I__1752 (
            .O(N__8357),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ));
    InMux I__1751 (
            .O(N__8354),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__1750 (
            .O(N__8351),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__1749 (
            .O(N__8348),
            .I(N__8345));
    LocalMux I__1748 (
            .O(N__8345),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO ));
    CascadeMux I__1747 (
            .O(N__8342),
            .I(\U409_CIA.CLK_CIA6_3_cascade_ ));
    InMux I__1746 (
            .O(N__8339),
            .I(N__8336));
    LocalMux I__1745 (
            .O(N__8336),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_2_1 ));
    InMux I__1744 (
            .O(N__8333),
            .I(N__8330));
    LocalMux I__1743 (
            .O(N__8330),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0 ));
    CascadeMux I__1742 (
            .O(N__8327),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ));
    InMux I__1741 (
            .O(N__8324),
            .I(N__8318));
    InMux I__1740 (
            .O(N__8323),
            .I(N__8318));
    LocalMux I__1739 (
            .O(N__8318),
            .I(\U409_CIA.CIA_CLK_COUNT11_3 ));
    CascadeMux I__1738 (
            .O(N__8315),
            .I(\U409_CIA.CLK_CIA6_0_cascade_ ));
    InMux I__1737 (
            .O(N__8312),
            .I(N__8309));
    LocalMux I__1736 (
            .O(N__8309),
            .I(\U409_CIA.CLK_CIA6_3 ));
    CascadeMux I__1735 (
            .O(N__8306),
            .I(\U409_CIA.CLK_CIA6_cascade_ ));
    InMux I__1734 (
            .O(N__8303),
            .I(N__8300));
    LocalMux I__1733 (
            .O(N__8300),
            .I(\U409_CIA.CLK_CIA_RNOZ0Z_1 ));
    InMux I__1732 (
            .O(N__8297),
            .I(N__8294));
    LocalMux I__1731 (
            .O(N__8294),
            .I(N__8290));
    InMux I__1730 (
            .O(N__8293),
            .I(N__8287));
    Span4Mux_h I__1729 (
            .O(N__8290),
            .I(N__8284));
    LocalMux I__1728 (
            .O(N__8287),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    Odrv4 I__1727 (
            .O(N__8284),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__1726 (
            .O(N__8279),
            .I(N__8275));
    InMux I__1725 (
            .O(N__8278),
            .I(N__8272));
    LocalMux I__1724 (
            .O(N__8275),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    LocalMux I__1723 (
            .O(N__8272),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    CascadeMux I__1722 (
            .O(N__8267),
            .I(N__8263));
    InMux I__1721 (
            .O(N__8266),
            .I(N__8260));
    InMux I__1720 (
            .O(N__8263),
            .I(N__8257));
    LocalMux I__1719 (
            .O(N__8260),
            .I(N__8254));
    LocalMux I__1718 (
            .O(N__8257),
            .I(N__8251));
    Span4Mux_v I__1717 (
            .O(N__8254),
            .I(N__8248));
    Span4Mux_h I__1716 (
            .O(N__8251),
            .I(N__8245));
    Sp12to4 I__1715 (
            .O(N__8248),
            .I(N__8242));
    Span4Mux_v I__1714 (
            .O(N__8245),
            .I(N__8239));
    Span12Mux_h I__1713 (
            .O(N__8242),
            .I(N__8236));
    Span4Mux_h I__1712 (
            .O(N__8239),
            .I(N__8233));
    Odrv12 I__1711 (
            .O(N__8236),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ));
    Odrv4 I__1710 (
            .O(N__8233),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ));
    InMux I__1709 (
            .O(N__8228),
            .I(N__8224));
    InMux I__1708 (
            .O(N__8227),
            .I(N__8221));
    LocalMux I__1707 (
            .O(N__8224),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    LocalMux I__1706 (
            .O(N__8221),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    InMux I__1705 (
            .O(N__8216),
            .I(N__8208));
    InMux I__1704 (
            .O(N__8215),
            .I(N__8208));
    InMux I__1703 (
            .O(N__8214),
            .I(N__8203));
    InMux I__1702 (
            .O(N__8213),
            .I(N__8203));
    LocalMux I__1701 (
            .O(N__8208),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__1700 (
            .O(N__8203),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    CascadeMux I__1699 (
            .O(N__8198),
            .I(N__8194));
    InMux I__1698 (
            .O(N__8197),
            .I(N__8189));
    InMux I__1697 (
            .O(N__8194),
            .I(N__8184));
    InMux I__1696 (
            .O(N__8193),
            .I(N__8184));
    InMux I__1695 (
            .O(N__8192),
            .I(N__8181));
    LocalMux I__1694 (
            .O(N__8189),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__1693 (
            .O(N__8184),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__1692 (
            .O(N__8181),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__1691 (
            .O(N__8174),
            .I(N__8167));
    InMux I__1690 (
            .O(N__8173),
            .I(N__8167));
    InMux I__1689 (
            .O(N__8172),
            .I(N__8164));
    LocalMux I__1688 (
            .O(N__8167),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    LocalMux I__1687 (
            .O(N__8164),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    IoInMux I__1686 (
            .O(N__8159),
            .I(N__8156));
    LocalMux I__1685 (
            .O(N__8156),
            .I(N__8153));
    IoSpan4Mux I__1684 (
            .O(N__8153),
            .I(N__8150));
    Span4Mux_s3_v I__1683 (
            .O(N__8150),
            .I(N__8147));
    Sp12to4 I__1682 (
            .O(N__8147),
            .I(N__8144));
    Span12Mux_v I__1681 (
            .O(N__8144),
            .I(N__8140));
    InMux I__1680 (
            .O(N__8143),
            .I(N__8137));
    Odrv12 I__1679 (
            .O(N__8140),
            .I(TACK_OUT));
    LocalMux I__1678 (
            .O(N__8137),
            .I(TACK_OUT));
    InMux I__1677 (
            .O(N__8132),
            .I(N__8126));
    InMux I__1676 (
            .O(N__8131),
            .I(N__8123));
    InMux I__1675 (
            .O(N__8130),
            .I(N__8118));
    InMux I__1674 (
            .O(N__8129),
            .I(N__8118));
    LocalMux I__1673 (
            .O(N__8126),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1672 (
            .O(N__8123),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1671 (
            .O(N__8118),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    InMux I__1670 (
            .O(N__8111),
            .I(N__8106));
    InMux I__1669 (
            .O(N__8110),
            .I(N__8101));
    InMux I__1668 (
            .O(N__8109),
            .I(N__8101));
    LocalMux I__1667 (
            .O(N__8106),
            .I(\U409_TRANSFER_ACK.N_62 ));
    LocalMux I__1666 (
            .O(N__8101),
            .I(\U409_TRANSFER_ACK.N_62 ));
    SRMux I__1665 (
            .O(N__8096),
            .I(N__8093));
    LocalMux I__1664 (
            .O(N__8093),
            .I(N__8088));
    SRMux I__1663 (
            .O(N__8092),
            .I(N__8085));
    SRMux I__1662 (
            .O(N__8091),
            .I(N__8081));
    Span4Mux_v I__1661 (
            .O(N__8088),
            .I(N__8078));
    LocalMux I__1660 (
            .O(N__8085),
            .I(N__8075));
    SRMux I__1659 (
            .O(N__8084),
            .I(N__8072));
    LocalMux I__1658 (
            .O(N__8081),
            .I(N__8069));
    Span4Mux_v I__1657 (
            .O(N__8078),
            .I(N__8064));
    Span4Mux_v I__1656 (
            .O(N__8075),
            .I(N__8064));
    LocalMux I__1655 (
            .O(N__8072),
            .I(N__8061));
    Odrv4 I__1654 (
            .O(N__8069),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv4 I__1653 (
            .O(N__8064),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv4 I__1652 (
            .O(N__8061),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    InMux I__1651 (
            .O(N__8054),
            .I(N__8051));
    LocalMux I__1650 (
            .O(N__8051),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1 ));
    InMux I__1649 (
            .O(N__8048),
            .I(N__8045));
    LocalMux I__1648 (
            .O(N__8045),
            .I(N__8038));
    InMux I__1647 (
            .O(N__8044),
            .I(N__8035));
    InMux I__1646 (
            .O(N__8043),
            .I(N__8028));
    InMux I__1645 (
            .O(N__8042),
            .I(N__8028));
    InMux I__1644 (
            .O(N__8041),
            .I(N__8025));
    Span4Mux_v I__1643 (
            .O(N__8038),
            .I(N__8020));
    LocalMux I__1642 (
            .O(N__8035),
            .I(N__8020));
    InMux I__1641 (
            .O(N__8034),
            .I(N__8015));
    InMux I__1640 (
            .O(N__8033),
            .I(N__8015));
    LocalMux I__1639 (
            .O(N__8028),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1638 (
            .O(N__8025),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    Odrv4 I__1637 (
            .O(N__8020),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1636 (
            .O(N__8015),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    InMux I__1635 (
            .O(N__8006),
            .I(N__8002));
    InMux I__1634 (
            .O(N__8005),
            .I(N__7997));
    LocalMux I__1633 (
            .O(N__8002),
            .I(N__7994));
    InMux I__1632 (
            .O(N__8001),
            .I(N__7991));
    CascadeMux I__1631 (
            .O(N__8000),
            .I(N__7988));
    LocalMux I__1630 (
            .O(N__7997),
            .I(N__7980));
    Span4Mux_v I__1629 (
            .O(N__7994),
            .I(N__7980));
    LocalMux I__1628 (
            .O(N__7991),
            .I(N__7980));
    InMux I__1627 (
            .O(N__7988),
            .I(N__7975));
    InMux I__1626 (
            .O(N__7987),
            .I(N__7975));
    Odrv4 I__1625 (
            .O(N__7980),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1624 (
            .O(N__7975),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    InMux I__1623 (
            .O(N__7970),
            .I(N__7964));
    InMux I__1622 (
            .O(N__7969),
            .I(N__7964));
    LocalMux I__1621 (
            .O(N__7964),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    IoInMux I__1620 (
            .O(N__7961),
            .I(N__7958));
    LocalMux I__1619 (
            .O(N__7958),
            .I(N__7955));
    Span12Mux_s2_v I__1618 (
            .O(N__7955),
            .I(N__7952));
    Odrv12 I__1617 (
            .O(N__7952),
            .I(RESETn_c_i));
    CascadeMux I__1616 (
            .O(N__7949),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_ ));
    InMux I__1615 (
            .O(N__7946),
            .I(N__7943));
    LocalMux I__1614 (
            .O(N__7943),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a3_3 ));
    InMux I__1613 (
            .O(N__7940),
            .I(N__7937));
    LocalMux I__1612 (
            .O(N__7937),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3 ));
    InMux I__1611 (
            .O(N__7934),
            .I(N__7930));
    InMux I__1610 (
            .O(N__7933),
            .I(N__7926));
    LocalMux I__1609 (
            .O(N__7930),
            .I(N__7923));
    InMux I__1608 (
            .O(N__7929),
            .I(N__7920));
    LocalMux I__1607 (
            .O(N__7926),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    Odrv4 I__1606 (
            .O(N__7923),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    LocalMux I__1605 (
            .O(N__7920),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    CascadeMux I__1604 (
            .O(N__7913),
            .I(N__7910));
    InMux I__1603 (
            .O(N__7910),
            .I(N__7907));
    LocalMux I__1602 (
            .O(N__7907),
            .I(N__7904));
    Odrv4 I__1601 (
            .O(N__7904),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out ));
    InMux I__1600 (
            .O(N__7901),
            .I(N__7891));
    InMux I__1599 (
            .O(N__7900),
            .I(N__7891));
    InMux I__1598 (
            .O(N__7899),
            .I(N__7891));
    InMux I__1597 (
            .O(N__7898),
            .I(N__7888));
    LocalMux I__1596 (
            .O(N__7891),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__1595 (
            .O(N__7888),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    CascadeMux I__1594 (
            .O(N__7883),
            .I(N__7878));
    InMux I__1593 (
            .O(N__7882),
            .I(N__7872));
    InMux I__1592 (
            .O(N__7881),
            .I(N__7869));
    InMux I__1591 (
            .O(N__7878),
            .I(N__7866));
    InMux I__1590 (
            .O(N__7877),
            .I(N__7861));
    InMux I__1589 (
            .O(N__7876),
            .I(N__7861));
    InMux I__1588 (
            .O(N__7875),
            .I(N__7858));
    LocalMux I__1587 (
            .O(N__7872),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1586 (
            .O(N__7869),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1585 (
            .O(N__7866),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1584 (
            .O(N__7861),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1583 (
            .O(N__7858),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    InMux I__1582 (
            .O(N__7847),
            .I(N__7840));
    InMux I__1581 (
            .O(N__7846),
            .I(N__7837));
    InMux I__1580 (
            .O(N__7845),
            .I(N__7832));
    InMux I__1579 (
            .O(N__7844),
            .I(N__7832));
    InMux I__1578 (
            .O(N__7843),
            .I(N__7829));
    LocalMux I__1577 (
            .O(N__7840),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1576 (
            .O(N__7837),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1575 (
            .O(N__7832),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__1574 (
            .O(N__7829),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    CascadeMux I__1573 (
            .O(N__7820),
            .I(N__7814));
    CascadeMux I__1572 (
            .O(N__7819),
            .I(N__7811));
    InMux I__1571 (
            .O(N__7818),
            .I(N__7806));
    InMux I__1570 (
            .O(N__7817),
            .I(N__7806));
    InMux I__1569 (
            .O(N__7814),
            .I(N__7803));
    InMux I__1568 (
            .O(N__7811),
            .I(N__7800));
    LocalMux I__1567 (
            .O(N__7806),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__1566 (
            .O(N__7803),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__1565 (
            .O(N__7800),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    InMux I__1564 (
            .O(N__7793),
            .I(N__7782));
    InMux I__1563 (
            .O(N__7792),
            .I(N__7782));
    InMux I__1562 (
            .O(N__7791),
            .I(N__7782));
    InMux I__1561 (
            .O(N__7790),
            .I(N__7777));
    InMux I__1560 (
            .O(N__7789),
            .I(N__7777));
    LocalMux I__1559 (
            .O(N__7782),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__1558 (
            .O(N__7777),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    CascadeMux I__1557 (
            .O(N__7772),
            .I(N__7769));
    InMux I__1556 (
            .O(N__7769),
            .I(N__7762));
    InMux I__1555 (
            .O(N__7768),
            .I(N__7762));
    InMux I__1554 (
            .O(N__7767),
            .I(N__7759));
    LocalMux I__1553 (
            .O(N__7762),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__1552 (
            .O(N__7759),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    IoInMux I__1551 (
            .O(N__7754),
            .I(N__7751));
    LocalMux I__1550 (
            .O(N__7751),
            .I(N__7748));
    Span4Mux_s2_v I__1549 (
            .O(N__7748),
            .I(N__7745));
    Span4Mux_v I__1548 (
            .O(N__7745),
            .I(N__7742));
    Odrv4 I__1547 (
            .O(N__7742),
            .I(GB_BUFFER_CLK40_IN_c_g_THRU_CO));
    CascadeMux I__1546 (
            .O(N__7739),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ));
    InMux I__1545 (
            .O(N__7736),
            .I(N__7732));
    InMux I__1544 (
            .O(N__7735),
            .I(N__7729));
    LocalMux I__1543 (
            .O(N__7732),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__1542 (
            .O(N__7729),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    InMux I__1541 (
            .O(N__7724),
            .I(N__7721));
    LocalMux I__1540 (
            .O(N__7721),
            .I(N__7717));
    InMux I__1539 (
            .O(N__7720),
            .I(N__7714));
    Odrv12 I__1538 (
            .O(N__7717),
            .I(AC_TACK));
    LocalMux I__1537 (
            .O(N__7714),
            .I(AC_TACK));
    CascadeMux I__1536 (
            .O(N__7709),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ));
    CascadeMux I__1535 (
            .O(N__7706),
            .I(N__7703));
    InMux I__1534 (
            .O(N__7703),
            .I(N__7700));
    LocalMux I__1533 (
            .O(N__7700),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    InMux I__1532 (
            .O(N__7697),
            .I(N__7694));
    LocalMux I__1531 (
            .O(N__7694),
            .I(N__7691));
    Span12Mux_h I__1530 (
            .O(N__7691),
            .I(N__7688));
    Span12Mux_v I__1529 (
            .O(N__7688),
            .I(N__7685));
    Odrv12 I__1528 (
            .O(N__7685),
            .I(CPUCONFn_c));
    InMux I__1527 (
            .O(N__7682),
            .I(N__7679));
    LocalMux I__1526 (
            .O(N__7679),
            .I(\U409_AUTOCONFIG.AC_STARTZ0 ));
    InMux I__1525 (
            .O(N__7676),
            .I(N__7672));
    InMux I__1524 (
            .O(N__7675),
            .I(N__7669));
    LocalMux I__1523 (
            .O(N__7672),
            .I(\U409_AUTOCONFIG.STATE4 ));
    LocalMux I__1522 (
            .O(N__7669),
            .I(\U409_AUTOCONFIG.STATE4 ));
    InMux I__1521 (
            .O(N__7664),
            .I(N__7661));
    LocalMux I__1520 (
            .O(N__7661),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_0 ));
    InMux I__1519 (
            .O(N__7658),
            .I(N__7655));
    LocalMux I__1518 (
            .O(N__7655),
            .I(N__7647));
    InMux I__1517 (
            .O(N__7654),
            .I(N__7642));
    InMux I__1516 (
            .O(N__7653),
            .I(N__7642));
    InMux I__1515 (
            .O(N__7652),
            .I(N__7639));
    InMux I__1514 (
            .O(N__7651),
            .I(N__7634));
    InMux I__1513 (
            .O(N__7650),
            .I(N__7634));
    Odrv4 I__1512 (
            .O(N__7647),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__1511 (
            .O(N__7642),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__1510 (
            .O(N__7639),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    LocalMux I__1509 (
            .O(N__7634),
            .I(\U409_AUTOCONFIG.STATEZ0Z_0 ));
    CascadeMux I__1508 (
            .O(N__7625),
            .I(N__7617));
    InMux I__1507 (
            .O(N__7624),
            .I(N__7614));
    CascadeMux I__1506 (
            .O(N__7623),
            .I(N__7608));
    CascadeMux I__1505 (
            .O(N__7622),
            .I(N__7605));
    InMux I__1504 (
            .O(N__7621),
            .I(N__7601));
    InMux I__1503 (
            .O(N__7620),
            .I(N__7598));
    InMux I__1502 (
            .O(N__7617),
            .I(N__7595));
    LocalMux I__1501 (
            .O(N__7614),
            .I(N__7592));
    InMux I__1500 (
            .O(N__7613),
            .I(N__7589));
    CascadeMux I__1499 (
            .O(N__7612),
            .I(N__7586));
    InMux I__1498 (
            .O(N__7611),
            .I(N__7579));
    InMux I__1497 (
            .O(N__7608),
            .I(N__7579));
    InMux I__1496 (
            .O(N__7605),
            .I(N__7579));
    CascadeMux I__1495 (
            .O(N__7604),
            .I(N__7576));
    LocalMux I__1494 (
            .O(N__7601),
            .I(N__7569));
    LocalMux I__1493 (
            .O(N__7598),
            .I(N__7569));
    LocalMux I__1492 (
            .O(N__7595),
            .I(N__7566));
    Span4Mux_v I__1491 (
            .O(N__7592),
            .I(N__7561));
    LocalMux I__1490 (
            .O(N__7589),
            .I(N__7561));
    InMux I__1489 (
            .O(N__7586),
            .I(N__7558));
    LocalMux I__1488 (
            .O(N__7579),
            .I(N__7555));
    InMux I__1487 (
            .O(N__7576),
            .I(N__7550));
    InMux I__1486 (
            .O(N__7575),
            .I(N__7550));
    InMux I__1485 (
            .O(N__7574),
            .I(N__7547));
    Span4Mux_v I__1484 (
            .O(N__7569),
            .I(N__7542));
    Span4Mux_v I__1483 (
            .O(N__7566),
            .I(N__7542));
    Span4Mux_v I__1482 (
            .O(N__7561),
            .I(N__7539));
    LocalMux I__1481 (
            .O(N__7558),
            .I(N__7532));
    Sp12to4 I__1480 (
            .O(N__7555),
            .I(N__7532));
    LocalMux I__1479 (
            .O(N__7550),
            .I(N__7532));
    LocalMux I__1478 (
            .O(N__7547),
            .I(N__7525));
    Sp12to4 I__1477 (
            .O(N__7542),
            .I(N__7525));
    Sp12to4 I__1476 (
            .O(N__7539),
            .I(N__7525));
    Span12Mux_h I__1475 (
            .O(N__7532),
            .I(N__7522));
    Span12Mux_h I__1474 (
            .O(N__7525),
            .I(N__7519));
    Span12Mux_v I__1473 (
            .O(N__7522),
            .I(N__7516));
    Span12Mux_v I__1472 (
            .O(N__7519),
            .I(N__7513));
    Odrv12 I__1471 (
            .O(N__7516),
            .I(RnW_c));
    Odrv12 I__1470 (
            .O(N__7513),
            .I(RnW_c));
    InMux I__1469 (
            .O(N__7508),
            .I(N__7505));
    LocalMux I__1468 (
            .O(N__7505),
            .I(N__7497));
    InMux I__1467 (
            .O(N__7504),
            .I(N__7492));
    InMux I__1466 (
            .O(N__7503),
            .I(N__7492));
    InMux I__1465 (
            .O(N__7502),
            .I(N__7489));
    InMux I__1464 (
            .O(N__7501),
            .I(N__7486));
    InMux I__1463 (
            .O(N__7500),
            .I(N__7483));
    Odrv4 I__1462 (
            .O(N__7497),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__1461 (
            .O(N__7492),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__1460 (
            .O(N__7489),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__1459 (
            .O(N__7486),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    LocalMux I__1458 (
            .O(N__7483),
            .I(\U409_AUTOCONFIG.STATEZ0Z_1 ));
    InMux I__1457 (
            .O(N__7472),
            .I(N__7469));
    LocalMux I__1456 (
            .O(N__7469),
            .I(N__7465));
    InMux I__1455 (
            .O(N__7468),
            .I(N__7462));
    Span4Mux_h I__1454 (
            .O(N__7465),
            .I(N__7458));
    LocalMux I__1453 (
            .O(N__7462),
            .I(N__7455));
    InMux I__1452 (
            .O(N__7461),
            .I(N__7452));
    Odrv4 I__1451 (
            .O(N__7458),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    Odrv12 I__1450 (
            .O(N__7455),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    LocalMux I__1449 (
            .O(N__7452),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    InMux I__1448 (
            .O(N__7445),
            .I(N__7441));
    InMux I__1447 (
            .O(N__7444),
            .I(N__7438));
    LocalMux I__1446 (
            .O(N__7441),
            .I(N__7433));
    LocalMux I__1445 (
            .O(N__7438),
            .I(N__7433));
    Span4Mux_v I__1444 (
            .O(N__7433),
            .I(N__7430));
    Odrv4 I__1443 (
            .O(N__7430),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn));
    InMux I__1442 (
            .O(N__7427),
            .I(N__7424));
    LocalMux I__1441 (
            .O(N__7424),
            .I(N__7421));
    Sp12to4 I__1440 (
            .O(N__7421),
            .I(N__7418));
    Span12Mux_v I__1439 (
            .O(N__7418),
            .I(N__7415));
    Span12Mux_h I__1438 (
            .O(N__7415),
            .I(N__7412));
    Odrv12 I__1437 (
            .O(N__7412),
            .I(TACKn_in));
    InMux I__1436 (
            .O(N__7409),
            .I(N__7406));
    LocalMux I__1435 (
            .O(N__7406),
            .I(\U409_TRANSFER_ACK.N_53 ));
    CascadeMux I__1434 (
            .O(N__7403),
            .I(\U409_TRANSFER_ACK.N_53_cascade_ ));
    InMux I__1433 (
            .O(N__7400),
            .I(N__7397));
    LocalMux I__1432 (
            .O(N__7397),
            .I(N__7394));
    Span4Mux_v I__1431 (
            .O(N__7394),
            .I(N__7390));
    InMux I__1430 (
            .O(N__7393),
            .I(N__7387));
    Odrv4 I__1429 (
            .O(N__7390),
            .I(ATA_SPACE));
    LocalMux I__1428 (
            .O(N__7387),
            .I(ATA_SPACE));
    IoInMux I__1427 (
            .O(N__7382),
            .I(N__7379));
    LocalMux I__1426 (
            .O(N__7379),
            .I(N__7376));
    Span12Mux_s3_v I__1425 (
            .O(N__7376),
            .I(N__7373));
    Span12Mux_v I__1424 (
            .O(N__7373),
            .I(N__7370));
    Span12Mux_h I__1423 (
            .O(N__7370),
            .I(N__7367));
    Odrv12 I__1422 (
            .O(N__7367),
            .I(BUFENn_c));
    InMux I__1421 (
            .O(N__7364),
            .I(N__7361));
    LocalMux I__1420 (
            .O(N__7361),
            .I(N__7353));
    InMux I__1419 (
            .O(N__7360),
            .I(N__7348));
    InMux I__1418 (
            .O(N__7359),
            .I(N__7348));
    InMux I__1417 (
            .O(N__7358),
            .I(N__7345));
    InMux I__1416 (
            .O(N__7357),
            .I(N__7342));
    InMux I__1415 (
            .O(N__7356),
            .I(N__7339));
    Odrv4 I__1414 (
            .O(N__7353),
            .I(\U409_AUTOCONFIG.D_OUT_sm0_0 ));
    LocalMux I__1413 (
            .O(N__7348),
            .I(\U409_AUTOCONFIG.D_OUT_sm0_0 ));
    LocalMux I__1412 (
            .O(N__7345),
            .I(\U409_AUTOCONFIG.D_OUT_sm0_0 ));
    LocalMux I__1411 (
            .O(N__7342),
            .I(\U409_AUTOCONFIG.D_OUT_sm0_0 ));
    LocalMux I__1410 (
            .O(N__7339),
            .I(\U409_AUTOCONFIG.D_OUT_sm0_0 ));
    IoInMux I__1409 (
            .O(N__7328),
            .I(N__7325));
    LocalMux I__1408 (
            .O(N__7325),
            .I(N__7322));
    Span4Mux_s3_v I__1407 (
            .O(N__7322),
            .I(N__7319));
    Span4Mux_v I__1406 (
            .O(N__7319),
            .I(N__7316));
    Sp12to4 I__1405 (
            .O(N__7316),
            .I(N__7313));
    Span12Mux_h I__1404 (
            .O(N__7313),
            .I(N__7309));
    InMux I__1403 (
            .O(N__7312),
            .I(N__7306));
    Odrv12 I__1402 (
            .O(N__7309),
            .I(CONFIGENn_c));
    LocalMux I__1401 (
            .O(N__7306),
            .I(CONFIGENn_c));
    InMux I__1400 (
            .O(N__7301),
            .I(N__7298));
    LocalMux I__1399 (
            .O(N__7298),
            .I(N__7290));
    InMux I__1398 (
            .O(N__7297),
            .I(N__7287));
    InMux I__1397 (
            .O(N__7296),
            .I(N__7284));
    InMux I__1396 (
            .O(N__7295),
            .I(N__7277));
    InMux I__1395 (
            .O(N__7294),
            .I(N__7277));
    InMux I__1394 (
            .O(N__7293),
            .I(N__7277));
    Odrv4 I__1393 (
            .O(N__7290),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__1392 (
            .O(N__7287),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__1391 (
            .O(N__7284),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    LocalMux I__1390 (
            .O(N__7277),
            .I(\U409_AUTOCONFIG.LIDE_CONFZ0 ));
    InMux I__1389 (
            .O(N__7268),
            .I(N__7265));
    LocalMux I__1388 (
            .O(N__7265),
            .I(N__7260));
    CascadeMux I__1387 (
            .O(N__7264),
            .I(N__7257));
    CascadeMux I__1386 (
            .O(N__7263),
            .I(N__7251));
    Span4Mux_v I__1385 (
            .O(N__7260),
            .I(N__7245));
    InMux I__1384 (
            .O(N__7257),
            .I(N__7242));
    InMux I__1383 (
            .O(N__7256),
            .I(N__7237));
    InMux I__1382 (
            .O(N__7255),
            .I(N__7237));
    InMux I__1381 (
            .O(N__7254),
            .I(N__7234));
    InMux I__1380 (
            .O(N__7251),
            .I(N__7225));
    InMux I__1379 (
            .O(N__7250),
            .I(N__7225));
    InMux I__1378 (
            .O(N__7249),
            .I(N__7225));
    InMux I__1377 (
            .O(N__7248),
            .I(N__7225));
    Odrv4 I__1376 (
            .O(N__7245),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1375 (
            .O(N__7242),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1374 (
            .O(N__7237),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1373 (
            .O(N__7234),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    LocalMux I__1372 (
            .O(N__7225),
            .I(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ));
    InMux I__1371 (
            .O(N__7214),
            .I(N__7210));
    InMux I__1370 (
            .O(N__7213),
            .I(N__7207));
    LocalMux I__1369 (
            .O(N__7210),
            .I(N__7204));
    LocalMux I__1368 (
            .O(N__7207),
            .I(\U409_AUTOCONFIG.STATE_d_2 ));
    Odrv4 I__1367 (
            .O(N__7204),
            .I(\U409_AUTOCONFIG.STATE_d_2 ));
    InMux I__1366 (
            .O(N__7199),
            .I(N__7195));
    InMux I__1365 (
            .O(N__7198),
            .I(N__7192));
    LocalMux I__1364 (
            .O(N__7195),
            .I(N__7187));
    LocalMux I__1363 (
            .O(N__7192),
            .I(N__7187));
    Span12Mux_v I__1362 (
            .O(N__7187),
            .I(N__7184));
    Odrv12 I__1361 (
            .O(N__7184),
            .I(\U409_AUTOCONFIG.un1_AZ0Z_13 ));
    InMux I__1360 (
            .O(N__7181),
            .I(N__7178));
    LocalMux I__1359 (
            .O(N__7178),
            .I(N__7175));
    Span4Mux_h I__1358 (
            .O(N__7175),
            .I(N__7170));
    InMux I__1357 (
            .O(N__7174),
            .I(N__7167));
    InMux I__1356 (
            .O(N__7173),
            .I(N__7164));
    Odrv4 I__1355 (
            .O(N__7170),
            .I(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1 ));
    LocalMux I__1354 (
            .O(N__7167),
            .I(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1 ));
    LocalMux I__1353 (
            .O(N__7164),
            .I(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1 ));
    CascadeMux I__1352 (
            .O(N__7157),
            .I(N__7153));
    CascadeMux I__1351 (
            .O(N__7156),
            .I(N__7149));
    InMux I__1350 (
            .O(N__7153),
            .I(N__7146));
    InMux I__1349 (
            .O(N__7152),
            .I(N__7143));
    InMux I__1348 (
            .O(N__7149),
            .I(N__7138));
    LocalMux I__1347 (
            .O(N__7146),
            .I(N__7135));
    LocalMux I__1346 (
            .O(N__7143),
            .I(N__7132));
    InMux I__1345 (
            .O(N__7142),
            .I(N__7129));
    InMux I__1344 (
            .O(N__7141),
            .I(N__7126));
    LocalMux I__1343 (
            .O(N__7138),
            .I(N__7121));
    Span4Mux_v I__1342 (
            .O(N__7135),
            .I(N__7112));
    Span4Mux_v I__1341 (
            .O(N__7132),
            .I(N__7112));
    LocalMux I__1340 (
            .O(N__7129),
            .I(N__7112));
    LocalMux I__1339 (
            .O(N__7126),
            .I(N__7112));
    InMux I__1338 (
            .O(N__7125),
            .I(N__7109));
    CascadeMux I__1337 (
            .O(N__7124),
            .I(N__7106));
    Span4Mux_v I__1336 (
            .O(N__7121),
            .I(N__7099));
    Span4Mux_v I__1335 (
            .O(N__7112),
            .I(N__7096));
    LocalMux I__1334 (
            .O(N__7109),
            .I(N__7093));
    InMux I__1333 (
            .O(N__7106),
            .I(N__7084));
    InMux I__1332 (
            .O(N__7105),
            .I(N__7084));
    InMux I__1331 (
            .O(N__7104),
            .I(N__7084));
    InMux I__1330 (
            .O(N__7103),
            .I(N__7084));
    InMux I__1329 (
            .O(N__7102),
            .I(N__7081));
    Odrv4 I__1328 (
            .O(N__7099),
            .I(AUTOCONFIG_SPACE));
    Odrv4 I__1327 (
            .O(N__7096),
            .I(AUTOCONFIG_SPACE));
    Odrv4 I__1326 (
            .O(N__7093),
            .I(AUTOCONFIG_SPACE));
    LocalMux I__1325 (
            .O(N__7084),
            .I(AUTOCONFIG_SPACE));
    LocalMux I__1324 (
            .O(N__7081),
            .I(AUTOCONFIG_SPACE));
    InMux I__1323 (
            .O(N__7070),
            .I(N__7067));
    LocalMux I__1322 (
            .O(N__7067),
            .I(N__7059));
    InMux I__1321 (
            .O(N__7066),
            .I(N__7055));
    InMux I__1320 (
            .O(N__7065),
            .I(N__7050));
    InMux I__1319 (
            .O(N__7064),
            .I(N__7050));
    InMux I__1318 (
            .O(N__7063),
            .I(N__7047));
    InMux I__1317 (
            .O(N__7062),
            .I(N__7044));
    Span4Mux_h I__1316 (
            .O(N__7059),
            .I(N__7041));
    InMux I__1315 (
            .O(N__7058),
            .I(N__7038));
    LocalMux I__1314 (
            .O(N__7055),
            .I(CONFIGURED));
    LocalMux I__1313 (
            .O(N__7050),
            .I(CONFIGURED));
    LocalMux I__1312 (
            .O(N__7047),
            .I(CONFIGURED));
    LocalMux I__1311 (
            .O(N__7044),
            .I(CONFIGURED));
    Odrv4 I__1310 (
            .O(N__7041),
            .I(CONFIGURED));
    LocalMux I__1309 (
            .O(N__7038),
            .I(CONFIGURED));
    CascadeMux I__1308 (
            .O(N__7025),
            .I(N__7020));
    InMux I__1307 (
            .O(N__7024),
            .I(N__7013));
    InMux I__1306 (
            .O(N__7023),
            .I(N__7013));
    InMux I__1305 (
            .O(N__7020),
            .I(N__7013));
    LocalMux I__1304 (
            .O(N__7013),
            .I(N__7009));
    InMux I__1303 (
            .O(N__7012),
            .I(N__7006));
    Span4Mux_v I__1302 (
            .O(N__7009),
            .I(N__7003));
    LocalMux I__1301 (
            .O(N__7006),
            .I(N__7000));
    Odrv4 I__1300 (
            .O(N__7003),
            .I(\U409_AUTOCONFIG.N_192 ));
    Odrv4 I__1299 (
            .O(N__7000),
            .I(\U409_AUTOCONFIG.N_192 ));
    InMux I__1298 (
            .O(N__6995),
            .I(N__6992));
    LocalMux I__1297 (
            .O(N__6992),
            .I(N__6989));
    Odrv4 I__1296 (
            .O(N__6989),
            .I(\U409_AUTOCONFIG.PR_OUTZ0Z_1 ));
    CEMux I__1295 (
            .O(N__6986),
            .I(N__6982));
    CEMux I__1294 (
            .O(N__6985),
            .I(N__6979));
    LocalMux I__1293 (
            .O(N__6982),
            .I(N__6975));
    LocalMux I__1292 (
            .O(N__6979),
            .I(N__6972));
    CEMux I__1291 (
            .O(N__6978),
            .I(N__6969));
    Span4Mux_v I__1290 (
            .O(N__6975),
            .I(N__6966));
    Span4Mux_v I__1289 (
            .O(N__6972),
            .I(N__6963));
    LocalMux I__1288 (
            .O(N__6969),
            .I(N__6960));
    Odrv4 I__1287 (
            .O(N__6966),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ));
    Odrv4 I__1286 (
            .O(N__6963),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ));
    Odrv4 I__1285 (
            .O(N__6960),
            .I(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ));
    CascadeMux I__1284 (
            .O(N__6953),
            .I(N__6950));
    InMux I__1283 (
            .O(N__6950),
            .I(N__6947));
    LocalMux I__1282 (
            .O(N__6947),
            .I(N__6944));
    Odrv4 I__1281 (
            .O(N__6944),
            .I(\U409_AUTOCONFIG.N_184_0 ));
    InMux I__1280 (
            .O(N__6941),
            .I(N__6935));
    InMux I__1279 (
            .O(N__6940),
            .I(N__6935));
    LocalMux I__1278 (
            .O(N__6935),
            .I(\U409_AUTOCONFIG.N_167 ));
    InMux I__1277 (
            .O(N__6932),
            .I(N__6926));
    InMux I__1276 (
            .O(N__6931),
            .I(N__6926));
    LocalMux I__1275 (
            .O(N__6926),
            .I(\U409_AUTOCONFIG.N_213_i ));
    InMux I__1274 (
            .O(N__6923),
            .I(N__6919));
    InMux I__1273 (
            .O(N__6922),
            .I(N__6915));
    LocalMux I__1272 (
            .O(N__6919),
            .I(N__6912));
    InMux I__1271 (
            .O(N__6918),
            .I(N__6909));
    LocalMux I__1270 (
            .O(N__6915),
            .I(\U409_AUTOCONFIG.N_182_0 ));
    Odrv4 I__1269 (
            .O(N__6912),
            .I(\U409_AUTOCONFIG.N_182_0 ));
    LocalMux I__1268 (
            .O(N__6909),
            .I(\U409_AUTOCONFIG.N_182_0 ));
    InMux I__1267 (
            .O(N__6902),
            .I(N__6896));
    InMux I__1266 (
            .O(N__6901),
            .I(N__6896));
    LocalMux I__1265 (
            .O(N__6896),
            .I(N__6892));
    InMux I__1264 (
            .O(N__6895),
            .I(N__6889));
    Odrv4 I__1263 (
            .O(N__6892),
            .I(\U409_AUTOCONFIG.N_223 ));
    LocalMux I__1262 (
            .O(N__6889),
            .I(\U409_AUTOCONFIG.N_223 ));
    InMux I__1261 (
            .O(N__6884),
            .I(N__6881));
    LocalMux I__1260 (
            .O(N__6881),
            .I(\U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_0_0 ));
    CascadeMux I__1259 (
            .O(N__6878),
            .I(N__6875));
    InMux I__1258 (
            .O(N__6875),
            .I(N__6870));
    InMux I__1257 (
            .O(N__6874),
            .I(N__6867));
    InMux I__1256 (
            .O(N__6873),
            .I(N__6864));
    LocalMux I__1255 (
            .O(N__6870),
            .I(N__6859));
    LocalMux I__1254 (
            .O(N__6867),
            .I(N__6859));
    LocalMux I__1253 (
            .O(N__6864),
            .I(N__6853));
    Span4Mux_v I__1252 (
            .O(N__6859),
            .I(N__6850));
    InMux I__1251 (
            .O(N__6858),
            .I(N__6847));
    InMux I__1250 (
            .O(N__6857),
            .I(N__6844));
    CascadeMux I__1249 (
            .O(N__6856),
            .I(N__6841));
    Span4Mux_v I__1248 (
            .O(N__6853),
            .I(N__6837));
    Span4Mux_v I__1247 (
            .O(N__6850),
            .I(N__6834));
    LocalMux I__1246 (
            .O(N__6847),
            .I(N__6829));
    LocalMux I__1245 (
            .O(N__6844),
            .I(N__6829));
    InMux I__1244 (
            .O(N__6841),
            .I(N__6824));
    InMux I__1243 (
            .O(N__6840),
            .I(N__6824));
    Sp12to4 I__1242 (
            .O(N__6837),
            .I(N__6821));
    Span4Mux_v I__1241 (
            .O(N__6834),
            .I(N__6818));
    Span4Mux_v I__1240 (
            .O(N__6829),
            .I(N__6813));
    LocalMux I__1239 (
            .O(N__6824),
            .I(N__6813));
    Span12Mux_h I__1238 (
            .O(N__6821),
            .I(N__6810));
    Span4Mux_v I__1237 (
            .O(N__6818),
            .I(N__6807));
    Sp12to4 I__1236 (
            .O(N__6813),
            .I(N__6804));
    Span12Mux_v I__1235 (
            .O(N__6810),
            .I(N__6801));
    Sp12to4 I__1234 (
            .O(N__6807),
            .I(N__6796));
    Span12Mux_v I__1233 (
            .O(N__6804),
            .I(N__6796));
    Odrv12 I__1232 (
            .O(N__6801),
            .I(A_c_3));
    Odrv12 I__1231 (
            .O(N__6796),
            .I(A_c_3));
    InMux I__1230 (
            .O(N__6791),
            .I(N__6788));
    LocalMux I__1229 (
            .O(N__6788),
            .I(N__6785));
    Odrv4 I__1228 (
            .O(N__6785),
            .I(\U409_AUTOCONFIG.N_190 ));
    InMux I__1227 (
            .O(N__6782),
            .I(N__6773));
    InMux I__1226 (
            .O(N__6781),
            .I(N__6770));
    InMux I__1225 (
            .O(N__6780),
            .I(N__6765));
    InMux I__1224 (
            .O(N__6779),
            .I(N__6755));
    InMux I__1223 (
            .O(N__6778),
            .I(N__6755));
    InMux I__1222 (
            .O(N__6777),
            .I(N__6750));
    InMux I__1221 (
            .O(N__6776),
            .I(N__6750));
    LocalMux I__1220 (
            .O(N__6773),
            .I(N__6745));
    LocalMux I__1219 (
            .O(N__6770),
            .I(N__6745));
    InMux I__1218 (
            .O(N__6769),
            .I(N__6740));
    InMux I__1217 (
            .O(N__6768),
            .I(N__6740));
    LocalMux I__1216 (
            .O(N__6765),
            .I(N__6737));
    InMux I__1215 (
            .O(N__6764),
            .I(N__6732));
    InMux I__1214 (
            .O(N__6763),
            .I(N__6732));
    InMux I__1213 (
            .O(N__6762),
            .I(N__6729));
    InMux I__1212 (
            .O(N__6761),
            .I(N__6724));
    InMux I__1211 (
            .O(N__6760),
            .I(N__6724));
    LocalMux I__1210 (
            .O(N__6755),
            .I(N__6715));
    LocalMux I__1209 (
            .O(N__6750),
            .I(N__6715));
    Span4Mux_h I__1208 (
            .O(N__6745),
            .I(N__6715));
    LocalMux I__1207 (
            .O(N__6740),
            .I(N__6715));
    Span4Mux_v I__1206 (
            .O(N__6737),
            .I(N__6712));
    LocalMux I__1205 (
            .O(N__6732),
            .I(N__6707));
    LocalMux I__1204 (
            .O(N__6729),
            .I(N__6707));
    LocalMux I__1203 (
            .O(N__6724),
            .I(N__6704));
    Span4Mux_v I__1202 (
            .O(N__6715),
            .I(N__6701));
    Span4Mux_v I__1201 (
            .O(N__6712),
            .I(N__6694));
    Span4Mux_v I__1200 (
            .O(N__6707),
            .I(N__6694));
    Span4Mux_v I__1199 (
            .O(N__6704),
            .I(N__6694));
    Sp12to4 I__1198 (
            .O(N__6701),
            .I(N__6689));
    Sp12to4 I__1197 (
            .O(N__6694),
            .I(N__6689));
    Odrv12 I__1196 (
            .O(N__6689),
            .I(A_c_4));
    InMux I__1195 (
            .O(N__6686),
            .I(N__6680));
    InMux I__1194 (
            .O(N__6685),
            .I(N__6680));
    LocalMux I__1193 (
            .O(N__6680),
            .I(N__6668));
    InMux I__1192 (
            .O(N__6679),
            .I(N__6665));
    InMux I__1191 (
            .O(N__6678),
            .I(N__6662));
    InMux I__1190 (
            .O(N__6677),
            .I(N__6657));
    InMux I__1189 (
            .O(N__6676),
            .I(N__6657));
    InMux I__1188 (
            .O(N__6675),
            .I(N__6652));
    InMux I__1187 (
            .O(N__6674),
            .I(N__6652));
    InMux I__1186 (
            .O(N__6673),
            .I(N__6647));
    InMux I__1185 (
            .O(N__6672),
            .I(N__6647));
    InMux I__1184 (
            .O(N__6671),
            .I(N__6644));
    Span4Mux_v I__1183 (
            .O(N__6668),
            .I(N__6631));
    LocalMux I__1182 (
            .O(N__6665),
            .I(N__6631));
    LocalMux I__1181 (
            .O(N__6662),
            .I(N__6631));
    LocalMux I__1180 (
            .O(N__6657),
            .I(N__6631));
    LocalMux I__1179 (
            .O(N__6652),
            .I(N__6631));
    LocalMux I__1178 (
            .O(N__6647),
            .I(N__6626));
    LocalMux I__1177 (
            .O(N__6644),
            .I(N__6626));
    InMux I__1176 (
            .O(N__6643),
            .I(N__6623));
    InMux I__1175 (
            .O(N__6642),
            .I(N__6620));
    Span4Mux_v I__1174 (
            .O(N__6631),
            .I(N__6617));
    Span4Mux_v I__1173 (
            .O(N__6626),
            .I(N__6614));
    LocalMux I__1172 (
            .O(N__6623),
            .I(N__6609));
    LocalMux I__1171 (
            .O(N__6620),
            .I(N__6609));
    Sp12to4 I__1170 (
            .O(N__6617),
            .I(N__6604));
    Sp12to4 I__1169 (
            .O(N__6614),
            .I(N__6604));
    Span12Mux_h I__1168 (
            .O(N__6609),
            .I(N__6601));
    Span12Mux_h I__1167 (
            .O(N__6604),
            .I(N__6598));
    Span12Mux_v I__1166 (
            .O(N__6601),
            .I(N__6595));
    Span12Mux_v I__1165 (
            .O(N__6598),
            .I(N__6592));
    Odrv12 I__1164 (
            .O(N__6595),
            .I(A_c_1));
    Odrv12 I__1163 (
            .O(N__6592),
            .I(A_c_1));
    CascadeMux I__1162 (
            .O(N__6587),
            .I(N__6579));
    InMux I__1161 (
            .O(N__6586),
            .I(N__6571));
    InMux I__1160 (
            .O(N__6585),
            .I(N__6571));
    InMux I__1159 (
            .O(N__6584),
            .I(N__6566));
    InMux I__1158 (
            .O(N__6583),
            .I(N__6566));
    InMux I__1157 (
            .O(N__6582),
            .I(N__6563));
    InMux I__1156 (
            .O(N__6579),
            .I(N__6559));
    InMux I__1155 (
            .O(N__6578),
            .I(N__6556));
    InMux I__1154 (
            .O(N__6577),
            .I(N__6551));
    InMux I__1153 (
            .O(N__6576),
            .I(N__6551));
    LocalMux I__1152 (
            .O(N__6571),
            .I(N__6546));
    LocalMux I__1151 (
            .O(N__6566),
            .I(N__6546));
    LocalMux I__1150 (
            .O(N__6563),
            .I(N__6543));
    CascadeMux I__1149 (
            .O(N__6562),
            .I(N__6540));
    LocalMux I__1148 (
            .O(N__6559),
            .I(N__6533));
    LocalMux I__1147 (
            .O(N__6556),
            .I(N__6533));
    LocalMux I__1146 (
            .O(N__6551),
            .I(N__6533));
    Span4Mux_v I__1145 (
            .O(N__6546),
            .I(N__6526));
    Span4Mux_v I__1144 (
            .O(N__6543),
            .I(N__6523));
    InMux I__1143 (
            .O(N__6540),
            .I(N__6520));
    Span4Mux_v I__1142 (
            .O(N__6533),
            .I(N__6517));
    InMux I__1141 (
            .O(N__6532),
            .I(N__6512));
    InMux I__1140 (
            .O(N__6531),
            .I(N__6512));
    InMux I__1139 (
            .O(N__6530),
            .I(N__6507));
    InMux I__1138 (
            .O(N__6529),
            .I(N__6507));
    Sp12to4 I__1137 (
            .O(N__6526),
            .I(N__6494));
    Sp12to4 I__1136 (
            .O(N__6523),
            .I(N__6494));
    LocalMux I__1135 (
            .O(N__6520),
            .I(N__6494));
    Sp12to4 I__1134 (
            .O(N__6517),
            .I(N__6494));
    LocalMux I__1133 (
            .O(N__6512),
            .I(N__6494));
    LocalMux I__1132 (
            .O(N__6507),
            .I(N__6494));
    Span12Mux_h I__1131 (
            .O(N__6494),
            .I(N__6491));
    Span12Mux_v I__1130 (
            .O(N__6491),
            .I(N__6488));
    Odrv12 I__1129 (
            .O(N__6488),
            .I(A_c_2));
    InMux I__1128 (
            .O(N__6485),
            .I(N__6479));
    InMux I__1127 (
            .O(N__6484),
            .I(N__6476));
    CascadeMux I__1126 (
            .O(N__6483),
            .I(N__6473));
    CascadeMux I__1125 (
            .O(N__6482),
            .I(N__6470));
    LocalMux I__1124 (
            .O(N__6479),
            .I(N__6465));
    LocalMux I__1123 (
            .O(N__6476),
            .I(N__6462));
    InMux I__1122 (
            .O(N__6473),
            .I(N__6457));
    InMux I__1121 (
            .O(N__6470),
            .I(N__6457));
    CascadeMux I__1120 (
            .O(N__6469),
            .I(N__6452));
    InMux I__1119 (
            .O(N__6468),
            .I(N__6449));
    Span4Mux_v I__1118 (
            .O(N__6465),
            .I(N__6442));
    Span4Mux_v I__1117 (
            .O(N__6462),
            .I(N__6442));
    LocalMux I__1116 (
            .O(N__6457),
            .I(N__6442));
    InMux I__1115 (
            .O(N__6456),
            .I(N__6439));
    InMux I__1114 (
            .O(N__6455),
            .I(N__6434));
    InMux I__1113 (
            .O(N__6452),
            .I(N__6434));
    LocalMux I__1112 (
            .O(N__6449),
            .I(\U409_AUTOCONFIG.N_198 ));
    Odrv4 I__1111 (
            .O(N__6442),
            .I(\U409_AUTOCONFIG.N_198 ));
    LocalMux I__1110 (
            .O(N__6439),
            .I(\U409_AUTOCONFIG.N_198 ));
    LocalMux I__1109 (
            .O(N__6434),
            .I(\U409_AUTOCONFIG.N_198 ));
    InMux I__1108 (
            .O(N__6425),
            .I(N__6419));
    InMux I__1107 (
            .O(N__6424),
            .I(N__6419));
    LocalMux I__1106 (
            .O(N__6419),
            .I(N__6416));
    Odrv4 I__1105 (
            .O(N__6416),
            .I(\U409_AUTOCONFIG.N_222 ));
    CascadeMux I__1104 (
            .O(N__6413),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNIMM061Z0Z_0_cascade_ ));
    IoInMux I__1103 (
            .O(N__6410),
            .I(N__6407));
    LocalMux I__1102 (
            .O(N__6407),
            .I(N__6404));
    IoSpan4Mux I__1101 (
            .O(N__6404),
            .I(N__6401));
    Sp12to4 I__1100 (
            .O(N__6401),
            .I(N__6398));
    Span12Mux_s7_v I__1099 (
            .O(N__6398),
            .I(N__6395));
    Odrv12 I__1098 (
            .O(N__6395),
            .I(D_OUT_0));
    InMux I__1097 (
            .O(N__6392),
            .I(N__6389));
    LocalMux I__1096 (
            .O(N__6389),
            .I(N__6386));
    Odrv12 I__1095 (
            .O(N__6386),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ));
    InMux I__1094 (
            .O(N__6383),
            .I(N__6380));
    LocalMux I__1093 (
            .O(N__6380),
            .I(N__6377));
    Odrv4 I__1092 (
            .O(N__6377),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ));
    InMux I__1091 (
            .O(N__6374),
            .I(N__6365));
    InMux I__1090 (
            .O(N__6373),
            .I(N__6365));
    InMux I__1089 (
            .O(N__6372),
            .I(N__6365));
    LocalMux I__1088 (
            .O(N__6365),
            .I(N__6361));
    InMux I__1087 (
            .O(N__6364),
            .I(N__6358));
    Odrv4 I__1086 (
            .O(N__6361),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxaZ0Z_1 ));
    LocalMux I__1085 (
            .O(N__6358),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxaZ0Z_1 ));
    InMux I__1084 (
            .O(N__6353),
            .I(N__6350));
    LocalMux I__1083 (
            .O(N__6350),
            .I(N__6347));
    Span4Mux_v I__1082 (
            .O(N__6347),
            .I(N__6344));
    Sp12to4 I__1081 (
            .O(N__6344),
            .I(N__6341));
    Span12Mux_h I__1080 (
            .O(N__6341),
            .I(N__6338));
    Span12Mux_h I__1079 (
            .O(N__6338),
            .I(N__6335));
    Span12Mux_v I__1078 (
            .O(N__6335),
            .I(N__6332));
    Odrv12 I__1077 (
            .O(N__6332),
            .I(AUTOBOOT_c));
    InMux I__1076 (
            .O(N__6329),
            .I(N__6326));
    LocalMux I__1075 (
            .O(N__6326),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ));
    InMux I__1074 (
            .O(N__6323),
            .I(N__6320));
    LocalMux I__1073 (
            .O(N__6320),
            .I(\U409_AUTOCONFIG.PR_OUTZ0Z_0 ));
    CascadeMux I__1072 (
            .O(N__6317),
            .I(N__6314));
    InMux I__1071 (
            .O(N__6314),
            .I(N__6311));
    LocalMux I__1070 (
            .O(N__6311),
            .I(N__6308));
    Span4Mux_v I__1069 (
            .O(N__6308),
            .I(N__6304));
    InMux I__1068 (
            .O(N__6307),
            .I(N__6301));
    Odrv4 I__1067 (
            .O(N__6304),
            .I(\U409_AUTOCONFIG.N_214_0 ));
    LocalMux I__1066 (
            .O(N__6301),
            .I(\U409_AUTOCONFIG.N_214_0 ));
    InMux I__1065 (
            .O(N__6296),
            .I(N__6290));
    InMux I__1064 (
            .O(N__6295),
            .I(N__6290));
    LocalMux I__1063 (
            .O(N__6290),
            .I(N__6287));
    Span4Mux_v I__1062 (
            .O(N__6287),
            .I(N__6282));
    InMux I__1061 (
            .O(N__6286),
            .I(N__6279));
    InMux I__1060 (
            .O(N__6285),
            .I(N__6276));
    Odrv4 I__1059 (
            .O(N__6282),
            .I(\U409_AUTOCONFIG.N_193_1 ));
    LocalMux I__1058 (
            .O(N__6279),
            .I(\U409_AUTOCONFIG.N_193_1 ));
    LocalMux I__1057 (
            .O(N__6276),
            .I(\U409_AUTOCONFIG.N_193_1 ));
    InMux I__1056 (
            .O(N__6269),
            .I(N__6266));
    LocalMux I__1055 (
            .O(N__6266),
            .I(N__6263));
    Odrv4 I__1054 (
            .O(N__6263),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ));
    InMux I__1053 (
            .O(N__6260),
            .I(N__6254));
    InMux I__1052 (
            .O(N__6259),
            .I(N__6254));
    LocalMux I__1051 (
            .O(N__6254),
            .I(N__6251));
    Span4Mux_v I__1050 (
            .O(N__6251),
            .I(N__6248));
    Odrv4 I__1049 (
            .O(N__6248),
            .I(\U409_AUTOCONFIG.N_159 ));
    CascadeMux I__1048 (
            .O(N__6245),
            .I(N__6242));
    InMux I__1047 (
            .O(N__6242),
            .I(N__6239));
    LocalMux I__1046 (
            .O(N__6239),
            .I(N__6235));
    CascadeMux I__1045 (
            .O(N__6238),
            .I(N__6232));
    Span4Mux_v I__1044 (
            .O(N__6235),
            .I(N__6229));
    InMux I__1043 (
            .O(N__6232),
            .I(N__6226));
    Odrv4 I__1042 (
            .O(N__6229),
            .I(\U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_2 ));
    LocalMux I__1041 (
            .O(N__6226),
            .I(\U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_2 ));
    InMux I__1040 (
            .O(N__6221),
            .I(N__6218));
    LocalMux I__1039 (
            .O(N__6218),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ));
    InMux I__1038 (
            .O(N__6215),
            .I(N__6212));
    LocalMux I__1037 (
            .O(N__6212),
            .I(N__6209));
    Odrv4 I__1036 (
            .O(N__6209),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ));
    InMux I__1035 (
            .O(N__6206),
            .I(N__6203));
    LocalMux I__1034 (
            .O(N__6203),
            .I(N__6200));
    Odrv4 I__1033 (
            .O(N__6200),
            .I(\U409_AUTOCONFIG.PR_OUTZ0Z_2 ));
    CascadeMux I__1032 (
            .O(N__6197),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2_cascade_ ));
    IoInMux I__1031 (
            .O(N__6194),
            .I(N__6191));
    LocalMux I__1030 (
            .O(N__6191),
            .I(N__6188));
    Span12Mux_s8_v I__1029 (
            .O(N__6188),
            .I(N__6185));
    Odrv12 I__1028 (
            .O(N__6185),
            .I(D_OUT_2));
    InMux I__1027 (
            .O(N__6182),
            .I(N__6174));
    InMux I__1026 (
            .O(N__6181),
            .I(N__6174));
    CascadeMux I__1025 (
            .O(N__6180),
            .I(N__6171));
    InMux I__1024 (
            .O(N__6179),
            .I(N__6167));
    LocalMux I__1023 (
            .O(N__6174),
            .I(N__6164));
    InMux I__1022 (
            .O(N__6171),
            .I(N__6161));
    InMux I__1021 (
            .O(N__6170),
            .I(N__6158));
    LocalMux I__1020 (
            .O(N__6167),
            .I(\U409_AUTOCONFIG.LIDE_BASE_10 ));
    Odrv12 I__1019 (
            .O(N__6164),
            .I(\U409_AUTOCONFIG.LIDE_BASE_10 ));
    LocalMux I__1018 (
            .O(N__6161),
            .I(\U409_AUTOCONFIG.LIDE_BASE_10 ));
    LocalMux I__1017 (
            .O(N__6158),
            .I(\U409_AUTOCONFIG.LIDE_BASE_10 ));
    InMux I__1016 (
            .O(N__6149),
            .I(N__6146));
    LocalMux I__1015 (
            .O(N__6146),
            .I(N__6143));
    Span4Mux_h I__1014 (
            .O(N__6143),
            .I(N__6139));
    InMux I__1013 (
            .O(N__6142),
            .I(N__6136));
    Span4Mux_v I__1012 (
            .O(N__6139),
            .I(N__6133));
    LocalMux I__1011 (
            .O(N__6136),
            .I(N__6130));
    Span4Mux_v I__1010 (
            .O(N__6133),
            .I(N__6127));
    Span12Mux_h I__1009 (
            .O(N__6130),
            .I(N__6124));
    Odrv4 I__1008 (
            .O(N__6127),
            .I(D_in_7));
    Odrv12 I__1007 (
            .O(N__6124),
            .I(D_in_7));
    CascadeMux I__1006 (
            .O(N__6119),
            .I(\U409_AUTOCONFIG.LIDE_BASE_10_cascade_ ));
    CascadeMux I__1005 (
            .O(N__6116),
            .I(N__6113));
    InMux I__1004 (
            .O(N__6113),
            .I(N__6110));
    LocalMux I__1003 (
            .O(N__6110),
            .I(N__6107));
    Odrv12 I__1002 (
            .O(N__6107),
            .I(\U409_AUTOCONFIG.N_78 ));
    InMux I__1001 (
            .O(N__6104),
            .I(N__6100));
    InMux I__1000 (
            .O(N__6103),
            .I(N__6091));
    LocalMux I__999 (
            .O(N__6100),
            .I(N__6088));
    InMux I__998 (
            .O(N__6099),
            .I(N__6085));
    InMux I__997 (
            .O(N__6098),
            .I(N__6082));
    InMux I__996 (
            .O(N__6097),
            .I(N__6075));
    InMux I__995 (
            .O(N__6096),
            .I(N__6075));
    InMux I__994 (
            .O(N__6095),
            .I(N__6075));
    InMux I__993 (
            .O(N__6094),
            .I(N__6072));
    LocalMux I__992 (
            .O(N__6091),
            .I(\U409_AUTOCONFIG.LIDE_BASE_10_2 ));
    Odrv12 I__991 (
            .O(N__6088),
            .I(\U409_AUTOCONFIG.LIDE_BASE_10_2 ));
    LocalMux I__990 (
            .O(N__6085),
            .I(\U409_AUTOCONFIG.LIDE_BASE_10_2 ));
    LocalMux I__989 (
            .O(N__6082),
            .I(\U409_AUTOCONFIG.LIDE_BASE_10_2 ));
    LocalMux I__988 (
            .O(N__6075),
            .I(\U409_AUTOCONFIG.LIDE_BASE_10_2 ));
    LocalMux I__987 (
            .O(N__6072),
            .I(\U409_AUTOCONFIG.LIDE_BASE_10_2 ));
    CascadeMux I__986 (
            .O(N__6059),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNIOO061Z0Z_1_cascade_ ));
    IoInMux I__985 (
            .O(N__6056),
            .I(N__6053));
    LocalMux I__984 (
            .O(N__6053),
            .I(N__6050));
    Span12Mux_s6_v I__983 (
            .O(N__6050),
            .I(N__6047));
    Odrv12 I__982 (
            .O(N__6047),
            .I(D_OUT_1));
    InMux I__981 (
            .O(N__6044),
            .I(N__6041));
    LocalMux I__980 (
            .O(N__6041),
            .I(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ));
    InMux I__979 (
            .O(N__6038),
            .I(N__6032));
    InMux I__978 (
            .O(N__6037),
            .I(N__6032));
    LocalMux I__977 (
            .O(N__6032),
            .I(\U409_AUTOCONFIG.N_225 ));
    CascadeMux I__976 (
            .O(N__6029),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_3_cascade_ ));
    InMux I__975 (
            .O(N__6026),
            .I(N__6023));
    LocalMux I__974 (
            .O(N__6023),
            .I(N__6020));
    Odrv4 I__973 (
            .O(N__6020),
            .I(\U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_3 ));
    InMux I__972 (
            .O(N__6017),
            .I(N__6010));
    InMux I__971 (
            .O(N__6016),
            .I(N__6003));
    InMux I__970 (
            .O(N__6015),
            .I(N__6003));
    InMux I__969 (
            .O(N__6014),
            .I(N__6003));
    CascadeMux I__968 (
            .O(N__6013),
            .I(N__5998));
    LocalMux I__967 (
            .O(N__6010),
            .I(N__5993));
    LocalMux I__966 (
            .O(N__6003),
            .I(N__5993));
    InMux I__965 (
            .O(N__6002),
            .I(N__5990));
    InMux I__964 (
            .O(N__6001),
            .I(N__5985));
    InMux I__963 (
            .O(N__5998),
            .I(N__5985));
    Span4Mux_v I__962 (
            .O(N__5993),
            .I(N__5980));
    LocalMux I__961 (
            .O(N__5990),
            .I(N__5980));
    LocalMux I__960 (
            .O(N__5985),
            .I(N__5975));
    Sp12to4 I__959 (
            .O(N__5980),
            .I(N__5975));
    Odrv12 I__958 (
            .O(N__5975),
            .I(A_c_6));
    CascadeMux I__957 (
            .O(N__5972),
            .I(N__5969));
    InMux I__956 (
            .O(N__5969),
            .I(N__5966));
    LocalMux I__955 (
            .O(N__5966),
            .I(N__5961));
    InMux I__954 (
            .O(N__5965),
            .I(N__5956));
    InMux I__953 (
            .O(N__5964),
            .I(N__5956));
    Span4Mux_v I__952 (
            .O(N__5961),
            .I(N__5950));
    LocalMux I__951 (
            .O(N__5956),
            .I(N__5950));
    CascadeMux I__950 (
            .O(N__5955),
            .I(N__5946));
    Span4Mux_v I__949 (
            .O(N__5950),
            .I(N__5941));
    InMux I__948 (
            .O(N__5949),
            .I(N__5938));
    InMux I__947 (
            .O(N__5946),
            .I(N__5931));
    InMux I__946 (
            .O(N__5945),
            .I(N__5931));
    InMux I__945 (
            .O(N__5944),
            .I(N__5931));
    Sp12to4 I__944 (
            .O(N__5941),
            .I(N__5924));
    LocalMux I__943 (
            .O(N__5938),
            .I(N__5924));
    LocalMux I__942 (
            .O(N__5931),
            .I(N__5924));
    Span12Mux_h I__941 (
            .O(N__5924),
            .I(N__5921));
    Odrv12 I__940 (
            .O(N__5921),
            .I(A_c_7));
    InMux I__939 (
            .O(N__5918),
            .I(N__5914));
    InMux I__938 (
            .O(N__5917),
            .I(N__5911));
    LocalMux I__937 (
            .O(N__5914),
            .I(N__5908));
    LocalMux I__936 (
            .O(N__5911),
            .I(\U409_AUTOCONFIG.un1_A_13Z0Z_3 ));
    Odrv4 I__935 (
            .O(N__5908),
            .I(\U409_AUTOCONFIG.un1_A_13Z0Z_3 ));
    CascadeMux I__934 (
            .O(N__5903),
            .I(\U409_AUTOCONFIG.un1_A_13Z0Z_0_cascade_ ));
    InMux I__933 (
            .O(N__5900),
            .I(N__5897));
    LocalMux I__932 (
            .O(N__5897),
            .I(\U409_AUTOCONFIG.N_70 ));
    InMux I__931 (
            .O(N__5894),
            .I(N__5890));
    InMux I__930 (
            .O(N__5893),
            .I(N__5887));
    LocalMux I__929 (
            .O(N__5890),
            .I(LIDE_BASE_7));
    LocalMux I__928 (
            .O(N__5887),
            .I(LIDE_BASE_7));
    InMux I__927 (
            .O(N__5882),
            .I(N__5879));
    LocalMux I__926 (
            .O(N__5879),
            .I(\U409_AUTOCONFIG.N_74 ));
    InMux I__925 (
            .O(N__5876),
            .I(N__5872));
    InMux I__924 (
            .O(N__5875),
            .I(N__5868));
    LocalMux I__923 (
            .O(N__5872),
            .I(N__5864));
    CascadeMux I__922 (
            .O(N__5871),
            .I(N__5861));
    LocalMux I__921 (
            .O(N__5868),
            .I(N__5858));
    InMux I__920 (
            .O(N__5867),
            .I(N__5855));
    Span4Mux_v I__919 (
            .O(N__5864),
            .I(N__5850));
    InMux I__918 (
            .O(N__5861),
            .I(N__5847));
    Span4Mux_v I__917 (
            .O(N__5858),
            .I(N__5844));
    LocalMux I__916 (
            .O(N__5855),
            .I(N__5841));
    InMux I__915 (
            .O(N__5854),
            .I(N__5836));
    InMux I__914 (
            .O(N__5853),
            .I(N__5836));
    Sp12to4 I__913 (
            .O(N__5850),
            .I(N__5830));
    LocalMux I__912 (
            .O(N__5847),
            .I(N__5830));
    Span4Mux_v I__911 (
            .O(N__5844),
            .I(N__5827));
    Span4Mux_h I__910 (
            .O(N__5841),
            .I(N__5822));
    LocalMux I__909 (
            .O(N__5836),
            .I(N__5822));
    InMux I__908 (
            .O(N__5835),
            .I(N__5819));
    Span12Mux_h I__907 (
            .O(N__5830),
            .I(N__5816));
    Span4Mux_v I__906 (
            .O(N__5827),
            .I(N__5813));
    Sp12to4 I__905 (
            .O(N__5822),
            .I(N__5808));
    LocalMux I__904 (
            .O(N__5819),
            .I(N__5808));
    Span12Mux_v I__903 (
            .O(N__5816),
            .I(N__5805));
    Sp12to4 I__902 (
            .O(N__5813),
            .I(N__5800));
    Span12Mux_v I__901 (
            .O(N__5808),
            .I(N__5800));
    Odrv12 I__900 (
            .O(N__5805),
            .I(A_c_22));
    Odrv12 I__899 (
            .O(N__5800),
            .I(A_c_22));
    CascadeMux I__898 (
            .O(N__5795),
            .I(N__5789));
    CascadeMux I__897 (
            .O(N__5794),
            .I(N__5786));
    CascadeMux I__896 (
            .O(N__5793),
            .I(N__5783));
    InMux I__895 (
            .O(N__5792),
            .I(N__5778));
    InMux I__894 (
            .O(N__5789),
            .I(N__5774));
    InMux I__893 (
            .O(N__5786),
            .I(N__5767));
    InMux I__892 (
            .O(N__5783),
            .I(N__5764));
    CascadeMux I__891 (
            .O(N__5782),
            .I(N__5761));
    CascadeMux I__890 (
            .O(N__5781),
            .I(N__5758));
    LocalMux I__889 (
            .O(N__5778),
            .I(N__5755));
    InMux I__888 (
            .O(N__5777),
            .I(N__5752));
    LocalMux I__887 (
            .O(N__5774),
            .I(N__5749));
    InMux I__886 (
            .O(N__5773),
            .I(N__5746));
    InMux I__885 (
            .O(N__5772),
            .I(N__5741));
    InMux I__884 (
            .O(N__5771),
            .I(N__5741));
    InMux I__883 (
            .O(N__5770),
            .I(N__5737));
    LocalMux I__882 (
            .O(N__5767),
            .I(N__5732));
    LocalMux I__881 (
            .O(N__5764),
            .I(N__5732));
    InMux I__880 (
            .O(N__5761),
            .I(N__5729));
    InMux I__879 (
            .O(N__5758),
            .I(N__5726));
    Span4Mux_h I__878 (
            .O(N__5755),
            .I(N__5721));
    LocalMux I__877 (
            .O(N__5752),
            .I(N__5721));
    Span4Mux_v I__876 (
            .O(N__5749),
            .I(N__5714));
    LocalMux I__875 (
            .O(N__5746),
            .I(N__5714));
    LocalMux I__874 (
            .O(N__5741),
            .I(N__5714));
    CascadeMux I__873 (
            .O(N__5740),
            .I(N__5711));
    LocalMux I__872 (
            .O(N__5737),
            .I(N__5702));
    Sp12to4 I__871 (
            .O(N__5732),
            .I(N__5702));
    LocalMux I__870 (
            .O(N__5729),
            .I(N__5702));
    LocalMux I__869 (
            .O(N__5726),
            .I(N__5702));
    Span4Mux_v I__868 (
            .O(N__5721),
            .I(N__5699));
    Span4Mux_v I__867 (
            .O(N__5714),
            .I(N__5696));
    InMux I__866 (
            .O(N__5711),
            .I(N__5693));
    Span12Mux_v I__865 (
            .O(N__5702),
            .I(N__5684));
    Sp12to4 I__864 (
            .O(N__5699),
            .I(N__5684));
    Sp12to4 I__863 (
            .O(N__5696),
            .I(N__5684));
    LocalMux I__862 (
            .O(N__5693),
            .I(N__5684));
    Odrv12 I__861 (
            .O(N__5684),
            .I(A_c_21));
    CascadeMux I__860 (
            .O(N__5681),
            .I(N__5678));
    InMux I__859 (
            .O(N__5678),
            .I(N__5675));
    LocalMux I__858 (
            .O(N__5675),
            .I(N__5671));
    InMux I__857 (
            .O(N__5674),
            .I(N__5668));
    Odrv4 I__856 (
            .O(N__5671),
            .I(LIDE_BASE_5));
    LocalMux I__855 (
            .O(N__5668),
            .I(LIDE_BASE_5));
    InMux I__854 (
            .O(N__5663),
            .I(N__5660));
    LocalMux I__853 (
            .O(N__5660),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ));
    InMux I__852 (
            .O(N__5657),
            .I(N__5654));
    LocalMux I__851 (
            .O(N__5654),
            .I(N__5651));
    Odrv4 I__850 (
            .O(N__5651),
            .I(\U409_AUTOCONFIG.N_72 ));
    CascadeMux I__849 (
            .O(N__5648),
            .I(N__5642));
    CascadeMux I__848 (
            .O(N__5647),
            .I(N__5638));
    CascadeMux I__847 (
            .O(N__5646),
            .I(N__5635));
    CascadeMux I__846 (
            .O(N__5645),
            .I(N__5630));
    InMux I__845 (
            .O(N__5642),
            .I(N__5623));
    InMux I__844 (
            .O(N__5641),
            .I(N__5623));
    InMux I__843 (
            .O(N__5638),
            .I(N__5623));
    InMux I__842 (
            .O(N__5635),
            .I(N__5616));
    InMux I__841 (
            .O(N__5634),
            .I(N__5616));
    InMux I__840 (
            .O(N__5633),
            .I(N__5616));
    InMux I__839 (
            .O(N__5630),
            .I(N__5613));
    LocalMux I__838 (
            .O(N__5623),
            .I(N__5610));
    LocalMux I__837 (
            .O(N__5616),
            .I(\U409_AUTOCONFIG.un1_STATE_6Z0Z_0 ));
    LocalMux I__836 (
            .O(N__5613),
            .I(\U409_AUTOCONFIG.un1_STATE_6Z0Z_0 ));
    Odrv4 I__835 (
            .O(N__5610),
            .I(\U409_AUTOCONFIG.un1_STATE_6Z0Z_0 ));
    InMux I__834 (
            .O(N__5603),
            .I(N__5597));
    InMux I__833 (
            .O(N__5602),
            .I(N__5597));
    LocalMux I__832 (
            .O(N__5597),
            .I(LIDE_BASE_6));
    CascadeMux I__831 (
            .O(N__5594),
            .I(N__5591));
    InMux I__830 (
            .O(N__5591),
            .I(N__5588));
    LocalMux I__829 (
            .O(N__5588),
            .I(N__5585));
    Odrv12 I__828 (
            .O(N__5585),
            .I(\U409_AUTOCONFIG.PR_OUTZ0Z_3 ));
    InMux I__827 (
            .O(N__5582),
            .I(N__5579));
    LocalMux I__826 (
            .O(N__5579),
            .I(N__5576));
    Odrv4 I__825 (
            .O(N__5576),
            .I(\U409_AUTOCONFIG.PR_OUT_cnst_i_0_2 ));
    InMux I__824 (
            .O(N__5573),
            .I(N__5570));
    LocalMux I__823 (
            .O(N__5570),
            .I(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ));
    InMux I__822 (
            .O(N__5567),
            .I(N__5564));
    LocalMux I__821 (
            .O(N__5564),
            .I(N__5561));
    Odrv12 I__820 (
            .O(N__5561),
            .I(\U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3 ));
    InMux I__819 (
            .O(N__5558),
            .I(N__5551));
    InMux I__818 (
            .O(N__5557),
            .I(N__5551));
    InMux I__817 (
            .O(N__5556),
            .I(N__5548));
    LocalMux I__816 (
            .O(N__5551),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_5 ));
    LocalMux I__815 (
            .O(N__5548),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_5 ));
    CascadeMux I__814 (
            .O(N__5543),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_4_cascade_ ));
    InMux I__813 (
            .O(N__5540),
            .I(N__5537));
    LocalMux I__812 (
            .O(N__5537),
            .I(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_1 ));
    IoInMux I__811 (
            .O(N__5534),
            .I(N__5531));
    LocalMux I__810 (
            .O(N__5531),
            .I(N__5528));
    IoSpan4Mux I__809 (
            .O(N__5528),
            .I(N__5525));
    Span4Mux_s1_v I__808 (
            .O(N__5525),
            .I(N__5522));
    Span4Mux_h I__807 (
            .O(N__5522),
            .I(N__5519));
    Sp12to4 I__806 (
            .O(N__5519),
            .I(N__5516));
    Span12Mux_v I__805 (
            .O(N__5516),
            .I(N__5513));
    Odrv12 I__804 (
            .O(N__5513),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn_i));
    IoInMux I__803 (
            .O(N__5510),
            .I(N__5507));
    LocalMux I__802 (
            .O(N__5507),
            .I(N__5502));
    IoInMux I__801 (
            .O(N__5506),
            .I(N__5499));
    IoInMux I__800 (
            .O(N__5505),
            .I(N__5496));
    IoSpan4Mux I__799 (
            .O(N__5502),
            .I(N__5493));
    LocalMux I__798 (
            .O(N__5499),
            .I(N__5488));
    LocalMux I__797 (
            .O(N__5496),
            .I(N__5488));
    Span4Mux_s3_v I__796 (
            .O(N__5493),
            .I(N__5482));
    Span4Mux_s3_v I__795 (
            .O(N__5488),
            .I(N__5482));
    IoInMux I__794 (
            .O(N__5487),
            .I(N__5479));
    Span4Mux_v I__793 (
            .O(N__5482),
            .I(N__5476));
    LocalMux I__792 (
            .O(N__5479),
            .I(N__5473));
    Odrv4 I__791 (
            .O(N__5476),
            .I(D_1_i));
    Odrv12 I__790 (
            .O(N__5473),
            .I(D_1_i));
    InMux I__789 (
            .O(N__5468),
            .I(N__5465));
    LocalMux I__788 (
            .O(N__5465),
            .I(N__5462));
    Odrv12 I__787 (
            .O(N__5462),
            .I(D_in_4));
    InMux I__786 (
            .O(N__5459),
            .I(N__5456));
    LocalMux I__785 (
            .O(N__5456),
            .I(\U409_AUTOCONFIG.N_76 ));
    InMux I__784 (
            .O(N__5453),
            .I(N__5447));
    InMux I__783 (
            .O(N__5452),
            .I(N__5447));
    LocalMux I__782 (
            .O(N__5447),
            .I(N__5444));
    Sp12to4 I__781 (
            .O(N__5444),
            .I(N__5441));
    Span12Mux_v I__780 (
            .O(N__5441),
            .I(N__5438));
    Odrv12 I__779 (
            .O(N__5438),
            .I(D_in_6));
    InMux I__778 (
            .O(N__5435),
            .I(N__5429));
    InMux I__777 (
            .O(N__5434),
            .I(N__5429));
    LocalMux I__776 (
            .O(N__5429),
            .I(N__5426));
    Span4Mux_v I__775 (
            .O(N__5426),
            .I(N__5423));
    Span4Mux_v I__774 (
            .O(N__5423),
            .I(N__5420));
    Odrv4 I__773 (
            .O(N__5420),
            .I(D_in_5));
    InMux I__772 (
            .O(N__5417),
            .I(N__5414));
    LocalMux I__771 (
            .O(N__5414),
            .I(\U409_AUTOCONFIG.N_82 ));
    IoInMux I__770 (
            .O(N__5411),
            .I(N__5408));
    LocalMux I__769 (
            .O(N__5408),
            .I(N__5405));
    Span4Mux_s3_v I__768 (
            .O(N__5405),
            .I(N__5402));
    Span4Mux_v I__767 (
            .O(N__5402),
            .I(N__5399));
    Span4Mux_h I__766 (
            .O(N__5399),
            .I(N__5396));
    Odrv4 I__765 (
            .O(N__5396),
            .I(D_OUT_3));
    InMux I__764 (
            .O(N__5393),
            .I(N__5390));
    LocalMux I__763 (
            .O(N__5390),
            .I(\U409_AUTOCONFIG.N_80 ));
    CascadeMux I__762 (
            .O(N__5387),
            .I(N__5384));
    InMux I__761 (
            .O(N__5384),
            .I(N__5380));
    InMux I__760 (
            .O(N__5383),
            .I(N__5377));
    LocalMux I__759 (
            .O(N__5380),
            .I(LIDE_BASE_2));
    LocalMux I__758 (
            .O(N__5377),
            .I(LIDE_BASE_2));
    InMux I__757 (
            .O(N__5372),
            .I(N__5368));
    InMux I__756 (
            .O(N__5371),
            .I(N__5365));
    LocalMux I__755 (
            .O(N__5368),
            .I(\U409_ADDRESS_DECODE.N_34_1 ));
    LocalMux I__754 (
            .O(N__5365),
            .I(\U409_ADDRESS_DECODE.N_34_1 ));
    CascadeMux I__753 (
            .O(N__5360),
            .I(N__5357));
    InMux I__752 (
            .O(N__5357),
            .I(N__5354));
    LocalMux I__751 (
            .O(N__5354),
            .I(\U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0Z0Z_0 ));
    InMux I__750 (
            .O(N__5351),
            .I(N__5347));
    InMux I__749 (
            .O(N__5350),
            .I(N__5344));
    LocalMux I__748 (
            .O(N__5347),
            .I(N__5341));
    LocalMux I__747 (
            .O(N__5344),
            .I(N__5338));
    Span4Mux_v I__746 (
            .O(N__5341),
            .I(N__5333));
    Span4Mux_h I__745 (
            .O(N__5338),
            .I(N__5333));
    Odrv4 I__744 (
            .O(N__5333),
            .I(N_100));
    InMux I__743 (
            .O(N__5330),
            .I(N__5327));
    LocalMux I__742 (
            .O(N__5327),
            .I(N__5323));
    InMux I__741 (
            .O(N__5326),
            .I(N__5320));
    Span12Mux_h I__740 (
            .O(N__5323),
            .I(N__5314));
    LocalMux I__739 (
            .O(N__5320),
            .I(N__5314));
    InMux I__738 (
            .O(N__5319),
            .I(N__5311));
    Odrv12 I__737 (
            .O(N__5314),
            .I(N_94));
    LocalMux I__736 (
            .O(N__5311),
            .I(N_94));
    CascadeMux I__735 (
            .O(N__5306),
            .I(\U409_AUTOCONFIG.PORTSIZEZ0Z_1_cascade_ ));
    IoInMux I__734 (
            .O(N__5303),
            .I(N__5300));
    LocalMux I__733 (
            .O(N__5300),
            .I(N__5297));
    Span4Mux_s3_v I__732 (
            .O(N__5297),
            .I(N__5294));
    Span4Mux_v I__731 (
            .O(N__5294),
            .I(N__5291));
    Span4Mux_v I__730 (
            .O(N__5291),
            .I(N__5288));
    Span4Mux_v I__729 (
            .O(N__5288),
            .I(N__5285));
    Odrv4 I__728 (
            .O(N__5285),
            .I(PORTSIZE_0_i));
    InMux I__727 (
            .O(N__5282),
            .I(N__5279));
    LocalMux I__726 (
            .O(N__5279),
            .I(N__5276));
    Odrv12 I__725 (
            .O(N__5276),
            .I(\U409_AUTOCONFIG.un1_STATE_6_0_0 ));
    InMux I__724 (
            .O(N__5273),
            .I(N__5266));
    InMux I__723 (
            .O(N__5272),
            .I(N__5257));
    InMux I__722 (
            .O(N__5271),
            .I(N__5257));
    InMux I__721 (
            .O(N__5270),
            .I(N__5257));
    InMux I__720 (
            .O(N__5269),
            .I(N__5257));
    LocalMux I__719 (
            .O(N__5266),
            .I(N__5254));
    LocalMux I__718 (
            .O(N__5257),
            .I(N__5251));
    Span4Mux_h I__717 (
            .O(N__5254),
            .I(N__5247));
    Span4Mux_v I__716 (
            .O(N__5251),
            .I(N__5244));
    InMux I__715 (
            .O(N__5250),
            .I(N__5241));
    Span4Mux_v I__714 (
            .O(N__5247),
            .I(N__5238));
    Sp12to4 I__713 (
            .O(N__5244),
            .I(N__5233));
    LocalMux I__712 (
            .O(N__5241),
            .I(N__5233));
    Sp12to4 I__711 (
            .O(N__5238),
            .I(N__5228));
    Span12Mux_h I__710 (
            .O(N__5233),
            .I(N__5228));
    Odrv12 I__709 (
            .O(N__5228),
            .I(A_c_5));
    InMux I__708 (
            .O(N__5225),
            .I(N__5221));
    InMux I__707 (
            .O(N__5224),
            .I(N__5217));
    LocalMux I__706 (
            .O(N__5221),
            .I(N__5214));
    InMux I__705 (
            .O(N__5220),
            .I(N__5211));
    LocalMux I__704 (
            .O(N__5217),
            .I(N__5206));
    Span4Mux_h I__703 (
            .O(N__5214),
            .I(N__5200));
    LocalMux I__702 (
            .O(N__5211),
            .I(N__5200));
    InMux I__701 (
            .O(N__5210),
            .I(N__5197));
    InMux I__700 (
            .O(N__5209),
            .I(N__5194));
    Span4Mux_v I__699 (
            .O(N__5206),
            .I(N__5191));
    InMux I__698 (
            .O(N__5205),
            .I(N__5188));
    Span4Mux_v I__697 (
            .O(N__5200),
            .I(N__5179));
    LocalMux I__696 (
            .O(N__5197),
            .I(N__5179));
    LocalMux I__695 (
            .O(N__5194),
            .I(N__5179));
    Span4Mux_v I__694 (
            .O(N__5191),
            .I(N__5176));
    LocalMux I__693 (
            .O(N__5188),
            .I(N__5173));
    InMux I__692 (
            .O(N__5187),
            .I(N__5170));
    InMux I__691 (
            .O(N__5186),
            .I(N__5167));
    Span4Mux_v I__690 (
            .O(N__5179),
            .I(N__5164));
    Span4Mux_v I__689 (
            .O(N__5176),
            .I(N__5157));
    Span4Mux_v I__688 (
            .O(N__5173),
            .I(N__5157));
    LocalMux I__687 (
            .O(N__5170),
            .I(N__5157));
    LocalMux I__686 (
            .O(N__5167),
            .I(N__5154));
    Sp12to4 I__685 (
            .O(N__5164),
            .I(N__5149));
    Sp12to4 I__684 (
            .O(N__5157),
            .I(N__5149));
    Span12Mux_v I__683 (
            .O(N__5154),
            .I(N__5146));
    Odrv12 I__682 (
            .O(N__5149),
            .I(A_c_20));
    Odrv12 I__681 (
            .O(N__5146),
            .I(A_c_20));
    CascadeMux I__680 (
            .O(N__5141),
            .I(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_1_cascade_ ));
    InMux I__679 (
            .O(N__5138),
            .I(N__5132));
    CascadeMux I__678 (
            .O(N__5137),
            .I(N__5129));
    CascadeMux I__677 (
            .O(N__5136),
            .I(N__5124));
    CascadeMux I__676 (
            .O(N__5135),
            .I(N__5121));
    LocalMux I__675 (
            .O(N__5132),
            .I(N__5118));
    InMux I__674 (
            .O(N__5129),
            .I(N__5115));
    InMux I__673 (
            .O(N__5128),
            .I(N__5110));
    InMux I__672 (
            .O(N__5127),
            .I(N__5110));
    InMux I__671 (
            .O(N__5124),
            .I(N__5107));
    InMux I__670 (
            .O(N__5121),
            .I(N__5103));
    Span4Mux_v I__669 (
            .O(N__5118),
            .I(N__5094));
    LocalMux I__668 (
            .O(N__5115),
            .I(N__5094));
    LocalMux I__667 (
            .O(N__5110),
            .I(N__5094));
    LocalMux I__666 (
            .O(N__5107),
            .I(N__5094));
    InMux I__665 (
            .O(N__5106),
            .I(N__5091));
    LocalMux I__664 (
            .O(N__5103),
            .I(N__5088));
    Span4Mux_v I__663 (
            .O(N__5094),
            .I(N__5083));
    LocalMux I__662 (
            .O(N__5091),
            .I(N__5083));
    Span4Mux_v I__661 (
            .O(N__5088),
            .I(N__5080));
    Span4Mux_v I__660 (
            .O(N__5083),
            .I(N__5077));
    Sp12to4 I__659 (
            .O(N__5080),
            .I(N__5072));
    Sp12to4 I__658 (
            .O(N__5077),
            .I(N__5072));
    Odrv12 I__657 (
            .O(N__5072),
            .I(A_c_23));
    InMux I__656 (
            .O(N__5069),
            .I(N__5063));
    InMux I__655 (
            .O(N__5068),
            .I(N__5063));
    LocalMux I__654 (
            .O(N__5063),
            .I(N__5058));
    InMux I__653 (
            .O(N__5062),
            .I(N__5055));
    InMux I__652 (
            .O(N__5061),
            .I(N__5052));
    Span4Mux_v I__651 (
            .O(N__5058),
            .I(N__5047));
    LocalMux I__650 (
            .O(N__5055),
            .I(N__5047));
    LocalMux I__649 (
            .O(N__5052),
            .I(N__5044));
    Span4Mux_h I__648 (
            .O(N__5047),
            .I(N__5041));
    Span12Mux_v I__647 (
            .O(N__5044),
            .I(N__5038));
    Odrv4 I__646 (
            .O(N__5041),
            .I(\U409_ADDRESS_DECODE.N_92 ));
    Odrv12 I__645 (
            .O(N__5038),
            .I(\U409_ADDRESS_DECODE.N_92 ));
    InMux I__644 (
            .O(N__5033),
            .I(N__5030));
    LocalMux I__643 (
            .O(N__5030),
            .I(N__5026));
    InMux I__642 (
            .O(N__5029),
            .I(N__5023));
    Odrv4 I__641 (
            .O(N__5026),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_4 ));
    LocalMux I__640 (
            .O(N__5023),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_4 ));
    InMux I__639 (
            .O(N__5018),
            .I(N__5015));
    LocalMux I__638 (
            .O(N__5015),
            .I(N__5012));
    Odrv4 I__637 (
            .O(N__5012),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE ));
    InMux I__636 (
            .O(N__5009),
            .I(N__5006));
    LocalMux I__635 (
            .O(N__5006),
            .I(\U409_ADDRESS_DECODE.N_34 ));
    InMux I__634 (
            .O(N__5003),
            .I(N__5000));
    LocalMux I__633 (
            .O(N__5000),
            .I(\U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_3 ));
    CascadeMux I__632 (
            .O(N__4997),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE_cascade_ ));
    InMux I__631 (
            .O(N__4994),
            .I(N__4991));
    LocalMux I__630 (
            .O(N__4991),
            .I(\U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_2 ));
    CascadeMux I__629 (
            .O(N__4988),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_0Z0Z_2_cascade_ ));
    InMux I__628 (
            .O(N__4985),
            .I(N__4982));
    LocalMux I__627 (
            .O(N__4982),
            .I(N__4979));
    Odrv4 I__626 (
            .O(N__4979),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_4 ));
    CascadeMux I__625 (
            .O(N__4976),
            .I(N__4972));
    InMux I__624 (
            .O(N__4975),
            .I(N__4967));
    InMux I__623 (
            .O(N__4972),
            .I(N__4967));
    LocalMux I__622 (
            .O(N__4967),
            .I(\U409_AUTOCONFIG.N_227_3 ));
    CascadeMux I__621 (
            .O(N__4964),
            .I(\U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_4_cascade_ ));
    InMux I__620 (
            .O(N__4961),
            .I(N__4958));
    LocalMux I__619 (
            .O(N__4958),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4 ));
    CascadeMux I__618 (
            .O(N__4955),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2_cascade_ ));
    InMux I__617 (
            .O(N__4952),
            .I(N__4949));
    LocalMux I__616 (
            .O(N__4949),
            .I(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1 ));
    CascadeMux I__615 (
            .O(N__4946),
            .I(ATA_SPACE_cascade_));
    InMux I__614 (
            .O(N__4943),
            .I(N__4939));
    InMux I__613 (
            .O(N__4942),
            .I(N__4936));
    LocalMux I__612 (
            .O(N__4939),
            .I(\U409_ADDRESS_DECODE.ATA_ENZ0 ));
    LocalMux I__611 (
            .O(N__4936),
            .I(\U409_ADDRESS_DECODE.ATA_ENZ0 ));
    InMux I__610 (
            .O(N__4931),
            .I(N__4928));
    LocalMux I__609 (
            .O(N__4928),
            .I(N__4924));
    InMux I__608 (
            .O(N__4927),
            .I(N__4921));
    Odrv12 I__607 (
            .O(N__4924),
            .I(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1 ));
    LocalMux I__606 (
            .O(N__4921),
            .I(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1 ));
    InMux I__605 (
            .O(N__4916),
            .I(N__4913));
    LocalMux I__604 (
            .O(N__4913),
            .I(N__4908));
    InMux I__603 (
            .O(N__4912),
            .I(N__4905));
    InMux I__602 (
            .O(N__4911),
            .I(N__4902));
    Span4Mux_v I__601 (
            .O(N__4908),
            .I(N__4895));
    LocalMux I__600 (
            .O(N__4905),
            .I(N__4895));
    LocalMux I__599 (
            .O(N__4902),
            .I(N__4895));
    Span4Mux_v I__598 (
            .O(N__4895),
            .I(N__4892));
    Span4Mux_v I__597 (
            .O(N__4892),
            .I(N__4889));
    Sp12to4 I__596 (
            .O(N__4889),
            .I(N__4886));
    Span12Mux_h I__595 (
            .O(N__4886),
            .I(N__4883));
    Odrv12 I__594 (
            .O(N__4883),
            .I(OVL_c));
    InMux I__593 (
            .O(N__4880),
            .I(N__4874));
    InMux I__592 (
            .O(N__4879),
            .I(N__4874));
    LocalMux I__591 (
            .O(N__4874),
            .I(N__4869));
    InMux I__590 (
            .O(N__4873),
            .I(N__4864));
    InMux I__589 (
            .O(N__4872),
            .I(N__4864));
    Span4Mux_h I__588 (
            .O(N__4869),
            .I(N__4858));
    LocalMux I__587 (
            .O(N__4864),
            .I(N__4858));
    CascadeMux I__586 (
            .O(N__4863),
            .I(N__4855));
    Span4Mux_v I__585 (
            .O(N__4858),
            .I(N__4852));
    InMux I__584 (
            .O(N__4855),
            .I(N__4849));
    Sp12to4 I__583 (
            .O(N__4852),
            .I(N__4844));
    LocalMux I__582 (
            .O(N__4849),
            .I(N__4844));
    Span12Mux_h I__581 (
            .O(N__4844),
            .I(N__4841));
    Span12Mux_v I__580 (
            .O(N__4841),
            .I(N__4838));
    Odrv12 I__579 (
            .O(N__4838),
            .I(A_c_19));
    CascadeMux I__578 (
            .O(N__4835),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_1_cascade_ ));
    InMux I__577 (
            .O(N__4832),
            .I(N__4829));
    LocalMux I__576 (
            .O(N__4829),
            .I(N__4824));
    CascadeMux I__575 (
            .O(N__4828),
            .I(N__4821));
    InMux I__574 (
            .O(N__4827),
            .I(N__4818));
    Span4Mux_v I__573 (
            .O(N__4824),
            .I(N__4813));
    InMux I__572 (
            .O(N__4821),
            .I(N__4810));
    LocalMux I__571 (
            .O(N__4818),
            .I(N__4807));
    InMux I__570 (
            .O(N__4817),
            .I(N__4802));
    InMux I__569 (
            .O(N__4816),
            .I(N__4802));
    Sp12to4 I__568 (
            .O(N__4813),
            .I(N__4799));
    LocalMux I__567 (
            .O(N__4810),
            .I(N__4796));
    Span4Mux_v I__566 (
            .O(N__4807),
            .I(N__4791));
    LocalMux I__565 (
            .O(N__4802),
            .I(N__4791));
    Span12Mux_s7_h I__564 (
            .O(N__4799),
            .I(N__4786));
    Span12Mux_h I__563 (
            .O(N__4796),
            .I(N__4786));
    Span4Mux_v I__562 (
            .O(N__4791),
            .I(N__4783));
    Span12Mux_v I__561 (
            .O(N__4786),
            .I(N__4780));
    Sp12to4 I__560 (
            .O(N__4783),
            .I(N__4777));
    Odrv12 I__559 (
            .O(N__4780),
            .I(A_c_16));
    Odrv12 I__558 (
            .O(N__4777),
            .I(A_c_16));
    IoInMux I__557 (
            .O(N__4772),
            .I(N__4769));
    LocalMux I__556 (
            .O(N__4769),
            .I(N__4766));
    IoSpan4Mux I__555 (
            .O(N__4766),
            .I(N__4763));
    Span4Mux_s2_v I__554 (
            .O(N__4763),
            .I(N__4760));
    Span4Mux_v I__553 (
            .O(N__4760),
            .I(N__4757));
    Span4Mux_v I__552 (
            .O(N__4757),
            .I(N__4754));
    Odrv4 I__551 (
            .O(N__4754),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn_i));
    InMux I__550 (
            .O(N__4751),
            .I(N__4744));
    InMux I__549 (
            .O(N__4750),
            .I(N__4744));
    InMux I__548 (
            .O(N__4749),
            .I(N__4741));
    LocalMux I__547 (
            .O(N__4744),
            .I(N__4735));
    LocalMux I__546 (
            .O(N__4741),
            .I(N__4732));
    InMux I__545 (
            .O(N__4740),
            .I(N__4729));
    InMux I__544 (
            .O(N__4739),
            .I(N__4726));
    InMux I__543 (
            .O(N__4738),
            .I(N__4723));
    Span4Mux_v I__542 (
            .O(N__4735),
            .I(N__4720));
    Span4Mux_v I__541 (
            .O(N__4732),
            .I(N__4717));
    LocalMux I__540 (
            .O(N__4729),
            .I(N__4714));
    LocalMux I__539 (
            .O(N__4726),
            .I(N__4709));
    LocalMux I__538 (
            .O(N__4723),
            .I(N__4709));
    Sp12to4 I__537 (
            .O(N__4720),
            .I(N__4704));
    Sp12to4 I__536 (
            .O(N__4717),
            .I(N__4704));
    Span4Mux_v I__535 (
            .O(N__4714),
            .I(N__4701));
    Span4Mux_v I__534 (
            .O(N__4709),
            .I(N__4698));
    Span12Mux_s11_h I__533 (
            .O(N__4704),
            .I(N__4695));
    Span4Mux_v I__532 (
            .O(N__4701),
            .I(N__4692));
    Span4Mux_v I__531 (
            .O(N__4698),
            .I(N__4689));
    Span12Mux_v I__530 (
            .O(N__4695),
            .I(N__4682));
    Sp12to4 I__529 (
            .O(N__4692),
            .I(N__4682));
    Sp12to4 I__528 (
            .O(N__4689),
            .I(N__4682));
    Odrv12 I__527 (
            .O(N__4682),
            .I(A_c_18));
    InMux I__526 (
            .O(N__4679),
            .I(N__4672));
    InMux I__525 (
            .O(N__4678),
            .I(N__4672));
    InMux I__524 (
            .O(N__4677),
            .I(N__4668));
    LocalMux I__523 (
            .O(N__4672),
            .I(N__4665));
    CascadeMux I__522 (
            .O(N__4671),
            .I(N__4662));
    LocalMux I__521 (
            .O(N__4668),
            .I(N__4659));
    Span4Mux_v I__520 (
            .O(N__4665),
            .I(N__4656));
    InMux I__519 (
            .O(N__4662),
            .I(N__4653));
    Span12Mux_v I__518 (
            .O(N__4659),
            .I(N__4650));
    Sp12to4 I__517 (
            .O(N__4656),
            .I(N__4645));
    LocalMux I__516 (
            .O(N__4653),
            .I(N__4645));
    Span12Mux_v I__515 (
            .O(N__4650),
            .I(N__4642));
    Span12Mux_v I__514 (
            .O(N__4645),
            .I(N__4639));
    Odrv12 I__513 (
            .O(N__4642),
            .I(A_c_17));
    Odrv12 I__512 (
            .O(N__4639),
            .I(A_c_17));
    InMux I__511 (
            .O(N__4634),
            .I(N__4628));
    InMux I__510 (
            .O(N__4633),
            .I(N__4628));
    LocalMux I__509 (
            .O(N__4628),
            .I(LIDE_BASE_1));
    InMux I__508 (
            .O(N__4625),
            .I(N__4621));
    InMux I__507 (
            .O(N__4624),
            .I(N__4618));
    LocalMux I__506 (
            .O(N__4621),
            .I(LIDE_BASE_4));
    LocalMux I__505 (
            .O(N__4618),
            .I(LIDE_BASE_4));
    InMux I__504 (
            .O(N__4613),
            .I(N__4609));
    InMux I__503 (
            .O(N__4612),
            .I(N__4606));
    LocalMux I__502 (
            .O(N__4609),
            .I(LIDE_BASE_3));
    LocalMux I__501 (
            .O(N__4606),
            .I(LIDE_BASE_3));
    CascadeMux I__500 (
            .O(N__4601),
            .I(N_89_cascade_));
    CascadeMux I__499 (
            .O(N__4598),
            .I(N_94_cascade_));
    InMux I__498 (
            .O(N__4595),
            .I(N__4592));
    LocalMux I__497 (
            .O(N__4592),
            .I(N__4589));
    Span4Mux_v I__496 (
            .O(N__4589),
            .I(N__4586));
    Odrv4 I__495 (
            .O(N__4586),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3Z0Z_1 ));
    InMux I__494 (
            .O(N__4583),
            .I(N__4580));
    LocalMux I__493 (
            .O(N__4580),
            .I(N__4577));
    Span4Mux_v I__492 (
            .O(N__4577),
            .I(N__4574));
    Span4Mux_h I__491 (
            .O(N__4574),
            .I(N__4571));
    Sp12to4 I__490 (
            .O(N__4571),
            .I(N__4568));
    Odrv12 I__489 (
            .O(N__4568),
            .I(TT_c_0));
    InMux I__488 (
            .O(N__4565),
            .I(N__4562));
    LocalMux I__487 (
            .O(N__4562),
            .I(N__4559));
    Span4Mux_v I__486 (
            .O(N__4559),
            .I(N__4556));
    Span4Mux_h I__485 (
            .O(N__4556),
            .I(N__4553));
    Sp12to4 I__484 (
            .O(N__4553),
            .I(N__4550));
    Odrv12 I__483 (
            .O(N__4550),
            .I(TT_c_1));
    CascadeMux I__482 (
            .O(N__4547),
            .I(N__4544));
    InMux I__481 (
            .O(N__4544),
            .I(N__4541));
    LocalMux I__480 (
            .O(N__4541),
            .I(N__4538));
    Odrv4 I__479 (
            .O(N__4538),
            .I(N_89));
    InMux I__478 (
            .O(N__4535),
            .I(N__4532));
    LocalMux I__477 (
            .O(N__4532),
            .I(N__4529));
    Odrv12 I__476 (
            .O(N__4529),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_8 ));
    CascadeMux I__475 (
            .O(N__4526),
            .I(N__4522));
    InMux I__474 (
            .O(N__4525),
            .I(N__4517));
    InMux I__473 (
            .O(N__4522),
            .I(N__4517));
    LocalMux I__472 (
            .O(N__4517),
            .I(N__4514));
    Span12Mux_v I__471 (
            .O(N__4514),
            .I(N__4511));
    Odrv12 I__470 (
            .O(N__4511),
            .I(A_c_15));
    CascadeMux I__469 (
            .O(N__4508),
            .I(N__4505));
    InMux I__468 (
            .O(N__4505),
            .I(N__4499));
    InMux I__467 (
            .O(N__4504),
            .I(N__4499));
    LocalMux I__466 (
            .O(N__4499),
            .I(N__4496));
    Span4Mux_v I__465 (
            .O(N__4496),
            .I(N__4493));
    Span4Mux_h I__464 (
            .O(N__4493),
            .I(N__4490));
    Odrv4 I__463 (
            .O(N__4490),
            .I(A_c_25));
    CascadeMux I__462 (
            .O(N__4487),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_3_cascade_ ));
    InMux I__461 (
            .O(N__4484),
            .I(N__4478));
    InMux I__460 (
            .O(N__4483),
            .I(N__4478));
    LocalMux I__459 (
            .O(N__4478),
            .I(N__4475));
    Span4Mux_v I__458 (
            .O(N__4475),
            .I(N__4472));
    Span4Mux_v I__457 (
            .O(N__4472),
            .I(N__4469));
    Sp12to4 I__456 (
            .O(N__4469),
            .I(N__4466));
    Odrv12 I__455 (
            .O(N__4466),
            .I(A_c_24));
    InMux I__454 (
            .O(N__4463),
            .I(N__4460));
    LocalMux I__453 (
            .O(N__4460),
            .I(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4 ));
    InMux I__452 (
            .O(N__4457),
            .I(N__4454));
    LocalMux I__451 (
            .O(N__4454),
            .I(N__4451));
    Span4Mux_v I__450 (
            .O(N__4451),
            .I(N__4447));
    InMux I__449 (
            .O(N__4450),
            .I(N__4444));
    Sp12to4 I__448 (
            .O(N__4447),
            .I(N__4439));
    LocalMux I__447 (
            .O(N__4444),
            .I(N__4439));
    Odrv12 I__446 (
            .O(N__4439),
            .I(A_c_27));
    InMux I__445 (
            .O(N__4436),
            .I(N__4430));
    InMux I__444 (
            .O(N__4435),
            .I(N__4430));
    LocalMux I__443 (
            .O(N__4430),
            .I(N__4427));
    Span4Mux_v I__442 (
            .O(N__4427),
            .I(N__4424));
    Sp12to4 I__441 (
            .O(N__4424),
            .I(N__4421));
    Odrv12 I__440 (
            .O(N__4421),
            .I(A_c_30));
    CascadeMux I__439 (
            .O(N__4418),
            .I(N__4415));
    InMux I__438 (
            .O(N__4415),
            .I(N__4409));
    InMux I__437 (
            .O(N__4414),
            .I(N__4409));
    LocalMux I__436 (
            .O(N__4409),
            .I(N__4406));
    Span4Mux_h I__435 (
            .O(N__4406),
            .I(N__4403));
    Span4Mux_v I__434 (
            .O(N__4403),
            .I(N__4400));
    Span4Mux_v I__433 (
            .O(N__4400),
            .I(N__4397));
    Odrv4 I__432 (
            .O(N__4397),
            .I(A_c_28));
    CascadeMux I__431 (
            .O(N__4394),
            .I(N__4390));
    InMux I__430 (
            .O(N__4393),
            .I(N__4385));
    InMux I__429 (
            .O(N__4390),
            .I(N__4385));
    LocalMux I__428 (
            .O(N__4385),
            .I(N__4382));
    Sp12to4 I__427 (
            .O(N__4382),
            .I(N__4379));
    Span12Mux_v I__426 (
            .O(N__4379),
            .I(N__4376));
    Odrv12 I__425 (
            .O(N__4376),
            .I(A_c_29));
    InMux I__424 (
            .O(N__4373),
            .I(N__4370));
    LocalMux I__423 (
            .O(N__4370),
            .I(N__4367));
    Span4Mux_v I__422 (
            .O(N__4367),
            .I(N__4363));
    InMux I__421 (
            .O(N__4366),
            .I(N__4360));
    Span4Mux_v I__420 (
            .O(N__4363),
            .I(N__4357));
    LocalMux I__419 (
            .O(N__4360),
            .I(N__4354));
    Sp12to4 I__418 (
            .O(N__4357),
            .I(N__4351));
    Span4Mux_v I__417 (
            .O(N__4354),
            .I(N__4348));
    Span12Mux_h I__416 (
            .O(N__4351),
            .I(N__4343));
    Sp12to4 I__415 (
            .O(N__4348),
            .I(N__4343));
    Odrv12 I__414 (
            .O(N__4343),
            .I(A_c_31));
    InMux I__413 (
            .O(N__4340),
            .I(N__4337));
    LocalMux I__412 (
            .O(N__4337),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_9 ));
    CascadeMux I__411 (
            .O(N__4334),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_11_cascade_ ));
    InMux I__410 (
            .O(N__4331),
            .I(N__4328));
    LocalMux I__409 (
            .O(N__4328),
            .I(N__4325));
    Odrv4 I__408 (
            .O(N__4325),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_10 ));
    IoInMux I__407 (
            .O(N__4322),
            .I(N__4319));
    LocalMux I__406 (
            .O(N__4319),
            .I(N__4316));
    Span12Mux_s11_h I__405 (
            .O(N__4316),
            .I(N__4313));
    Span12Mux_h I__404 (
            .O(N__4313),
            .I(N__4310));
    Odrv12 I__403 (
            .O(N__4310),
            .I(N_61_i));
    IoInMux I__402 (
            .O(N__4307),
            .I(N__4304));
    LocalMux I__401 (
            .O(N__4304),
            .I(N__4301));
    Span12Mux_s2_h I__400 (
            .O(N__4301),
            .I(N__4298));
    Span12Mux_v I__399 (
            .O(N__4298),
            .I(N__4295));
    Odrv12 I__398 (
            .O(N__4295),
            .I(SPIO_c));
    InMux I__397 (
            .O(N__4292),
            .I(N__4286));
    InMux I__396 (
            .O(N__4291),
            .I(N__4286));
    LocalMux I__395 (
            .O(N__4286),
            .I(N__4283));
    Span4Mux_v I__394 (
            .O(N__4283),
            .I(N__4280));
    Span4Mux_v I__393 (
            .O(N__4280),
            .I(N__4277));
    Sp12to4 I__392 (
            .O(N__4277),
            .I(N__4274));
    Odrv12 I__391 (
            .O(N__4274),
            .I(A_c_26));
    IoInMux I__390 (
            .O(N__4271),
            .I(N__4268));
    LocalMux I__389 (
            .O(N__4268),
            .I(N__4265));
    IoSpan4Mux I__388 (
            .O(N__4265),
            .I(N__4262));
    Sp12to4 I__387 (
            .O(N__4262),
            .I(N__4259));
    Span12Mux_s1_h I__386 (
            .O(N__4259),
            .I(N__4256));
    Span12Mux_v I__385 (
            .O(N__4256),
            .I(N__4253));
    Odrv12 I__384 (
            .O(N__4253),
            .I(PPIO_c));
    ClkMux I__383 (
            .O(N__4250),
            .I(N__4211));
    ClkMux I__382 (
            .O(N__4249),
            .I(N__4211));
    ClkMux I__381 (
            .O(N__4248),
            .I(N__4211));
    ClkMux I__380 (
            .O(N__4247),
            .I(N__4211));
    ClkMux I__379 (
            .O(N__4246),
            .I(N__4211));
    ClkMux I__378 (
            .O(N__4245),
            .I(N__4211));
    ClkMux I__377 (
            .O(N__4244),
            .I(N__4211));
    ClkMux I__376 (
            .O(N__4243),
            .I(N__4211));
    ClkMux I__375 (
            .O(N__4242),
            .I(N__4211));
    ClkMux I__374 (
            .O(N__4241),
            .I(N__4211));
    ClkMux I__373 (
            .O(N__4240),
            .I(N__4211));
    ClkMux I__372 (
            .O(N__4239),
            .I(N__4211));
    ClkMux I__371 (
            .O(N__4238),
            .I(N__4211));
    GlobalMux I__370 (
            .O(N__4211),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.LASTCLK_1C  (
            .O(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .I(N__4250));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ),
            .I(N__4249));
    INV \INVU409_TRANSFER_ACK.CIA_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .I(N__4246));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_0C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .I(N__4243));
    INV \INVU409_TRANSFER_ACK.ROMENnC  (
            .O(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .I(N__4248));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .I(N__4242));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .I(N__4240));
    INV \INVU409_TRANSFER_ACK.TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .I(N__4239));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .I(N__4238));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .I(N__4245));
    INV \INVU409_TRANSFER_ACK.TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .I(N__4241));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .I(N__4247));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .I(N__4244));
    INV \INVU409_AUTOCONFIG.AC_TACKC  (
            .O(\INVU409_AUTOCONFIG.AC_TACKC_net ),
            .I(N__9889));
    INV \INVU409_AUTOCONFIG.STATE_0C  (
            .O(\INVU409_AUTOCONFIG.STATE_0C_net ),
            .I(N__9891));
    INV \INVU409_AUTOCONFIG.CONFIGENnC  (
            .O(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .I(N__9898));
    INV \INVU409_AUTOCONFIG.LIDE_OUT_1C  (
            .O(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .I(N__9896));
    INV \INVU409_AUTOCONFIG.LIDE_OUT_3C  (
            .O(\INVU409_AUTOCONFIG.LIDE_OUT_3C_net ),
            .I(N__9895));
    INV \INVU409_AUTOCONFIG.PR_OUT_3C  (
            .O(\INVU409_AUTOCONFIG.PR_OUT_3C_net ),
            .I(N__9897));
    INV \INVU409_AUTOCONFIG.LIDE_BASE_6C  (
            .O(\INVU409_AUTOCONFIG.LIDE_BASE_6C_net ),
            .I(N__9899));
    INV \INVU409_AUTOCONFIG.LIDE_BASE_2C  (
            .O(\INVU409_AUTOCONFIG.LIDE_BASE_2C_net ),
            .I(N__9904));
    INV \INVU409_AUTOCONFIG.LIDE_BASE_1C  (
            .O(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .I(N__9905));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_17_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_6_0_));
    defparam IN_MUX_bfv_17_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_7_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_17_7_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_9_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7961),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_9_LC_1_15_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_9_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_9_LC_1_15_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_9_LC_1_15_1  (
            .in0(N__4292),
            .in1(N__5351),
            .in2(N__4508),
            .in3(N__4484),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_3_LC_1_15_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_3_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_3_LC_1_15_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_3_LC_1_15_2  (
            .in0(N__4457),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4291),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_15_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_15_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_15_3  (
            .in0(N__4504),
            .in1(N__4463),
            .in2(N__4487),
            .in3(N__4483),
            .lcout(\U409_ADDRESS_DECODE.N_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_16_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_16_0  (
            .in0(N__4435),
            .in1(N__4366),
            .in2(N__4394),
            .in3(N__4414),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_10_LC_1_16_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_10_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_10_LC_1_16_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_10_LC_1_16_3  (
            .in0(N__4450),
            .in1(N__4436),
            .in2(N__4418),
            .in3(N__4393),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_0_LC_2_11_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_0_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_0_LC_2_11_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_0_LC_2_11_0  (
            .in0(N__4749),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5186),
            .lcout(N_100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_11_LC_2_14_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_11_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_11_LC_2_14_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_11_LC_2_14_1  (
            .in0(N__4677),
            .in1(N__4535),
            .in2(N__5740),
            .in3(N__4373),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_2_14_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_2_14_2 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_2_14_2  (
            .in0(N__4595),
            .in1(N__4340),
            .in2(N__4334),
            .in3(N__4331),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.N_61_i_LC_5_5_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.N_61_i_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.N_61_i_LC_5_5_6 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U409_ADDRESS_DECODE.N_61_i_LC_5_5_6  (
            .in0(N__4740),
            .in1(N__5326),
            .in2(N__5793),
            .in3(N__5220),
            .lcout(N_61_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_5_8_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_5_8_3 .LUT_INIT=16'b1100111101000111;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_5_8_3  (
            .in0(N__6286),
            .in1(N__6781),
            .in2(N__6238),
            .in3(N__6582),
            .lcout(\U409_AUTOCONFIG.PR_OUT_cnst_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_0_0_LC_5_9_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_0_0_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_0_0_LC_5_9_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_0_0_LC_5_9_0  (
            .in0(N__6642),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6468),
            .lcout(\U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_0_1_LC_5_10_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_0_1_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_0_1_LC_5_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a3_0_1_LC_5_10_2  (
            .in0(N__5792),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5210),
            .lcout(\U409_ADDRESS_DECODE.N_34_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_5_0_a3_LC_5_11_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_5_0_a3_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_5_0_a3_LC_5_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_5_0_a3_LC_5_11_0  (
            .in0(N__4879),
            .in1(N__4750),
            .in2(N__4828),
            .in3(N__4678),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACE_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_LC_5_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_LC_5_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_LC_5_11_4  (
            .in0(N__4880),
            .in1(N__10412),
            .in2(N__5135),
            .in3(N__5875),
            .lcout(N_89),
            .ltout(N_89_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_5_11_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_5_11_5 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_5_11_5  (
            .in0(N__4679),
            .in1(_gnd_net_),
            .in2(N__4601),
            .in3(N__5062),
            .lcout(N_94),
            .ltout(N_94_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_1_LC_5_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_1_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_1_LC_5_11_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_1_LC_5_11_6  (
            .in0(N__5209),
            .in1(N__5777),
            .in2(N__4598),
            .in3(N__4751),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_8_LC_5_14_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_8_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_8_LC_5_14_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_8_LC_5_14_1  (
            .in0(N__4583),
            .in1(N__4565),
            .in2(N__4547),
            .in3(N__4832),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CS0_LC_6_3_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CS0_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CS0_LC_6_3_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_ADDRESS_DECODE.CS0_LC_6_3_2  (
            .in0(N__8460),
            .in1(N__4816),
            .in2(N__4526),
            .in3(N__8518),
            .lcout(\U409_ADDRESS_DECODE.CSZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CS1_LC_6_3_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CS1_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CS1_LC_6_3_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_ADDRESS_DECODE.CS1_LC_6_3_3  (
            .in0(N__4817),
            .in1(N__4525),
            .in2(N__8522),
            .in3(N__8461),
            .lcout(\U409_ADDRESS_DECODE.CSZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_1_LC_6_4_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_1_LC_6_4_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_1_LC_6_4_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_1_LC_6_4_5  (
            .in0(N__4738),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5225),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_4_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_4_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_4_6  (
            .in0(N__5770),
            .in1(N__5330),
            .in2(N__4835),
            .in3(N__4827),
            .lcout(AUTOCONFIG_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_6_5_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_6_5_4 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_6_5_4  (
            .in0(N__4931),
            .in1(N__4911),
            .in2(N__5794),
            .in3(N__5138),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_6_6_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_6_6_1 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_6_6_1  (
            .in0(N__4739),
            .in1(N__5383),
            .in2(N__4671),
            .in3(N__4633),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_1_LC_6_6_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_1_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_1_LC_6_6_2 .LUT_INIT=16'b1111101000101010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_1_LC_6_6_2  (
            .in0(N__4634),
            .in1(N__6182),
            .in2(N__5647),
            .in3(N__5417),
            .lcout(LIDE_BASE_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .ce(),
            .sr(N__10130));
    defparam \U409_AUTOCONFIG.LIDE_BASE_3_LC_6_6_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_3_LC_6_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_3_LC_6_6_5 .LUT_INIT=16'b1111011111000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_3_LC_6_6_5  (
            .in0(N__6181),
            .in1(N__5641),
            .in2(N__6116),
            .in3(N__4613),
            .lcout(LIDE_BASE_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .ce(),
            .sr(N__10130));
    defparam \U409_AUTOCONFIG.LIDE_BASE_4_LC_6_6_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_4_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_4_LC_6_6_6 .LUT_INIT=16'b1101111111000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_4_LC_6_6_6  (
            .in0(N__6104),
            .in1(N__5459),
            .in2(N__5648),
            .in3(N__4625),
            .lcout(LIDE_BASE_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_1C_net ),
            .ce(),
            .sr(N__10130));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_6_7_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_6_7_1 .LUT_INIT=16'b1000001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_6_7_1  (
            .in0(N__5018),
            .in1(N__5893),
            .in2(N__5137),
            .in3(N__7058),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_6_7_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_6_7_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_6_7_2  (
            .in0(N__7214),
            .in1(N__5273),
            .in2(N__5972),
            .in3(N__5282),
            .lcout(\U409_AUTOCONFIG.un1_STATE_6Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_6_7_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_6_7_4 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_6_7_4  (
            .in0(N__5224),
            .in1(N__4624),
            .in2(N__4863),
            .in3(N__4612),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_6_7_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_LC_6_7_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_LC_6_7_5  (
            .in0(N__4961),
            .in1(N__5663),
            .in2(N__4955),
            .in3(N__4952),
            .lcout(ATA_SPACE),
            .ltout(ATA_SPACE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_6_7_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_LC_6_7_6 .LUT_INIT=16'b1010101000100000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_LC_6_7_6  (
            .in0(N__10393),
            .in1(N__7613),
            .in2(N__4946),
            .in3(N__4942),
            .lcout(\U409_ADDRESS_DECODE.ATA_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9903),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_6_8_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_6_8_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_6_8_1  (
            .in0(N__4927),
            .in1(N__5128),
            .in2(N__5782),
            .in3(N__4912),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_2_LC_6_8_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_2_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_2_LC_6_8_3 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a3_2_LC_6_8_3  (
            .in0(N__5867),
            .in1(N__5127),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_6_8_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_6_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_6_8_5  (
            .in0(_gnd_net_),
            .in1(N__7393),
            .in2(_gnd_net_),
            .in3(N__4943),
            .lcout(U409_ADDRESS_DECODE_un1_ATA_ENn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_0_1_LC_6_9_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_0_1_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_0_1_LC_6_9_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_0_1_LC_6_9_0  (
            .in0(N__6456),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6643),
            .lcout(\U409_AUTOCONFIG.N_193_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_1_LC_6_9_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_1_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_1_LC_6_9_1 .LUT_INIT=16'b0100000001000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_1_LC_6_9_1  (
            .in0(N__5854),
            .in1(N__5069),
            .in2(N__10424),
            .in3(_gnd_net_),
            .lcout(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_3_LC_6_9_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_3_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_3_LC_6_9_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a3_3_LC_6_9_2  (
            .in0(N__4873),
            .in1(N__4916),
            .in2(N__5781),
            .in3(N__5205),
            .lcout(\U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_0_LC_6_9_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_0_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a3_0_LC_6_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a3_0_LC_6_9_3  (
            .in0(N__5853),
            .in1(N__5372),
            .in2(N__5136),
            .in3(N__4872),
            .lcout(\U409_ADDRESS_DECODE.N_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_14_2_LC_6_9_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_14_2_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_14_2_LC_6_9_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_AUTOCONFIG.un1_A_14_2_LC_6_9_4  (
            .in0(N__6578),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6780),
            .lcout(\U409_AUTOCONFIG.N_227_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a3_LC_6_9_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a3_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_0_a3_LC_6_9_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_0_a3_LC_6_9_5  (
            .in0(N__10420),
            .in1(N__5068),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACE ),
            .ltout(\U409_ADDRESS_DECODE.Z2_SPACE_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_6_9_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_6_9_6 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_6_9_6  (
            .in0(N__5009),
            .in1(N__5003),
            .in2(N__4997),
            .in3(N__4994),
            .lcout(ROMEN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_0_2_LC_6_10_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_0_2_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_0_2_LC_6_10_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_0_2_LC_6_10_0  (
            .in0(N__5945),
            .in1(N__6015),
            .in2(N__4976),
            .in3(N__5269),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_o3_2_LC_6_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_o3_2_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_o3_2_LC_6_10_1 .LUT_INIT=16'b1100110001001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_o3_2_LC_6_10_1  (
            .in0(N__6857),
            .in1(N__10394),
            .in2(N__4988),
            .in3(N__6672),
            .lcout(\U409_AUTOCONFIG.N_214_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_LC_6_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_LC_6_10_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_LC_6_10_2  (
            .in0(N__4985),
            .in1(N__5272),
            .in2(N__5360),
            .in3(N__6762),
            .lcout(\U409_AUTOCONFIG.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_4_LC_6_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_4_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_4_LC_6_10_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_4_LC_6_10_4  (
            .in0(N__5944),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6014),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_4 ),
            .ltout(\U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_2_LC_6_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_2_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_2_LC_6_10_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_2_LC_6_10_5  (
            .in0(N__5271),
            .in1(N__4975),
            .in2(N__4964),
            .in3(N__6673),
            .lcout(\U409_AUTOCONFIG.N_192 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a2_1_LC_6_10_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a2_1_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a2_1_LC_6_10_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a2_1_LC_6_10_6  (
            .in0(N__6858),
            .in1(N__5270),
            .in2(N__5955),
            .in3(N__6016),
            .lcout(\U409_AUTOCONFIG.N_198 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_10_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_10_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_10_7  (
            .in0(N__5371),
            .in1(N__5556),
            .in2(N__5871),
            .in3(N__5033),
            .lcout(CIA_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_0_LC_6_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_0_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_0_LC_6_11_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_0_LC_6_11_3  (
            .in0(N__6529),
            .in1(N__6840),
            .in2(_gnd_net_),
            .in3(N__6671),
            .lcout(\U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PORTSIZE_1_LC_6_11_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PORTSIZE_1_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PORTSIZE_1_LC_6_11_4 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \U409_AUTOCONFIG.PORTSIZE_1_LC_6_11_4  (
            .in0(N__5350),
            .in1(N__5319),
            .in2(N__7156),
            .in3(N__5773),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.PORTSIZEZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PORTSIZE_0_i_LC_6_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PORTSIZE_0_i_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PORTSIZE_0_i_LC_6_11_5 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U409_AUTOCONFIG.PORTSIZE_0_i_LC_6_11_5  (
            .in0(N__10717),
            .in1(N__7461),
            .in2(N__5306),
            .in3(N__8605),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_STATE_6_0_LC_6_11_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_STATE_6_0_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_STATE_6_0_LC_6_11_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_AUTOCONFIG.un1_STATE_6_0_LC_6_11_6  (
            .in0(N__6002),
            .in1(N__6761),
            .in2(N__6856),
            .in3(N__6530),
            .lcout(\U409_AUTOCONFIG.un1_STATE_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_13_3_LC_6_11_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_13_3_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_13_3_LC_6_11_7 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U409_AUTOCONFIG.un1_A_13_3_LC_6_11_7  (
            .in0(N__6760),
            .in1(N__5250),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_AUTOCONFIG.un1_A_13Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_1_LC_6_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_1_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_1_LC_6_12_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_1_LC_6_12_3  (
            .in0(N__5835),
            .in1(N__5187),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_1 ),
            .ltout(\U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_12_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_12_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_12_4  (
            .in0(N__5771),
            .in1(N__5557),
            .in2(N__5141),
            .in3(N__5029),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_0_a3_LC_6_12_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_0_a3_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_0_a3_LC_6_12_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_4_0_a3_LC_6_12_6  (
            .in0(N__5106),
            .in1(N__5061),
            .in2(_gnd_net_),
            .in3(N__10413),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACE_4 ),
            .ltout(\U409_ADDRESS_DECODE.CIA_SPACE_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_12_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_12_7 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_12_7  (
            .in0(N__5558),
            .in1(N__5772),
            .in2(N__5543),
            .in3(N__5540),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_4_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.D_1_i_LC_7_4_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.D_1_i_LC_7_4_0  (
            .in0(N__7102),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7624),
            .lcout(D_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_4_LC_7_5_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_4_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_4_LC_7_5_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_4_LC_7_5_0  (
            .in0(N__5468),
            .in1(N__7104),
            .in2(N__7622),
            .in3(N__6095),
            .lcout(\U409_AUTOCONFIG.N_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_6_LC_7_5_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_6_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_6_LC_7_5_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_6_LC_7_5_1  (
            .in0(N__6097),
            .in1(N__7611),
            .in2(N__7124),
            .in3(N__5453),
            .lcout(\U409_AUTOCONFIG.N_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_2_LC_7_5_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_2_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_2_LC_7_5_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_2_LC_7_5_3  (
            .in0(N__6170),
            .in1(N__7125),
            .in2(N__7604),
            .in3(N__5452),
            .lcout(\U409_AUTOCONFIG.N_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_5_LC_7_5_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_5_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_5_LC_7_5_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_5_LC_7_5_4  (
            .in0(N__5435),
            .in1(N__7105),
            .in2(N__7623),
            .in3(N__6096),
            .lcout(\U409_AUTOCONFIG.N_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_1_LC_7_5_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_1_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_1_LC_7_5_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_1_LC_7_5_6  (
            .in0(N__5434),
            .in1(N__7575),
            .in2(N__6180),
            .in3(N__7103),
            .lcout(\U409_AUTOCONFIG.N_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_7_5_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_7_5_7 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_7_5_7  (
            .in0(N__5567),
            .in1(N__7358),
            .in2(N__5594),
            .in3(N__7063),
            .lcout(D_OUT_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_2_LC_7_6_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_2_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_2_LC_7_6_1 .LUT_INIT=16'b1011101011110000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_2_LC_7_6_1  (
            .in0(N__5393),
            .in1(N__6179),
            .in2(N__5387),
            .in3(N__5633),
            .lcout(LIDE_BASE_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_2C_net ),
            .ce(),
            .sr(N__10129));
    defparam \U409_AUTOCONFIG.LIDE_BASE_7_LC_7_6_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_7_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_7_LC_7_6_2 .LUT_INIT=16'b1101111111000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_7_LC_7_6_2  (
            .in0(N__6099),
            .in1(N__5900),
            .in2(N__5646),
            .in3(N__5894),
            .lcout(LIDE_BASE_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_2C_net ),
            .ce(),
            .sr(N__10129));
    defparam \U409_AUTOCONFIG.LIDE_BASE_5_LC_7_6_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_5_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_5_LC_7_6_3 .LUT_INIT=16'b1101110011110000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_5_LC_7_6_3  (
            .in0(N__6098),
            .in1(N__5882),
            .in2(N__5681),
            .in3(N__5634),
            .lcout(LIDE_BASE_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_2C_net ),
            .ce(),
            .sr(N__10129));
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_7_6_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.CONFIGURED_LC_7_6_7 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U409_AUTOCONFIG.CONFIGURED_LC_7_6_7  (
            .in0(N__7181),
            .in1(N__7357),
            .in2(_gnd_net_),
            .in3(N__7062),
            .lcout(CONFIGURED),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_2C_net ),
            .ce(),
            .sr(N__10129));
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_7_7_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_7_7_0 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_7_7_0  (
            .in0(N__5876),
            .in1(N__5602),
            .in2(N__5795),
            .in3(N__5674),
            .lcout(\U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_6_LC_7_7_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_6_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_6_LC_7_7_2 .LUT_INIT=16'b1101111111000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_6_LC_7_7_2  (
            .in0(N__6103),
            .in1(N__5657),
            .in2(N__5645),
            .in3(N__5603),
            .lcout(LIDE_BASE_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_BASE_6C_net ),
            .ce(),
            .sr(N__10128));
    defparam \U409_AUTOCONFIG.PR_OUT_3_LC_7_8_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_3_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PR_OUT_3_LC_7_8_4 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_3_LC_7_8_4  (
            .in0(N__6026),
            .in1(N__10375),
            .in2(N__6587),
            .in3(N__6285),
            .lcout(\U409_AUTOCONFIG.PR_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.PR_OUT_3C_net ),
            .ce(N__6986),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_2_LC_7_8_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_2_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PR_OUT_2_LC_7_8_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_2_LC_7_8_7  (
            .in0(N__10374),
            .in1(N__5582),
            .in2(_gnd_net_),
            .in3(N__7012),
            .lcout(\U409_AUTOCONFIG.PR_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.PR_OUT_3C_net ),
            .ce(N__6986),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_9_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_9_3 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_9_3  (
            .in0(N__6364),
            .in1(N__6038),
            .in2(_gnd_net_),
            .in3(N__6922),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_3C_net ),
            .ce(N__6978),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_7_9_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_7_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_7_9_4  (
            .in0(N__6044),
            .in1(N__5573),
            .in2(_gnd_net_),
            .in3(N__7268),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_9_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_9_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(N__6307),
            .in2(_gnd_net_),
            .in3(N__6037),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_3C_net ),
            .ce(N__6978),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_3_LC_7_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_3_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_3_LC_7_10_1 .LUT_INIT=16'b1001000000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_3_LC_7_10_1  (
            .in0(N__6577),
            .in1(N__6763),
            .in2(N__6469),
            .in3(N__6677),
            .lcout(\U409_AUTOCONFIG.N_225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_3_LC_7_10_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_3_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_3_LC_7_10_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_3_LC_7_10_2  (
            .in0(N__6676),
            .in1(N__10377),
            .in2(N__6878),
            .in3(N__6576),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_LC_7_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_LC_7_10_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_LC_7_10_3  (
            .in0(N__6017),
            .in1(N__5949),
            .in2(N__6029),
            .in3(N__5917),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxaZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_3_LC_7_10_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_3_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNO_0_3_LC_7_10_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNO_0_3_LC_7_10_4  (
            .in0(N__6764),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6455),
            .lcout(\U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_7_11_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_7_11_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_7_11_0  (
            .in0(N__5964),
            .in1(N__6674),
            .in2(N__6013),
            .in3(N__6531),
            .lcout(\U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_13_0_LC_7_11_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_13_0_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_13_0_LC_7_11_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U409_AUTOCONFIG.un1_A_13_0_LC_7_11_5  (
            .in0(N__6675),
            .in1(N__6001),
            .in2(_gnd_net_),
            .in3(N__6874),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.un1_A_13Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.un1_A_13_LC_7_11_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.un1_A_13_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.un1_A_13_LC_7_11_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_AUTOCONFIG.un1_A_13_LC_7_11_6  (
            .in0(N__5965),
            .in1(N__5918),
            .in2(N__5903),
            .in3(N__6532),
            .lcout(\U409_AUTOCONFIG.un1_AZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_7_LC_8_5_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_7_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_7_LC_8_5_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_7_LC_8_5_1  (
            .in0(N__6142),
            .in1(N__7141),
            .in2(N__7612),
            .in3(N__6094),
            .lcout(\U409_AUTOCONFIG.N_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_5_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_5_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_5_6  (
            .in0(_gnd_net_),
            .in1(N__7296),
            .in2(_gnd_net_),
            .in3(N__7254),
            .lcout(\U409_AUTOCONFIG.D_OUT_sm0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_8_6_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_8_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_8_6_0  (
            .in0(N__7250),
            .in1(N__6383),
            .in2(_gnd_net_),
            .in3(N__6269),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_8_6_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_8_6_1 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_8_6_1  (
            .in0(N__6206),
            .in1(N__7360),
            .in2(N__6197),
            .in3(N__7065),
            .lcout(D_OUT_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_LC_8_6_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_LC_8_6_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_LC_8_6_3  (
            .in0(N__6686),
            .in1(N__7294),
            .in2(_gnd_net_),
            .in3(N__7249),
            .lcout(\U409_AUTOCONFIG.LIDE_BASE_10 ),
            .ltout(\U409_AUTOCONFIG.LIDE_BASE_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_3_LC_8_6_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_3_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_BASE_RNO_0_3_LC_8_6_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_BASE_RNO_0_3_LC_8_6_4  (
            .in0(N__6149),
            .in1(N__7142),
            .in2(N__6119),
            .in3(N__7621),
            .lcout(\U409_AUTOCONFIG.N_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_0_LC_8_6_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_0_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_0_LC_8_6_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_0_LC_8_6_5  (
            .in0(N__6685),
            .in1(N__7293),
            .in2(_gnd_net_),
            .in3(N__7248),
            .lcout(\U409_AUTOCONFIG.LIDE_BASE_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_8_6_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_8_6_6 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_8_6_6  (
            .in0(N__7295),
            .in1(N__6392),
            .in2(N__7263),
            .in3(N__6215),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.LIDE_OUT_RNIOO061Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNID8KD2_1_LC_8_6_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNID8KD2_1_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNID8KD2_1_LC_8_6_7 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNID8KD2_1_LC_8_6_7  (
            .in0(N__6995),
            .in1(N__7359),
            .in2(N__6059),
            .in3(N__7064),
            .lcout(D_OUT_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_8_7_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_8_7_6 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_8_7_6  (
            .in0(N__6329),
            .in1(N__6221),
            .in2(N__7264),
            .in3(N__7301),
            .lcout(),
            .ltout(\U409_AUTOCONFIG.LIDE_OUT_RNIMM061Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_RNIA5KD2_0_LC_8_7_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_RNIA5KD2_0_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_RNIA5KD2_0_LC_8_7_7 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_RNIA5KD2_0_LC_8_7_7  (
            .in0(N__7364),
            .in1(N__6323),
            .in2(N__6413),
            .in3(N__7066),
            .lcout(D_OUT_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_8_8_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_1_LC_8_8_0 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_1_LC_8_8_0  (
            .in0(N__6932),
            .in1(N__6373),
            .in2(N__10405),
            .in3(N__6296),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(N__6985),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_8_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_8_1 .LUT_INIT=16'b1010101110101010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_8_1  (
            .in0(N__6374),
            .in1(N__6902),
            .in2(N__7025),
            .in3(N__6923),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(N__6985),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_8_8_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_0_LC_8_8_2 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_0_LC_8_8_2  (
            .in0(N__6791),
            .in1(N__6372),
            .in2(N__6953),
            .in3(N__6353),
            .lcout(\U409_AUTOCONFIG.LIDE_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(N__6985),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_0_LC_8_8_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_0_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PR_OUT_0_LC_8_8_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_0_LC_8_8_3  (
            .in0(N__7023),
            .in1(N__6260),
            .in2(N__10403),
            .in3(N__6940),
            .lcout(\U409_AUTOCONFIG.PR_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(N__6985),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_8_8_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_8_8_4 .LUT_INIT=16'b0100000001010000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_8_8_4  (
            .in0(N__6901),
            .in1(N__6782),
            .in2(N__6317),
            .in3(N__6295),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(N__6985),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_8_8_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_8_8_5 .LUT_INIT=16'b0010001000000010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_8_8_5  (
            .in0(N__10363),
            .in1(N__6259),
            .in2(N__6245),
            .in3(N__6931),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(N__6985),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_8_8_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_8_8_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_8_8_6  (
            .in0(N__6424),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10364),
            .lcout(\U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(N__6985),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_1_LC_8_8_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_1_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.PR_OUT_1_LC_8_8_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_1_LC_8_8_7  (
            .in0(N__7024),
            .in1(N__6425),
            .in2(N__10404),
            .in3(N__6941),
            .lcout(\U409_AUTOCONFIG.PR_OUTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.LIDE_OUT_1C_net ),
            .ce(N__6985),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNI10V92_1_LC_8_9_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNI10V92_1_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNI10V92_1_LC_8_9_1 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNI10V92_1_LC_8_9_1  (
            .in0(N__7664),
            .in1(N__7502),
            .in2(N__10408),
            .in3(N__7675),
            .lcout(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_8_9_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_8_9_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_8_9_2  (
            .in0(N__6918),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6895),
            .lcout(\U409_AUTOCONFIG.N_184_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_a2_0_LC_8_9_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_a2_0_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.PR_OUT_cnst_i_a2_0_LC_8_9_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_AUTOCONFIG.PR_OUT_cnst_i_a2_0_LC_8_9_4  (
            .in0(N__6586),
            .in1(N__6779),
            .in2(_gnd_net_),
            .in3(N__6485),
            .lcout(\U409_AUTOCONFIG.N_167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_x3_0_LC_8_9_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_x3_0_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_x3_0_LC_8_9_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_x3_0_LC_8_9_5  (
            .in0(N__6778),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6585),
            .lcout(\U409_AUTOCONFIG.N_213_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_i_o3_3_LC_8_10_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_i_o3_3_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_cnst_i_o3_3_LC_8_10_3 .LUT_INIT=16'b1100110010001100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_cnst_i_o3_3_LC_8_10_3  (
            .in0(N__6777),
            .in1(N__10376),
            .in2(N__6483),
            .in3(N__6584),
            .lcout(\U409_AUTOCONFIG.N_182_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_2_LC_8_10_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_2_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_2_LC_8_10_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_2_LC_8_10_5  (
            .in0(N__6776),
            .in1(N__6583),
            .in2(N__6482),
            .in3(N__6679),
            .lcout(\U409_AUTOCONFIG.N_223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_8_11_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_8_11_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_8_11_1  (
            .in0(N__6769),
            .in1(N__6884),
            .in2(_gnd_net_),
            .in3(N__6873),
            .lcout(\U409_AUTOCONFIG.N_190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_LC_8_11_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_LC_8_11_3 .LUT_INIT=16'b0000110100000000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_LC_8_11_3  (
            .in0(N__6768),
            .in1(N__6678),
            .in2(N__6562),
            .in3(N__6484),
            .lcout(\U409_AUTOCONFIG.N_222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.LV_SPACE_LC_8_11_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LV_SPACE_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.LV_SPACE_LC_8_11_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_AUTOCONFIG.LV_SPACE_LC_8_11_7  (
            .in0(N__7444),
            .in1(N__7472),
            .in2(N__7157),
            .in3(N__7400),
            .lcout(BUFENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_9_6_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_9_6_0 .SEQ_MODE=4'b1001;
    defparam \U409_AUTOCONFIG.CONFIGENn_LC_9_6_0 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \U409_AUTOCONFIG.CONFIGENn_LC_9_6_0  (
            .in0(N__7356),
            .in1(N__7312),
            .in2(_gnd_net_),
            .in3(N__7173),
            .lcout(CONFIGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .ce(),
            .sr(N__10127));
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_9_6_5 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.LIDE_CONF_LC_9_6_5 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U409_AUTOCONFIG.LIDE_CONF_LC_9_6_5  (
            .in0(N__7255),
            .in1(N__7174),
            .in2(_gnd_net_),
            .in3(N__7297),
            .lcout(\U409_AUTOCONFIG.LIDE_CONFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .ce(),
            .sr(N__10127));
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_9_6_6 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.BRIDGE_CONF_LC_9_6_6 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U409_AUTOCONFIG.BRIDGE_CONF_LC_9_6_6  (
            .in0(N__7199),
            .in1(N__7213),
            .in2(_gnd_net_),
            .in3(N__7256),
            .lcout(\U409_AUTOCONFIG.BRIDGE_CONFZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.CONFIGENnC_net ),
            .ce(),
            .sr(N__10127));
    defparam \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_9_7_4 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_9_7_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__7500),
            .in2(_gnd_net_),
            .in3(N__7650),
            .lcout(\U409_AUTOCONFIG.STATE_d_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIDEFO1_0_LC_9_7_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIDEFO1_0_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIDEFO1_0_LC_9_7_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIDEFO1_0_LC_9_7_7  (
            .in0(N__7651),
            .in1(N__7198),
            .in2(_gnd_net_),
            .in3(N__7501),
            .lcout(\U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_0_LC_9_8_0 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_0_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.STATE_0_LC_9_8_0 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \U409_AUTOCONFIG.STATE_0_LC_9_8_0  (
            .in0(N__7503),
            .in1(N__7653),
            .in2(N__10406),
            .in3(N__7676),
            .lcout(\U409_AUTOCONFIG.STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_1_LC_9_8_2 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_1_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.STATE_1_LC_9_8_2 .LUT_INIT=16'b0001000010100000;
    LogicCell40 \U409_AUTOCONFIG.STATE_1_LC_9_8_2  (
            .in0(N__7504),
            .in1(N__7620),
            .in2(N__10407),
            .in3(N__7654),
            .lcout(\U409_AUTOCONFIG.STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_LC_9_9_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_START_LC_9_9_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_AUTOCONFIG.AC_START_LC_9_9_1  (
            .in0(N__7152),
            .in1(N__8578),
            .in2(_gnd_net_),
            .in3(N__7070),
            .lcout(\U409_AUTOCONFIG.AC_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9890),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_START_RNI04BC_LC_9_9_3 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_START_RNI04BC_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.AC_START_RNI04BC_LC_9_9_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_AUTOCONFIG.AC_START_RNI04BC_LC_9_9_3  (
            .in0(N__7697),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7682),
            .lcout(\U409_AUTOCONFIG.STATE4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.STATE_RNIJFAU_0_LC_9_9_7 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.STATE_RNIJFAU_0_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_AUTOCONFIG.STATE_RNIJFAU_0_LC_9_9_7 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \U409_AUTOCONFIG.STATE_RNIJFAU_0_LC_9_9_7  (
            .in0(N__7574),
            .in1(N__7652),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_AUTOCONFIG.AC_TACK_LC_9_10_1 .C_ON=1'b0;
    defparam \U409_AUTOCONFIG.AC_TACK_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_AUTOCONFIG.AC_TACK_LC_9_10_1 .LUT_INIT=16'b1110111011001000;
    LogicCell40 \U409_AUTOCONFIG.AC_TACK_LC_9_10_1  (
            .in0(N__7720),
            .in1(N__7658),
            .in2(N__7625),
            .in3(N__7508),
            .lcout(AC_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_AUTOCONFIG.AC_TACKC_net ),
            .ce(),
            .sr(N__10124));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_12_0 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_12_0  (
            .in0(N__7468),
            .in1(N__7445),
            .in2(N__10419),
            .in3(N__7427),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_9_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_9_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__7881),
            .in2(_gnd_net_),
            .in3(N__7846),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_11_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_11_2 .LUT_INIT=16'b0011001110111011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_11_2  (
            .in0(N__7736),
            .in1(N__7409),
            .in2(_gnd_net_),
            .in3(N__8110),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .ce(),
            .sr(N__8091));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_10_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_10_11_5 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_10_11_5  (
            .in0(N__7876),
            .in1(N__8044),
            .in2(N__7706),
            .in3(N__7940),
            .lcout(\U409_TRANSFER_ACK.N_53 ),
            .ltout(\U409_TRANSFER_ACK.N_53_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_10_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_10_11_6 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_10_11_6  (
            .in0(N__9931),
            .in1(N__8569),
            .in2(N__7403),
            .in3(N__8109),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_11_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_11_7 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_11_7  (
            .in0(N__7877),
            .in1(N__7934),
            .in2(N__7739),
            .in3(N__7847),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .ce(),
            .sr(N__8091));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_12_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_12_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_12_1  (
            .in0(N__8048),
            .in1(N__8005),
            .in2(_gnd_net_),
            .in3(N__7790),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__8084));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_12_5 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_12_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_12_5  (
            .in0(N__7929),
            .in1(N__7882),
            .in2(_gnd_net_),
            .in3(N__7789),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__8084));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_10_3 .LUT_INIT=16'b0100000001010000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_10_3  (
            .in0(N__8197),
            .in1(N__8216),
            .in2(N__10362),
            .in3(N__8172),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_10_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_10_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_10_5  (
            .in0(N__10305),
            .in1(N__8192),
            .in2(_gnd_net_),
            .in3(N__8215),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_11_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_11_10_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(N__8227),
            .in2(_gnd_net_),
            .in3(N__7735),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_10_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_10_7  (
            .in0(N__7724),
            .in1(N__8297),
            .in2(N__7709),
            .in3(N__8966),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_11_2 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_11_2  (
            .in0(N__8034),
            .in1(N__8130),
            .in2(N__8000),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_11_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_11_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_11_11_5  (
            .in0(N__7898),
            .in1(N__7843),
            .in2(N__7819),
            .in3(N__7767),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_11_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_11_6  (
            .in0(N__7987),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8129),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_11_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_11_11_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_11_11_7  (
            .in0(N__7875),
            .in1(N__8033),
            .in2(N__7949),
            .in3(N__7946),
            .lcout(\U409_TRANSFER_ACK.N_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_12_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_12_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_12_2  (
            .in0(N__7817),
            .in1(N__7969),
            .in2(_gnd_net_),
            .in3(N__7792),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__8092));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_11_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_11_12_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_11_12_3  (
            .in0(N__7900),
            .in1(N__7844),
            .in2(N__7820),
            .in3(N__7768),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_12_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_12_4 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_12_4  (
            .in0(N__7933),
            .in1(N__7901),
            .in2(N__7913),
            .in3(N__7791),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__8092));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_11_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_11_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_11_12_5  (
            .in0(N__7899),
            .in1(N__8131),
            .in2(N__7883),
            .in3(N__7845),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_12_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_12_6 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_12_6  (
            .in0(N__7818),
            .in1(N__7970),
            .in2(N__7772),
            .in3(N__7793),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net ),
            .ce(),
            .sr(N__8092));
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_6.C_ON=1'b0;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9933),
            .lcout(GB_BUFFER_CLK40_IN_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_9_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_9_7  (
            .in0(N__8582),
            .in1(N__8266),
            .in2(N__9935),
            .in3(N__8278),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_12_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_LC_12_10_2 .LUT_INIT=16'b0011000011110001;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_LC_12_10_2  (
            .in0(N__8174),
            .in1(N__8193),
            .in2(N__9100),
            .in3(N__8213),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .ce(),
            .sr(N__10120));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_10_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_10_4  (
            .in0(N__8947),
            .in1(N__8279),
            .in2(N__8267),
            .in3(N__8228),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .ce(),
            .sr(N__10120));
    defparam \U409_TRANSFER_ACK.TACK_OUT_LC_12_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUT_LC_12_10_5 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.TACK_OUT_LC_12_10_5 .LUT_INIT=16'b1100111011001010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUT_LC_12_10_5  (
            .in0(N__8214),
            .in1(N__8143),
            .in2(N__8198),
            .in3(N__8173),
            .lcout(TACK_OUT),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_ENC_net ),
            .ce(),
            .sr(N__10120));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_11_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_11_1  (
            .in0(N__8043),
            .in1(N__8132),
            .in2(_gnd_net_),
            .in3(N__8006),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__8096));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_11_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_11_6 .LUT_INIT=16'b1101110000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_11_6  (
            .in0(N__8576),
            .in1(N__8042),
            .in2(N__9934),
            .in3(N__8111),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net ),
            .ce(),
            .sr(N__8096));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_12_12_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_12_12_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_12_12_0  (
            .in0(N__8054),
            .in1(N__8041),
            .in2(_gnd_net_),
            .in3(N__8001),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_5.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_5.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_19_5 (
            .in0(N__10271),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_13_9_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_13_9_0 .LUT_INIT=16'b0001001001011010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_13_9_0  (
            .in0(N__8387),
            .in1(N__8333),
            .in2(N__8363),
            .in3(N__8324),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10912),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMUMD1_7_LC_13_9_2 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMUMD1_7_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMUMD1_7_LC_13_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIMUMD1_7_LC_13_9_2  (
            .in0(N__8756),
            .in1(N__8701),
            .in2(N__8734),
            .in3(N__8636),
            .lcout(\U409_CIA.CLK_CIA6_3 ),
            .ltout(\U409_CIA.CLK_CIA6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_13_9_3 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_13_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_1_LC_13_9_3  (
            .in0(N__8672),
            .in1(N__8385),
            .in2(N__8342),
            .in3(N__8339),
            .lcout(\U409_CIA.CLK_CIA_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_13_9_4 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_13_9_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_2_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__8790),
            .in2(_gnd_net_),
            .in3(N__8411),
            .lcout(\U409_CIA.un1_CIA_CLK_COUNT_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_13_9_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_13_9_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_13_9_6  (
            .in0(N__8386),
            .in1(N__8791),
            .in2(N__8417),
            .in3(N__8702),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_2_0 ),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_13_9_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_13_9_7 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_13_9_7  (
            .in0(N__8323),
            .in1(N__8795),
            .in2(N__8327),
            .in3(N__8348),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10912),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_13_10_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_13_10_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_13_10_4  (
            .in0(N__8729),
            .in1(N__8637),
            .in2(N__8762),
            .in3(N__8674),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNI9DRM_2_LC_13_10_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNI9DRM_2_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNI9DRM_2_LC_13_10_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNI9DRM_2_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__8383),
            .in2(_gnd_net_),
            .in3(N__8413),
            .lcout(\U409_CIA.CLK_CIA6_0 ),
            .ltout(\U409_CIA.CLK_CIA6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_13_10_6 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_13_10_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_0_LC_13_10_6  (
            .in0(N__8794),
            .in1(N__8673),
            .in2(N__8315),
            .in3(N__8312),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_LC_13_10_7 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_LC_13_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLK_CIA_LC_13_10_7 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \U409_CIA.CLK_CIA_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__8895),
            .in2(N__8306),
            .in3(N__8303),
            .lcout(CLK_CIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10910),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_11_6 .LUT_INIT=16'b1010001110100010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_11_6  (
            .in0(N__8293),
            .in1(N__9213),
            .in2(N__8591),
            .in3(N__9305),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(N__10121));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a4_1_LC_13_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a4_1_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a4_1_LC_13_12_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a4_1_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__8577),
            .in2(_gnd_net_),
            .in3(N__9927),
            .lcout(\U409_TRANSFER_ACK.N_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNI692L_0_LC_14_5_1 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNI692L_0_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNI692L_0_LC_14_5_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_CIA.VMA_RNI692L_0_LC_14_5_1  (
            .in0(N__10290),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10175),
            .lcout(CIA_ENABLE),
            .ltout(CIA_ENABLE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_14_5_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_14_5_2 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8525),
            .in3(N__8517),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_14_5_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_14_5_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_14_5_4  (
            .in0(_gnd_net_),
            .in1(N__8471),
            .in2(_gnd_net_),
            .in3(N__8465),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_14_9_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_14_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__8634),
            .in2(N__8705),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_14_9_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_14_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__8412),
            .in2(_gnd_net_),
            .in3(N__8390),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__10911),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_14_9_2 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_14_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__8384),
            .in2(_gnd_net_),
            .in3(N__8354),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_14_9_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_14_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__8671),
            .in2(_gnd_net_),
            .in3(N__8351),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__10911),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_14_9_4 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_14_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__8793),
            .in2(_gnd_net_),
            .in3(N__8804),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_14_9_5 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_14_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_6_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__8761),
            .in2(_gnd_net_),
            .in3(N__8801),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ),
            .clk(N__10911),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_14_9_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_14_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_7_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__8733),
            .in2(_gnd_net_),
            .in3(N__8798),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10911),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_14_9_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_14_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_14_9_7  (
            .in0(N__8635),
            .in1(N__8700),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10911),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_14_10_0 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_14_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_14_10_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_14_10_0  (
            .in0(N__8704),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10909),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_1_LC_14_10_5 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_1_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_1_LC_14_10_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_CIA.VMA_RNO_1_LC_14_10_5  (
            .in0(N__8792),
            .in1(N__8760),
            .in2(N__8735),
            .in3(N__8703),
            .lcout(),
            .ltout(\U409_CIA.un1_CIA_CLK_COUNT_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_14_10_6 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_14_10_6 .LUT_INIT=16'b0100000010000000;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_14_10_6  (
            .in0(N__8675),
            .in1(N__8648),
            .in2(N__8642),
            .in3(N__8638),
            .lcout(),
            .ltout(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_14_10_7 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_14_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_14_10_7 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \U409_CIA.VMA_LC_14_10_7  (
            .in0(N__8639),
            .in1(N__8609),
            .in2(N__8594),
            .in3(N__10164),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10909),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_14_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_14_11_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_14_11_2  (
            .in0(N__9236),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9268),
            .lcout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_14_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_14_11_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_14_11_5  (
            .in0(N__9298),
            .in1(N__9266),
            .in2(N__9212),
            .in3(N__9235),
            .lcout(\U409_TRANSFER_ACK.N_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI1MEE_1_LC_14_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI1MEE_1_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI1MEE_1_LC_14_11_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI1MEE_1_LC_14_11_6  (
            .in0(N__9234),
            .in1(N__9198),
            .in2(_gnd_net_),
            .in3(N__9297),
            .lcout(\U409_TRANSFER_ACK.N_19 ),
            .ltout(\U409_TRANSFER_ACK.N_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_14_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_14_11_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_14_11_7  (
            .in0(N__8940),
            .in1(N__9171),
            .in2(N__8855),
            .in3(N__9267),
            .lcout(\U409_TRANSFER_ACK.N_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_LC_14_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_14_12_3 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_14_12_3 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_LC_14_12_3  (
            .in0(N__8827),
            .in1(N__8852),
            .in2(_gnd_net_),
            .in3(N__8846),
            .lcout(ROMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROMENnC_net ),
            .ce(),
            .sr(N__10122));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_15_7_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_15_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_15_7_0  (
            .in0(_gnd_net_),
            .in1(N__9405),
            .in2(N__9487),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_15_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_15_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_15_7_1  (
            .in0(_gnd_net_),
            .in1(N__9421),
            .in2(_gnd_net_),
            .in3(N__8816),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__10786),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_15_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_15_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_15_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(N__9502),
            .in2(_gnd_net_),
            .in3(N__8813),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__10786),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_15_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_15_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_15_7_3  (
            .in0(_gnd_net_),
            .in1(N__9364),
            .in2(_gnd_net_),
            .in3(N__8810),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_15_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_15_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_15_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_15_7_4  (
            .in0(_gnd_net_),
            .in1(N__9532),
            .in2(_gnd_net_),
            .in3(N__8807),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__10786),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_15_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_15_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(N__9445),
            .in2(_gnd_net_),
            .in3(N__8882),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_15_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_15_7_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_15_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(N__8998),
            .in2(_gnd_net_),
            .in3(N__8879),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__10786),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_15_7_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_15_7_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(N__9964),
            .in2(_gnd_net_),
            .in3(N__8876),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_15_8_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_15_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__9679),
            .in2(_gnd_net_),
            .in3(N__8873),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_15_8_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_15_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_15_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__9016),
            .in2(_gnd_net_),
            .in3(N__8870),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__10788),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_15_8_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_15_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_15_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__9517),
            .in2(_gnd_net_),
            .in3(N__8867),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__10788),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_15_8_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_15_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_15_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(N__9433),
            .in2(_gnd_net_),
            .in3(N__8864),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__10788),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_15_8_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_15_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_15_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(N__9028),
            .in2(_gnd_net_),
            .in3(N__8861),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__10788),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_15_8_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_15_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(N__9946),
            .in2(_gnd_net_),
            .in3(N__8858),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_15_8_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_15_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_15_8_6  (
            .in0(_gnd_net_),
            .in1(N__9805),
            .in2(_gnd_net_),
            .in3(N__9035),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_15_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_15_8_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(N__9389),
            .in2(_gnd_net_),
            .in3(N__9032),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10788),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_15_9_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_15_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_15_9_0 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_15_9_0  (
            .in0(N__8986),
            .in1(N__9632),
            .in2(N__10402),
            .in3(N__9827),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_15_9_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_15_9_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_15_9_2  (
            .in0(N__9029),
            .in1(N__9017),
            .in2(N__9005),
            .in3(N__9806),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_15_9_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_15_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_15_9_3  (
            .in0(N__9965),
            .in1(N__9680),
            .in2(N__9452),
            .in3(N__9947),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_15_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_15_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_15_9_7 .LUT_INIT=16'b0100000011001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_15_9_7  (
            .in0(N__8985),
            .in1(N__10361),
            .in2(N__9668),
            .in3(N__9818),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_15_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_15_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_15_10_1 .LUT_INIT=16'b0100111001001100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_15_10_1  (
            .in0(N__9661),
            .in1(N__8965),
            .in2(N__8987),
            .in3(N__9836),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__10125));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_15_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_15_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_15_10_2 .LUT_INIT=16'b0011001100100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_15_10_2  (
            .in0(N__8951),
            .in1(N__9274),
            .in2(N__9175),
            .in3(N__8924),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__10125));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_15_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_15_10_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_15_10_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_15_10_6  (
            .in0(N__8902),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_TACK_ENC_net ),
            .ce(),
            .sr(N__10125));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_15_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_15_11_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_15_11_2 .LUT_INIT=16'b0000111101110000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_15_11_2  (
            .in0(N__9237),
            .in1(N__9205),
            .in2(N__9275),
            .in3(N__9302),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__10123));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_15_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_15_11_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_15_11_3 .LUT_INIT=16'b0011111110000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_15_11_3  (
            .in0(N__9304),
            .in1(N__9273),
            .in2(N__9215),
            .in3(N__9239),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__10123));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_15_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_15_11_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_15_11_7 .LUT_INIT=16'b0011100001111000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_15_11_7  (
            .in0(N__9303),
            .in1(N__9272),
            .in2(N__9214),
            .in3(N__9238),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net ),
            .ce(),
            .sr(N__10123));
    defparam \U409_TRANSFER_ACK.TACK_EN_RNIPUKQ5_LC_15_16_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNIPUKQ5_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_RNIPUKQ5_LC_15_16_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_RNIPUKQ5_LC_15_16_4  (
            .in0(N__9176),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9112),
            .lcout(TCIn_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_16_6_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_16_6_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_16_6_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_16_6_0  (
            .in0(N__9338),
            .in1(N__9588),
            .in2(N__10604),
            .in3(N__9625),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10787),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_16_6_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_16_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_16_6_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_16_6_1  (
            .in0(N__10065),
            .in1(_gnd_net_),
            .in2(N__10091),
            .in3(_gnd_net_),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10787),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_16_6_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_16_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_16_6_2 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_16_6_2  (
            .in0(N__9336),
            .in1(N__9586),
            .in2(N__10070),
            .in3(N__9623),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10787),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_16_6_3 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_16_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_16_6_3 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \U409_TICK.TICK50_LC_16_6_3  (
            .in0(N__9585),
            .in1(N__9339),
            .in2(N__9626),
            .in3(N__9046),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10787),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_16_6_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_16_6_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_16_6_4 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_16_6_4  (
            .in0(N__9337),
            .in1(N__9587),
            .in2(N__9986),
            .in3(N__9624),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10787),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_16_6_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_16_6_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_16_6_5  (
            .in0(N__10043),
            .in1(N__10574),
            .in2(N__10090),
            .in3(N__10804),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_16_6_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_16_6_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_16_6_6  (
            .in0(N__10028),
            .in1(N__9998),
            .in2(_gnd_net_),
            .in3(N__10064),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_16_6_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_16_6_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_16_6_7  (
            .in0(N__9353),
            .in1(N__10499),
            .in2(N__9347),
            .in3(N__10535),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_16_7_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_16_7_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_16_7_0  (
            .in0(N__10013),
            .in1(N__10853),
            .in2(N__10592),
            .in3(N__10829),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_16_7_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_16_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_16_7_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_16_7_1  (
            .in0(N__9328),
            .in1(N__9590),
            .in2(N__9344),
            .in3(N__10508),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10789),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_16_7_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_16_7_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_16_7_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_16_7_2  (
            .in0(N__9589),
            .in1(N__9619),
            .in2(N__10841),
            .in3(N__9335),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10789),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_16_7_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_16_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_16_7_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_16_7_3  (
            .in0(N__9617),
            .in1(N__9592),
            .in2(N__9340),
            .in3(N__10817),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10789),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_16_7_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_16_7_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_16_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(N__9483),
            .in2(_gnd_net_),
            .in3(N__9409),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10789),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_16_7_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_16_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_16_7_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_16_7_5  (
            .in0(N__9618),
            .in1(N__9593),
            .in2(N__9341),
            .in3(N__10544),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10789),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_16_7_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_16_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_16_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_16_7_6  (
            .in0(N__10520),
            .in1(N__10556),
            .in2(N__10619),
            .in3(N__10484),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_16_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_16_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_16_7_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_16_7_7  (
            .in0(N__9616),
            .in1(N__9591),
            .in2(N__9560),
            .in3(N__10472),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10789),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_16_8_0 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_16_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_16_8_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \U409_TICK.TICK60_LC_16_8_0  (
            .in0(N__9714),
            .in1(N__9790),
            .in2(N__9767),
            .in3(N__9544),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10791),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_16_8_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_16_8_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_16_8_1  (
            .in0(N__9533),
            .in1(N__9365),
            .in2(_gnd_net_),
            .in3(N__9482),
            .lcout(),
            .ltout(\U409_TICK.TICK603_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_16_8_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_16_8_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_16_8_2  (
            .in0(N__9377),
            .in1(N__9521),
            .in2(N__9506),
            .in3(N__9503),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_16_8_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_16_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_16_8_3 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_16_8_3  (
            .in0(N__9488),
            .in1(N__9753),
            .in2(N__9491),
            .in3(N__9716),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10791),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_16_8_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_16_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_16_8_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_16_8_4  (
            .in0(N__9713),
            .in1(N__9789),
            .in2(N__9766),
            .in3(N__9458),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10791),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_16_8_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_16_8_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_16_8_5  (
            .in0(N__9434),
            .in1(N__9422),
            .in2(N__9410),
            .in3(N__9388),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_16_8_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_16_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_16_8_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_16_8_6  (
            .in0(N__9712),
            .in1(N__9788),
            .in2(N__9765),
            .in3(N__9371),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10791),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_16_8_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_16_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_16_8_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_16_8_7  (
            .in0(N__9791),
            .in1(N__9715),
            .in2(N__9974),
            .in3(N__9763),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10791),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_16_9_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_16_9_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_16_9_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_16_9_0  (
            .in0(N__9792),
            .in1(N__9748),
            .in2(N__9724),
            .in3(N__9953),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10793),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_16_9_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_16_9_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_16_9_1  (
            .in0(N__9932),
            .in1(N__10447),
            .in2(_gnd_net_),
            .in3(N__10462),
            .lcout(\U409_TRANSFER_ACK.N_17_mux ),
            .ltout(\U409_TRANSFER_ACK.N_17_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_16_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_16_9_2 .LUT_INIT=16'b0001101101011111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_16_9_2  (
            .in0(N__9660),
            .in1(N__10434),
            .in2(N__9830),
            .in3(N__10145),
            .lcout(\U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_16_9_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_16_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__10448),
            .in2(_gnd_net_),
            .in3(N__10461),
            .lcout(\U409_TRANSFER_ACK.N_3_0 ),
            .ltout(\U409_TRANSFER_ACK.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_16_9_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_16_9_4 .LUT_INIT=16'b0000010100100111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_16_9_4  (
            .in0(N__9659),
            .in1(N__10435),
            .in2(N__9821),
            .in3(N__10146),
            .lcout(\U409_TRANSFER_ACK.N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_16_9_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_16_9_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_16_9_5 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_16_9_5  (
            .in0(N__9812),
            .in1(N__9720),
            .in2(N__9764),
            .in3(N__9794),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10793),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_16_9_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_16_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_16_9_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_16_9_6  (
            .in0(N__9793),
            .in1(N__9749),
            .in2(N__9725),
            .in3(N__9686),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10793),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_16_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_16_9_7 .LUT_INIT=16'b0011011100000100;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_16_9_7  (
            .in0(N__10147),
            .in1(N__9658),
            .in2(N__10439),
            .in3(N__9638),
            .lcout(\U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_16_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_16_10_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_16_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10463),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(N__10126));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_16_10_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_16_10_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_16_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10148),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(N__10126));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_16_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_16_10_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_16_10_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_16_10_7  (
            .in0(N__10398),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10171),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.LASTCLK_1C_net ),
            .ce(),
            .sr(N__10126));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_17_6_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_17_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_17_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_17_6_0  (
            .in0(_gnd_net_),
            .in1(N__10083),
            .in2(N__10069),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_6_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_17_6_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_17_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_17_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_17_6_1  (
            .in0(_gnd_net_),
            .in1(N__10042),
            .in2(_gnd_net_),
            .in3(N__10031),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__10790),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_17_6_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_17_6_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_17_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_17_6_2  (
            .in0(_gnd_net_),
            .in1(N__10027),
            .in2(_gnd_net_),
            .in3(N__10016),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__10790),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_17_6_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_17_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_17_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_17_6_3  (
            .in0(_gnd_net_),
            .in1(N__10012),
            .in2(_gnd_net_),
            .in3(N__10001),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__10790),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_17_6_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_17_6_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_17_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_17_6_4  (
            .in0(_gnd_net_),
            .in1(N__9997),
            .in2(_gnd_net_),
            .in3(N__9977),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_17_6_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_17_6_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_17_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_17_6_5  (
            .in0(_gnd_net_),
            .in1(N__10615),
            .in2(_gnd_net_),
            .in3(N__10595),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_17_6_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_17_6_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_17_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_17_6_6  (
            .in0(_gnd_net_),
            .in1(N__10588),
            .in2(_gnd_net_),
            .in3(N__10577),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__10790),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_17_6_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_17_6_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_17_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_17_6_7  (
            .in0(_gnd_net_),
            .in1(N__10570),
            .in2(_gnd_net_),
            .in3(N__10559),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__10790),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_17_7_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_17_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_17_7_0  (
            .in0(_gnd_net_),
            .in1(N__10555),
            .in2(_gnd_net_),
            .in3(N__10538),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_17_7_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_17_7_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_17_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_17_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_17_7_1  (
            .in0(_gnd_net_),
            .in1(N__10534),
            .in2(_gnd_net_),
            .in3(N__10523),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__10792),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_17_7_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_17_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_17_7_2  (
            .in0(_gnd_net_),
            .in1(N__10519),
            .in2(_gnd_net_),
            .in3(N__10502),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_17_7_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_17_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_17_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_17_7_3  (
            .in0(_gnd_net_),
            .in1(N__10498),
            .in2(_gnd_net_),
            .in3(N__10487),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__10792),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_17_7_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_17_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_17_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_17_7_4  (
            .in0(_gnd_net_),
            .in1(N__10483),
            .in2(_gnd_net_),
            .in3(N__10466),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_17_7_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_17_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_17_7_5  (
            .in0(_gnd_net_),
            .in1(N__10852),
            .in2(_gnd_net_),
            .in3(N__10832),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_17_7_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_17_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_17_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_17_7_6  (
            .in0(_gnd_net_),
            .in1(N__10828),
            .in2(_gnd_net_),
            .in3(N__10811),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_17_7_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_17_7_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_17_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_17_7_7  (
            .in0(_gnd_net_),
            .in1(N__10805),
            .in2(_gnd_net_),
            .in3(N__10808),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10792),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_18_12_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_18_12_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_18_12_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_18_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_0_LC_23_9_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_0_LC_23_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_0_LC_23_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_0_LC_23_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10727),
            .lcout(U409_ADDRESS_DECODE_un1_ATA_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PCS1_LC_24_2_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PCS1_LC_24_2_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PCS1_LC_24_2_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.PCS1_LC_24_2_3  (
            .in0(N__10955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10676),
            .lcout(PCS1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PCS0_LC_24_3_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PCS0_LC_24_3_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PCS0_LC_24_3_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U409_ADDRESS_DECODE.PCS0_LC_24_3_1  (
            .in0(_gnd_net_),
            .in1(N__10672),
            .in2(_gnd_net_),
            .in3(N__10956),
            .lcout(PCS0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.SCS0_LC_24_3_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.SCS0_LC_24_3_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.SCS0_LC_24_3_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U409_ADDRESS_DECODE.SCS0_LC_24_3_5  (
            .in0(N__10975),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10957),
            .lcout(SCS0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.SCS1_LC_24_3_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.SCS1_LC_24_3_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.SCS1_LC_24_3_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.SCS1_LC_24_3_7  (
            .in0(N__10976),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10958),
            .lcout(SCS1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam AGNUS_CLK_obuf_RNO_LC_24_14_6.C_ON=1'b0;
    defparam AGNUS_CLK_obuf_RNO_LC_24_14_6.SEQ_MODE=4'b0000;
    defparam AGNUS_CLK_obuf_RNO_LC_24_14_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 AGNUS_CLK_obuf_RNO_LC_24_14_6 (
            .in0(N__10916),
            .in1(N__10889),
            .in2(_gnd_net_),
            .in3(N__10877),
            .lcout(AGNUS_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 28 2025 13:13:51

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    DRA,
    CMA,
    DA,
    A,
    DBRn,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    TCIn,
    TBIn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    input [9:0] DRA;
    output [10:0] CMA;
    output [2:0] DA;
    input [20:0] A;
    input DBRn;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    output TCIn;
    output TBIn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__12519;
    wire N__12518;
    wire N__12517;
    wire N__12510;
    wire N__12509;
    wire N__12508;
    wire N__12501;
    wire N__12500;
    wire N__12499;
    wire N__12492;
    wire N__12491;
    wire N__12490;
    wire N__12483;
    wire N__12482;
    wire N__12481;
    wire N__12474;
    wire N__12473;
    wire N__12472;
    wire N__12465;
    wire N__12464;
    wire N__12463;
    wire N__12456;
    wire N__12455;
    wire N__12454;
    wire N__12447;
    wire N__12446;
    wire N__12445;
    wire N__12438;
    wire N__12437;
    wire N__12436;
    wire N__12429;
    wire N__12428;
    wire N__12427;
    wire N__12420;
    wire N__12419;
    wire N__12418;
    wire N__12411;
    wire N__12410;
    wire N__12409;
    wire N__12402;
    wire N__12401;
    wire N__12400;
    wire N__12393;
    wire N__12392;
    wire N__12391;
    wire N__12384;
    wire N__12383;
    wire N__12382;
    wire N__12375;
    wire N__12374;
    wire N__12373;
    wire N__12366;
    wire N__12365;
    wire N__12364;
    wire N__12357;
    wire N__12356;
    wire N__12355;
    wire N__12348;
    wire N__12347;
    wire N__12346;
    wire N__12339;
    wire N__12338;
    wire N__12337;
    wire N__12330;
    wire N__12329;
    wire N__12328;
    wire N__12321;
    wire N__12320;
    wire N__12319;
    wire N__12312;
    wire N__12311;
    wire N__12310;
    wire N__12303;
    wire N__12302;
    wire N__12301;
    wire N__12294;
    wire N__12293;
    wire N__12292;
    wire N__12285;
    wire N__12284;
    wire N__12283;
    wire N__12276;
    wire N__12275;
    wire N__12274;
    wire N__12267;
    wire N__12266;
    wire N__12265;
    wire N__12258;
    wire N__12257;
    wire N__12256;
    wire N__12249;
    wire N__12248;
    wire N__12247;
    wire N__12240;
    wire N__12239;
    wire N__12238;
    wire N__12231;
    wire N__12230;
    wire N__12229;
    wire N__12222;
    wire N__12221;
    wire N__12220;
    wire N__12213;
    wire N__12212;
    wire N__12211;
    wire N__12204;
    wire N__12203;
    wire N__12202;
    wire N__12195;
    wire N__12194;
    wire N__12193;
    wire N__12186;
    wire N__12185;
    wire N__12184;
    wire N__12177;
    wire N__12176;
    wire N__12175;
    wire N__12168;
    wire N__12167;
    wire N__12166;
    wire N__12159;
    wire N__12158;
    wire N__12157;
    wire N__12150;
    wire N__12149;
    wire N__12148;
    wire N__12141;
    wire N__12140;
    wire N__12139;
    wire N__12132;
    wire N__12131;
    wire N__12130;
    wire N__12123;
    wire N__12122;
    wire N__12121;
    wire N__12114;
    wire N__12113;
    wire N__12112;
    wire N__12105;
    wire N__12104;
    wire N__12103;
    wire N__12096;
    wire N__12095;
    wire N__12094;
    wire N__12087;
    wire N__12086;
    wire N__12085;
    wire N__12078;
    wire N__12077;
    wire N__12076;
    wire N__12069;
    wire N__12068;
    wire N__12067;
    wire N__12060;
    wire N__12059;
    wire N__12058;
    wire N__12051;
    wire N__12050;
    wire N__12049;
    wire N__12042;
    wire N__12041;
    wire N__12040;
    wire N__12033;
    wire N__12032;
    wire N__12031;
    wire N__12024;
    wire N__12023;
    wire N__12022;
    wire N__12015;
    wire N__12014;
    wire N__12013;
    wire N__12006;
    wire N__12005;
    wire N__12004;
    wire N__11997;
    wire N__11996;
    wire N__11995;
    wire N__11988;
    wire N__11987;
    wire N__11986;
    wire N__11979;
    wire N__11978;
    wire N__11977;
    wire N__11970;
    wire N__11969;
    wire N__11968;
    wire N__11961;
    wire N__11960;
    wire N__11959;
    wire N__11952;
    wire N__11951;
    wire N__11950;
    wire N__11943;
    wire N__11942;
    wire N__11941;
    wire N__11934;
    wire N__11933;
    wire N__11932;
    wire N__11925;
    wire N__11924;
    wire N__11923;
    wire N__11916;
    wire N__11915;
    wire N__11914;
    wire N__11907;
    wire N__11906;
    wire N__11905;
    wire N__11898;
    wire N__11897;
    wire N__11896;
    wire N__11889;
    wire N__11888;
    wire N__11887;
    wire N__11880;
    wire N__11879;
    wire N__11878;
    wire N__11871;
    wire N__11870;
    wire N__11869;
    wire N__11862;
    wire N__11861;
    wire N__11860;
    wire N__11853;
    wire N__11852;
    wire N__11851;
    wire N__11844;
    wire N__11843;
    wire N__11842;
    wire N__11835;
    wire N__11834;
    wire N__11833;
    wire N__11826;
    wire N__11825;
    wire N__11824;
    wire N__11817;
    wire N__11816;
    wire N__11815;
    wire N__11808;
    wire N__11807;
    wire N__11806;
    wire N__11799;
    wire N__11798;
    wire N__11797;
    wire N__11790;
    wire N__11789;
    wire N__11788;
    wire N__11781;
    wire N__11780;
    wire N__11779;
    wire N__11772;
    wire N__11771;
    wire N__11770;
    wire N__11763;
    wire N__11762;
    wire N__11761;
    wire N__11754;
    wire N__11753;
    wire N__11752;
    wire N__11745;
    wire N__11744;
    wire N__11743;
    wire N__11736;
    wire N__11735;
    wire N__11734;
    wire N__11727;
    wire N__11726;
    wire N__11725;
    wire N__11718;
    wire N__11717;
    wire N__11716;
    wire N__11709;
    wire N__11708;
    wire N__11707;
    wire N__11700;
    wire N__11699;
    wire N__11698;
    wire N__11691;
    wire N__11690;
    wire N__11689;
    wire N__11682;
    wire N__11681;
    wire N__11680;
    wire N__11673;
    wire N__11672;
    wire N__11671;
    wire N__11654;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11644;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11625;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11594;
    wire N__11593;
    wire N__11590;
    wire N__11589;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11579;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11552;
    wire N__11549;
    wire N__11548;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11523;
    wire N__11522;
    wire N__11517;
    wire N__11514;
    wire N__11511;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11480;
    wire N__11477;
    wire N__11474;
    wire N__11471;
    wire N__11468;
    wire N__11465;
    wire N__11462;
    wire N__11459;
    wire N__11456;
    wire N__11455;
    wire N__11452;
    wire N__11451;
    wire N__11448;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11435;
    wire N__11430;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11416;
    wire N__11411;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11395;
    wire N__11394;
    wire N__11393;
    wire N__11390;
    wire N__11387;
    wire N__11382;
    wire N__11379;
    wire N__11374;
    wire N__11369;
    wire N__11366;
    wire N__11365;
    wire N__11362;
    wire N__11359;
    wire N__11358;
    wire N__11353;
    wire N__11352;
    wire N__11349;
    wire N__11346;
    wire N__11343;
    wire N__11340;
    wire N__11337;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11323;
    wire N__11318;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11293;
    wire N__11292;
    wire N__11291;
    wire N__11290;
    wire N__11289;
    wire N__11288;
    wire N__11287;
    wire N__11286;
    wire N__11285;
    wire N__11284;
    wire N__11283;
    wire N__11282;
    wire N__11281;
    wire N__11280;
    wire N__11279;
    wire N__11276;
    wire N__11275;
    wire N__11274;
    wire N__11269;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11234;
    wire N__11233;
    wire N__11230;
    wire N__11229;
    wire N__11226;
    wire N__11223;
    wire N__11220;
    wire N__11217;
    wire N__11210;
    wire N__11207;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11182;
    wire N__11171;
    wire N__11166;
    wire N__11161;
    wire N__11158;
    wire N__11151;
    wire N__11148;
    wire N__11143;
    wire N__11140;
    wire N__11137;
    wire N__11132;
    wire N__11131;
    wire N__11128;
    wire N__11125;
    wire N__11124;
    wire N__11123;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11089;
    wire N__11086;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11068;
    wire N__11067;
    wire N__11066;
    wire N__11065;
    wire N__11064;
    wire N__11063;
    wire N__11062;
    wire N__11061;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11035;
    wire N__11034;
    wire N__11033;
    wire N__11032;
    wire N__11031;
    wire N__11030;
    wire N__11029;
    wire N__11028;
    wire N__11027;
    wire N__11026;
    wire N__11025;
    wire N__11024;
    wire N__11023;
    wire N__11022;
    wire N__11021;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10981;
    wire N__10980;
    wire N__10979;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10966;
    wire N__10965;
    wire N__10964;
    wire N__10963;
    wire N__10962;
    wire N__10959;
    wire N__10958;
    wire N__10957;
    wire N__10956;
    wire N__10955;
    wire N__10954;
    wire N__10953;
    wire N__10952;
    wire N__10951;
    wire N__10950;
    wire N__10949;
    wire N__10948;
    wire N__10947;
    wire N__10946;
    wire N__10945;
    wire N__10944;
    wire N__10943;
    wire N__10942;
    wire N__10941;
    wire N__10940;
    wire N__10939;
    wire N__10938;
    wire N__10935;
    wire N__10934;
    wire N__10933;
    wire N__10932;
    wire N__10931;
    wire N__10930;
    wire N__10929;
    wire N__10928;
    wire N__10927;
    wire N__10926;
    wire N__10925;
    wire N__10924;
    wire N__10923;
    wire N__10922;
    wire N__10919;
    wire N__10918;
    wire N__10917;
    wire N__10914;
    wire N__10913;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10806;
    wire N__10805;
    wire N__10802;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10789;
    wire N__10786;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10761;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10726;
    wire N__10725;
    wire N__10724;
    wire N__10723;
    wire N__10722;
    wire N__10721;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10700;
    wire N__10697;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10666;
    wire N__10665;
    wire N__10662;
    wire N__10661;
    wire N__10656;
    wire N__10653;
    wire N__10650;
    wire N__10647;
    wire N__10644;
    wire N__10641;
    wire N__10638;
    wire N__10637;
    wire N__10636;
    wire N__10633;
    wire N__10630;
    wire N__10627;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10611;
    wire N__10608;
    wire N__10603;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10588;
    wire N__10585;
    wire N__10584;
    wire N__10581;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10562;
    wire N__10559;
    wire N__10558;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10524;
    wire N__10521;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10465;
    wire N__10464;
    wire N__10457;
    wire N__10456;
    wire N__10455;
    wire N__10454;
    wire N__10451;
    wire N__10444;
    wire N__10439;
    wire N__10438;
    wire N__10437;
    wire N__10436;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10412;
    wire N__10411;
    wire N__10408;
    wire N__10403;
    wire N__10400;
    wire N__10399;
    wire N__10398;
    wire N__10395;
    wire N__10390;
    wire N__10387;
    wire N__10384;
    wire N__10379;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10339;
    wire N__10338;
    wire N__10337;
    wire N__10336;
    wire N__10335;
    wire N__10334;
    wire N__10333;
    wire N__10332;
    wire N__10331;
    wire N__10330;
    wire N__10329;
    wire N__10328;
    wire N__10327;
    wire N__10326;
    wire N__10325;
    wire N__10324;
    wire N__10323;
    wire N__10322;
    wire N__10321;
    wire N__10320;
    wire N__10319;
    wire N__10318;
    wire N__10317;
    wire N__10316;
    wire N__10315;
    wire N__10314;
    wire N__10313;
    wire N__10312;
    wire N__10311;
    wire N__10310;
    wire N__10309;
    wire N__10308;
    wire N__10307;
    wire N__10306;
    wire N__10305;
    wire N__10304;
    wire N__10301;
    wire N__10300;
    wire N__10299;
    wire N__10298;
    wire N__10297;
    wire N__10296;
    wire N__10295;
    wire N__10294;
    wire N__10293;
    wire N__10202;
    wire N__10199;
    wire N__10198;
    wire N__10197;
    wire N__10194;
    wire N__10191;
    wire N__10190;
    wire N__10187;
    wire N__10182;
    wire N__10179;
    wire N__10178;
    wire N__10177;
    wire N__10174;
    wire N__10171;
    wire N__10168;
    wire N__10165;
    wire N__10162;
    wire N__10159;
    wire N__10152;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10133;
    wire N__10132;
    wire N__10131;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10111;
    wire N__10108;
    wire N__10105;
    wire N__10102;
    wire N__10099;
    wire N__10096;
    wire N__10093;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10081;
    wire N__10080;
    wire N__10079;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10060;
    wire N__10057;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10045;
    wire N__10044;
    wire N__10043;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9868;
    wire N__9865;
    wire N__9864;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9856;
    wire N__9853;
    wire N__9850;
    wire N__9847;
    wire N__9844;
    wire N__9843;
    wire N__9840;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9788;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9776;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9768;
    wire N__9767;
    wire N__9762;
    wire N__9759;
    wire N__9758;
    wire N__9757;
    wire N__9756;
    wire N__9753;
    wire N__9750;
    wire N__9747;
    wire N__9744;
    wire N__9741;
    wire N__9738;
    wire N__9735;
    wire N__9730;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9706;
    wire N__9705;
    wire N__9704;
    wire N__9703;
    wire N__9700;
    wire N__9699;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9691;
    wire N__9690;
    wire N__9687;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9670;
    wire N__9669;
    wire N__9664;
    wire N__9661;
    wire N__9660;
    wire N__9659;
    wire N__9652;
    wire N__9647;
    wire N__9644;
    wire N__9643;
    wire N__9642;
    wire N__9641;
    wire N__9638;
    wire N__9633;
    wire N__9630;
    wire N__9629;
    wire N__9628;
    wire N__9627;
    wire N__9626;
    wire N__9625;
    wire N__9624;
    wire N__9617;
    wire N__9612;
    wire N__9609;
    wire N__9602;
    wire N__9597;
    wire N__9594;
    wire N__9589;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9571;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9541;
    wire N__9538;
    wire N__9535;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9523;
    wire N__9518;
    wire N__9515;
    wire N__9514;
    wire N__9511;
    wire N__9508;
    wire N__9505;
    wire N__9500;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9490;
    wire N__9487;
    wire N__9486;
    wire N__9485;
    wire N__9480;
    wire N__9477;
    wire N__9474;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9436;
    wire N__9433;
    wire N__9430;
    wire N__9429;
    wire N__9424;
    wire N__9421;
    wire N__9420;
    wire N__9417;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9344;
    wire N__9343;
    wire N__9342;
    wire N__9341;
    wire N__9340;
    wire N__9339;
    wire N__9338;
    wire N__9337;
    wire N__9334;
    wire N__9333;
    wire N__9332;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9314;
    wire N__9313;
    wire N__9310;
    wire N__9309;
    wire N__9308;
    wire N__9307;
    wire N__9306;
    wire N__9305;
    wire N__9304;
    wire N__9303;
    wire N__9300;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9288;
    wire N__9285;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9265;
    wire N__9258;
    wire N__9251;
    wire N__9250;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9225;
    wire N__9222;
    wire N__9219;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9194;
    wire N__9187;
    wire N__9184;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9043;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8992;
    wire N__8991;
    wire N__8988;
    wire N__8983;
    wire N__8980;
    wire N__8977;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8875;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8863;
    wire N__8860;
    wire N__8857;
    wire N__8854;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8806;
    wire N__8801;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8779;
    wire N__8776;
    wire N__8773;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8761;
    wire N__8758;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8719;
    wire N__8718;
    wire N__8715;
    wire N__8710;
    wire N__8707;
    wire N__8704;
    wire N__8703;
    wire N__8700;
    wire N__8697;
    wire N__8694;
    wire N__8687;
    wire N__8686;
    wire N__8683;
    wire N__8680;
    wire N__8679;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8667;
    wire N__8664;
    wire N__8661;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8515;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8501;
    wire N__8500;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8476;
    wire N__8475;
    wire N__8474;
    wire N__8473;
    wire N__8472;
    wire N__8471;
    wire N__8468;
    wire N__8467;
    wire N__8466;
    wire N__8465;
    wire N__8460;
    wire N__8459;
    wire N__8458;
    wire N__8457;
    wire N__8454;
    wire N__8449;
    wire N__8448;
    wire N__8445;
    wire N__8442;
    wire N__8439;
    wire N__8436;
    wire N__8433;
    wire N__8430;
    wire N__8425;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8377;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8362;
    wire N__8357;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8338;
    wire N__8337;
    wire N__8334;
    wire N__8331;
    wire N__8330;
    wire N__8329;
    wire N__8328;
    wire N__8327;
    wire N__8326;
    wire N__8323;
    wire N__8322;
    wire N__8321;
    wire N__8320;
    wire N__8319;
    wire N__8318;
    wire N__8315;
    wire N__8312;
    wire N__8307;
    wire N__8304;
    wire N__8303;
    wire N__8302;
    wire N__8301;
    wire N__8298;
    wire N__8297;
    wire N__8294;
    wire N__8291;
    wire N__8286;
    wire N__8279;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8257;
    wire N__8240;
    wire N__8239;
    wire N__8238;
    wire N__8235;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8227;
    wire N__8226;
    wire N__8225;
    wire N__8224;
    wire N__8221;
    wire N__8220;
    wire N__8219;
    wire N__8216;
    wire N__8215;
    wire N__8214;
    wire N__8213;
    wire N__8212;
    wire N__8209;
    wire N__8204;
    wire N__8201;
    wire N__8200;
    wire N__8199;
    wire N__8198;
    wire N__8197;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8187;
    wire N__8184;
    wire N__8181;
    wire N__8176;
    wire N__8169;
    wire N__8162;
    wire N__8159;
    wire N__8154;
    wire N__8149;
    wire N__8126;
    wire N__8125;
    wire N__8122;
    wire N__8121;
    wire N__8118;
    wire N__8117;
    wire N__8114;
    wire N__8113;
    wire N__8112;
    wire N__8109;
    wire N__8108;
    wire N__8103;
    wire N__8100;
    wire N__8093;
    wire N__8092;
    wire N__8091;
    wire N__8090;
    wire N__8089;
    wire N__8088;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8076;
    wire N__8073;
    wire N__8070;
    wire N__8063;
    wire N__8060;
    wire N__8045;
    wire N__8044;
    wire N__8043;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8035;
    wire N__8034;
    wire N__8031;
    wire N__8030;
    wire N__8029;
    wire N__8028;
    wire N__8027;
    wire N__8026;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8015;
    wire N__8012;
    wire N__8011;
    wire N__8010;
    wire N__8009;
    wire N__8006;
    wire N__8001;
    wire N__7998;
    wire N__7995;
    wire N__7988;
    wire N__7981;
    wire N__7978;
    wire N__7977;
    wire N__7974;
    wire N__7973;
    wire N__7970;
    wire N__7969;
    wire N__7968;
    wire N__7965;
    wire N__7962;
    wire N__7959;
    wire N__7956;
    wire N__7945;
    wire N__7944;
    wire N__7943;
    wire N__7942;
    wire N__7939;
    wire N__7936;
    wire N__7933;
    wire N__7930;
    wire N__7927;
    wire N__7922;
    wire N__7919;
    wire N__7912;
    wire N__7905;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7879;
    wire N__7878;
    wire N__7877;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7863;
    wire N__7860;
    wire N__7855;
    wire N__7854;
    wire N__7853;
    wire N__7852;
    wire N__7851;
    wire N__7850;
    wire N__7849;
    wire N__7848;
    wire N__7847;
    wire N__7846;
    wire N__7845;
    wire N__7840;
    wire N__7837;
    wire N__7834;
    wire N__7829;
    wire N__7826;
    wire N__7821;
    wire N__7820;
    wire N__7813;
    wire N__7812;
    wire N__7807;
    wire N__7806;
    wire N__7805;
    wire N__7804;
    wire N__7803;
    wire N__7798;
    wire N__7793;
    wire N__7792;
    wire N__7791;
    wire N__7790;
    wire N__7787;
    wire N__7786;
    wire N__7785;
    wire N__7784;
    wire N__7783;
    wire N__7782;
    wire N__7779;
    wire N__7776;
    wire N__7773;
    wire N__7766;
    wire N__7763;
    wire N__7762;
    wire N__7761;
    wire N__7756;
    wire N__7751;
    wire N__7746;
    wire N__7739;
    wire N__7734;
    wire N__7731;
    wire N__7722;
    wire N__7717;
    wire N__7706;
    wire N__7699;
    wire N__7696;
    wire N__7693;
    wire N__7688;
    wire N__7685;
    wire N__7682;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7657;
    wire N__7656;
    wire N__7653;
    wire N__7650;
    wire N__7647;
    wire N__7640;
    wire N__7637;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7619;
    wire N__7618;
    wire N__7617;
    wire N__7616;
    wire N__7615;
    wire N__7614;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7602;
    wire N__7597;
    wire N__7594;
    wire N__7583;
    wire N__7580;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7570;
    wire N__7565;
    wire N__7564;
    wire N__7561;
    wire N__7560;
    wire N__7559;
    wire N__7558;
    wire N__7555;
    wire N__7554;
    wire N__7551;
    wire N__7548;
    wire N__7547;
    wire N__7546;
    wire N__7545;
    wire N__7544;
    wire N__7543;
    wire N__7542;
    wire N__7541;
    wire N__7538;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7525;
    wire N__7522;
    wire N__7517;
    wire N__7508;
    wire N__7505;
    wire N__7500;
    wire N__7481;
    wire N__7480;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7427;
    wire N__7424;
    wire N__7421;
    wire N__7418;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7397;
    wire N__7396;
    wire N__7395;
    wire N__7394;
    wire N__7391;
    wire N__7388;
    wire N__7387;
    wire N__7384;
    wire N__7381;
    wire N__7380;
    wire N__7379;
    wire N__7376;
    wire N__7375;
    wire N__7374;
    wire N__7371;
    wire N__7368;
    wire N__7365;
    wire N__7362;
    wire N__7359;
    wire N__7356;
    wire N__7353;
    wire N__7348;
    wire N__7343;
    wire N__7334;
    wire N__7325;
    wire N__7322;
    wire N__7321;
    wire N__7318;
    wire N__7315;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7301;
    wire N__7300;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7290;
    wire N__7283;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7270;
    wire N__7269;
    wire N__7268;
    wire N__7267;
    wire N__7264;
    wire N__7261;
    wire N__7258;
    wire N__7257;
    wire N__7252;
    wire N__7249;
    wire N__7248;
    wire N__7247;
    wire N__7244;
    wire N__7241;
    wire N__7238;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7220;
    wire N__7217;
    wire N__7208;
    wire N__7205;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7197;
    wire N__7196;
    wire N__7193;
    wire N__7190;
    wire N__7187;
    wire N__7184;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7166;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7147;
    wire N__7146;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7124;
    wire N__7121;
    wire N__7120;
    wire N__7119;
    wire N__7118;
    wire N__7115;
    wire N__7110;
    wire N__7107;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7090;
    wire N__7085;
    wire N__7084;
    wire N__7081;
    wire N__7080;
    wire N__7077;
    wire N__7074;
    wire N__7071;
    wire N__7064;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7012;
    wire N__7011;
    wire N__7010;
    wire N__7009;
    wire N__7008;
    wire N__7003;
    wire N__7002;
    wire N__6999;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6983;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6971;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6957;
    wire N__6954;
    wire N__6951;
    wire N__6948;
    wire N__6943;
    wire N__6940;
    wire N__6935;
    wire N__6934;
    wire N__6933;
    wire N__6932;
    wire N__6931;
    wire N__6930;
    wire N__6923;
    wire N__6920;
    wire N__6915;
    wire N__6908;
    wire N__6905;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6895;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6885;
    wire N__6880;
    wire N__6877;
    wire N__6876;
    wire N__6875;
    wire N__6870;
    wire N__6867;
    wire N__6864;
    wire N__6863;
    wire N__6862;
    wire N__6859;
    wire N__6852;
    wire N__6849;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6827;
    wire N__6824;
    wire N__6823;
    wire N__6822;
    wire N__6819;
    wire N__6818;
    wire N__6817;
    wire N__6816;
    wire N__6815;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6786;
    wire N__6781;
    wire N__6778;
    wire N__6775;
    wire N__6774;
    wire N__6771;
    wire N__6768;
    wire N__6765;
    wire N__6762;
    wire N__6759;
    wire N__6756;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6710;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6614;
    wire N__6611;
    wire N__6608;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6587;
    wire N__6584;
    wire N__6583;
    wire N__6582;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6545;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6491;
    wire N__6490;
    wire N__6487;
    wire N__6484;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6455;
    wire N__6452;
    wire N__6449;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6437;
    wire N__6434;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6391;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6381;
    wire N__6374;
    wire N__6373;
    wire N__6372;
    wire N__6369;
    wire N__6366;
    wire N__6363;
    wire N__6356;
    wire N__6355;
    wire N__6354;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6332;
    wire N__6331;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6314;
    wire N__6311;
    wire N__6310;
    wire N__6307;
    wire N__6306;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6290;
    wire N__6287;
    wire N__6284;
    wire N__6283;
    wire N__6282;
    wire N__6277;
    wire N__6274;
    wire N__6273;
    wire N__6270;
    wire N__6267;
    wire N__6264;
    wire N__6259;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6220;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6198;
    wire N__6197;
    wire N__6196;
    wire N__6193;
    wire N__6190;
    wire N__6183;
    wire N__6180;
    wire N__6175;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6157;
    wire N__6154;
    wire N__6153;
    wire N__6152;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6128;
    wire N__6119;
    wire N__6118;
    wire N__6117;
    wire N__6114;
    wire N__6109;
    wire N__6104;
    wire N__6101;
    wire N__6100;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6074;
    wire N__6073;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6065;
    wire N__6062;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6048;
    wire N__6045;
    wire N__6038;
    wire N__6037;
    wire N__6036;
    wire N__6029;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6008;
    wire N__6005;
    wire N__6002;
    wire N__5999;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5953;
    wire N__5952;
    wire N__5951;
    wire N__5950;
    wire N__5949;
    wire N__5948;
    wire N__5941;
    wire N__5938;
    wire N__5931;
    wire N__5924;
    wire N__5921;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5903;
    wire N__5902;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5888;
    wire N__5885;
    wire N__5880;
    wire N__5877;
    wire N__5874;
    wire N__5871;
    wire N__5868;
    wire N__5865;
    wire N__5862;
    wire N__5859;
    wire N__5856;
    wire N__5853;
    wire N__5850;
    wire N__5843;
    wire N__5840;
    wire N__5837;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5815;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5803;
    wire N__5802;
    wire N__5799;
    wire N__5794;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5765;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5753;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5741;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5729;
    wire N__5728;
    wire N__5727;
    wire N__5726;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5705;
    wire N__5704;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5671;
    wire N__5670;
    wire N__5669;
    wire N__5666;
    wire N__5661;
    wire N__5658;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5639;
    wire N__5636;
    wire N__5633;
    wire N__5630;
    wire N__5629;
    wire N__5628;
    wire N__5627;
    wire N__5626;
    wire N__5625;
    wire N__5624;
    wire N__5623;
    wire N__5622;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5585;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5573;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5558;
    wire N__5557;
    wire N__5554;
    wire N__5551;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5533;
    wire N__5532;
    wire N__5531;
    wire N__5530;
    wire N__5527;
    wire N__5526;
    wire N__5525;
    wire N__5524;
    wire N__5523;
    wire N__5522;
    wire N__5521;
    wire N__5518;
    wire N__5517;
    wire N__5514;
    wire N__5513;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5501;
    wire N__5496;
    wire N__5489;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5474;
    wire N__5471;
    wire N__5466;
    wire N__5461;
    wire N__5458;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5323;
    wire N__5320;
    wire N__5319;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5307;
    wire N__5304;
    wire N__5301;
    wire N__5298;
    wire N__5295;
    wire N__5292;
    wire N__5289;
    wire N__5286;
    wire N__5283;
    wire N__5280;
    wire N__5277;
    wire N__5274;
    wire N__5273;
    wire N__5266;
    wire N__5263;
    wire N__5258;
    wire N__5257;
    wire N__5254;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5213;
    wire N__5206;
    wire N__5203;
    wire N__5198;
    wire N__5195;
    wire N__5194;
    wire N__5191;
    wire N__5188;
    wire N__5183;
    wire N__5182;
    wire N__5179;
    wire N__5176;
    wire N__5171;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5140;
    wire N__5137;
    wire N__5134;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5119;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5109;
    wire N__5102;
    wire N__5101;
    wire N__5098;
    wire N__5095;
    wire N__5092;
    wire N__5089;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5070;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5032;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5020;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5008;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4996;
    wire N__4991;
    wire N__4990;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4946;
    wire N__4945;
    wire N__4944;
    wire N__4939;
    wire N__4936;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4915;
    wire N__4914;
    wire N__4913;
    wire N__4912;
    wire N__4911;
    wire N__4908;
    wire N__4907;
    wire N__4904;
    wire N__4903;
    wire N__4902;
    wire N__4899;
    wire N__4898;
    wire N__4895;
    wire N__4890;
    wire N__4887;
    wire N__4886;
    wire N__4885;
    wire N__4882;
    wire N__4879;
    wire N__4872;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4855;
    wire N__4852;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4825;
    wire N__4824;
    wire N__4821;
    wire N__4820;
    wire N__4819;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4802;
    wire N__4793;
    wire N__4790;
    wire N__4789;
    wire N__4786;
    wire N__4785;
    wire N__4784;
    wire N__4783;
    wire N__4780;
    wire N__4777;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4744;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4727;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4690;
    wire N__4687;
    wire N__4684;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4615;
    wire N__4614;
    wire N__4613;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4586;
    wire N__4585;
    wire N__4582;
    wire N__4581;
    wire N__4580;
    wire N__4579;
    wire N__4576;
    wire N__4573;
    wire N__4570;
    wire N__4565;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4546;
    wire N__4543;
    wire N__4540;
    wire N__4535;
    wire N__4534;
    wire N__4531;
    wire N__4530;
    wire N__4529;
    wire N__4528;
    wire N__4525;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4502;
    wire N__4499;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4469;
    wire N__4466;
    wire N__4465;
    wire N__4462;
    wire N__4459;
    wire N__4454;
    wire N__4453;
    wire N__4450;
    wire N__4447;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4385;
    wire N__4384;
    wire N__4381;
    wire N__4378;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4342;
    wire N__4339;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire DBRn_c_i_0;
    wire CLK80_PLL_i_i;
    wire DBR_SYNCZ0Z_0;
    wire DBRn_c;
    wire REGENn_c;
    wire \U712_REG_SM.START_RSTZ0 ;
    wire \U712_REG_SM.un6_REG_CYCLE_START_cascade_ ;
    wire REGSPACEn_c;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNT_1_sqmuxa_1 ;
    wire \U712_REG_SM.N_188 ;
    wire \U712_REG_SM.WRITE_CYCLEZ0 ;
    wire \U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ;
    wire \U712_REG_SM.N_157_cascade_ ;
    wire \U712_REG_SM.N_109_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTc_0_0_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_REG_SM.REG_CYCLE_0_sqmuxa_cascade_ ;
    wire \U712_REG_SM.N_185 ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.N_109_0 ;
    wire \U712_REG_SM.N_105_0 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_1 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.N_166 ;
    wire LDSn_c;
    wire DBDIR_c;
    wire bfn_8_11_0_;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_2 ;
    wire \U712_CHIP_RAM.un2_DBR_COUNT_cry_1 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_3 ;
    wire \U712_CHIP_RAM.un2_DBR_COUNT_cry_2 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_4 ;
    wire \U712_CHIP_RAM.un2_DBR_COUNT_cry_3 ;
    wire \U712_CHIP_RAM.un2_DBR_COUNT_cry_4 ;
    wire \U712_CHIP_RAM.un2_DBR_COUNT_cry_5 ;
    wire \U712_CHIP_RAM.un2_DBR_COUNT_cry_6 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_0 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_1 ;
    wire \U712_REG_SM.N_159 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_0 ;
    wire \U712_REG_SM.N_109 ;
    wire \U712_REG_SM.N_164 ;
    wire \U712_REG_SM.N_80 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_96 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_96_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire UDSn_c;
    wire U712_BYTE_ENABLE_UDS_0;
    wire \U712_REG_SM.N_163 ;
    wire CLK40_PLL_i_i;
    wire \U712_CYCLE_TERM.N_51_cascade_ ;
    wire \U712_CHIP_RAM.BANK0_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_5 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_6 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_7 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0_cascade_ ;
    wire LATCH_CLK_c;
    wire \U712_CHIP_RAM.N_144_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_4 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_3 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire ASn_c;
    wire \U712_REG_SM.N_163_0 ;
    wire TSn_c;
    wire RAMENn_c;
    wire VBENn_c;
    wire \U712_CYCLE_TERM.N_47_0 ;
    wire TACK_EN;
    wire TACK_OUTn;
    wire bfn_10_9_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH5lto1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_START_2_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.N_9 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_ ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER33_1_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_2_cascade_ ;
    wire \U712_CHIP_RAM.N_64_cascade_ ;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER18 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_1 ;
    wire \U712_CHIP_RAM.LATCH_CLK_6 ;
    wire bfn_10_13_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_64 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire CLK40_PLL_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ1Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire CLMBEn_c;
    wire \U712_CHIP_RAM.LATCH_CLK_0_sqmuxa ;
    wire \U712_CHIP_RAM.LATCH_CLK_0_sqmuxa_cascade_ ;
    wire REG_TACK;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0_cascade_ ;
    wire AWEn_c;
    wire DBR_SYNCZ0Z_1;
    wire \U712_CHIP_RAM.N_152 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.N_108_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_a3_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_0_cascade_ ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_331_3_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER37_0_a3_1_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_7_2 ;
    wire \U712_CHIP_RAM.BANK0_7_0_cascade_ ;
    wire BANK0_c;
    wire A_c_20;
    wire \U712_CHIP_RAM.A_m_20 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ;
    wire \U712_CHIP_RAM.A_m_2_20 ;
    wire \U712_CHIP_RAM.N_94_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1_cascade_ ;
    wire \U712_CHIP_RAM.N_187 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1_1_cascade_ ;
    wire \U712_CHIP_RAM.N_155 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1 ;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ;
    wire \U712_BYTE_ENABLE.N_58 ;
    wire N_56_i;
    wire SIZ_c_0;
    wire A_c_1;
    wire A_c_0;
    wire SIZ_c_1;
    wire N_58_i;
    wire DMA_LATCH_EN_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0_0 ;
    wire A_c_8;
    wire A_c_15;
    wire A_c_16;
    wire A_c_18;
    wire A_c_13;
    wire A_c_6;
    wire \U712_CHIP_RAM.CLK_EN_5_0 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_DISABLEZ0 ;
    wire \U712_CHIP_RAM.N_95 ;
    wire \U712_CHIP_RAM.N_119 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.N_95_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_3_sqmuxa_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_3_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_7 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER38_1_0 ;
    wire \U712_CHIP_RAM.N_94 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_cascade_ ;
    wire \U712_CHIP_RAM.CPU_TACK_7_0 ;
    wire CPU_TACKm;
    wire A_c_7;
    wire A_c_14;
    wire \U712_CHIP_RAM.N_173 ;
    wire \U712_CHIP_RAM.un3_CPU_CYCLE_START ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_177 ;
    wire \U712_CHIP_RAM.N_172 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_1_sqmuxa_1_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.N_186 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER34 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER34_cascade_ ;
    wire A_c_2;
    wire A_c_9;
    wire \U712_CHIP_RAM.SDRAM_COUNTER16_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER17_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER15 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER17_0_cascade_ ;
    wire \U712_CHIP_RAM.N_33 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER19_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER17_1_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa ;
    wire \U712_CHIP_RAM.N_38_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_i_1_1 ;
    wire \U712_CHIP_RAM.N_151 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER19_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_i ;
    wire \U712_CHIP_RAM.N_331_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_29_i_a2_i_1 ;
    wire \U712_CHIP_RAM.N_61_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1 ;
    wire \U712_CHIP_RAM.N_218 ;
    wire \U712_CHIP_RAM.N_154 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_29_i_a2_i_1_0 ;
    wire RESETn_c;
    wire RESETn_c_i;
    wire UMBEn_c;
    wire \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_1_cascade_ ;
    wire CUMBEn_c;
    wire UUBEn_c;
    wire \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_1 ;
    wire CUUBEn_c;
    wire DBENn_c;
    wire DMA_CYCLEm;
    wire \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_0 ;
    wire \U712_BYTE_ENABLE.N_56 ;
    wire \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_0_cascade_ ;
    wire CLLBEn_c;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire A_c_3;
    wire \U712_CHIP_RAM.N_11_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ;
    wire A_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire A_c_5;
    wire A_c_12;
    wire A_c_4;
    wire A_c_11;
    wire CMA_c_10;
    wire A_c_17;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire CPU_CYCLEm;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire WEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_4;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire DRA_c_1;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_7;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire RAS0n_c;
    wire AGNUS_REV_c;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire RnW_c;
    wire WRITE_CYCLEm;
    wire DRDDIR_c;
    wire CASLn_c;
    wire CASUn_c;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__4259),
            .RESETB(N__5831),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__12519),
            .DIN(N__12518),
            .DOUT(N__12517),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__12519),
            .PADOUT(N__12518),
            .PADIN(N__12517),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8723),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__12510),
            .DIN(N__12509),
            .DOUT(N__12508),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__12510),
            .PADOUT(N__12509),
            .PADIN(N__12508),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__12501),
            .DIN(N__12500),
            .DOUT(N__12499),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__12501),
            .PADOUT(N__12500),
            .PADIN(N__12499),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9554),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__12492),
            .DIN(N__12491),
            .DOUT(N__12490),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__12492),
            .PADOUT(N__12491),
            .PADIN(N__12490),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10682),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__12483),
            .DIN(N__12482),
            .DOUT(N__12481),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__12483),
            .PADOUT(N__12482),
            .PADIN(N__12481),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__12474),
            .DIN(N__12473),
            .DOUT(N__12472),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__12474),
            .PADOUT(N__12473),
            .PADIN(N__12472),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__12465),
            .DIN(N__12464),
            .DOUT(N__12463),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__12465),
            .PADOUT(N__12464),
            .PADIN(N__12463),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__12456),
            .DIN(N__12455),
            .DOUT(N__12454),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__12456),
            .PADOUT(N__12455),
            .PADIN(N__12454),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__12447),
            .DIN(N__12446),
            .DOUT(N__12445),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__12447),
            .PADOUT(N__12446),
            .PADIN(N__12445),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__12438),
            .DIN(N__12437),
            .DOUT(N__12436),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__12438),
            .PADOUT(N__12437),
            .PADIN(N__12436),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__12429),
            .DIN(N__12428),
            .DOUT(N__12427),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__12429),
            .PADOUT(N__12428),
            .PADIN(N__12427),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10364),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__12420),
            .DIN(N__12419),
            .DOUT(N__12418),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__12420),
            .PADOUT(N__12419),
            .PADIN(N__12418),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8779),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__12411),
            .DIN(N__12410),
            .DOUT(N__12409),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__12411),
            .PADOUT(N__12410),
            .PADIN(N__12409),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__12402),
            .DIN(N__12401),
            .DOUT(N__12400),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__12402),
            .PADOUT(N__12401),
            .PADIN(N__12400),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5371),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__12393),
            .DIN(N__12392),
            .DOUT(N__12391),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__12393),
            .PADOUT(N__12392),
            .PADIN(N__12391),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__12384),
            .DIN(N__12383),
            .DOUT(N__12382),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__12384),
            .PADOUT(N__12383),
            .PADIN(N__12382),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__12375),
            .DIN(N__12374),
            .DOUT(N__12373),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__12375),
            .PADOUT(N__12374),
            .PADIN(N__12373),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5348),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__12366),
            .DIN(N__12365),
            .DOUT(N__12364),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__12366),
            .PADOUT(N__12365),
            .PADIN(N__12364),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__12357),
            .DIN(N__12356),
            .DOUT(N__12355),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__12357),
            .PADOUT(N__12356),
            .PADIN(N__12355),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__12348),
            .DIN(N__12347),
            .DOUT(N__12346),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__12348),
            .PADOUT(N__12347),
            .PADIN(N__12346),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9143),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__12339),
            .DIN(N__12338),
            .DOUT(N__12337),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__12339),
            .PADOUT(N__12338),
            .PADIN(N__12337),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__12330),
            .DIN(N__12329),
            .DOUT(N__12328),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__12330),
            .PADOUT(N__12329),
            .PADIN(N__12328),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9455),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__12321),
            .DIN(N__12320),
            .DOUT(N__12319),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__12321),
            .PADOUT(N__12320),
            .PADIN(N__12319),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__12312),
            .DIN(N__12311),
            .DOUT(N__12310),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__12312),
            .PADOUT(N__12311),
            .PADIN(N__12310),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7031),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__12303),
            .DIN(N__12302),
            .DOUT(N__12301),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__12303),
            .PADOUT(N__12302),
            .PADIN(N__12301),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5319),
            .DIN0(),
            .DOUT0(N__5257),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__12294),
            .DIN(N__12293),
            .DOUT(N__12292),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__12294),
            .PADOUT(N__12293),
            .PADIN(N__12292),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__12285),
            .DIN(N__12284),
            .DOUT(N__12283),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__12285),
            .PADOUT(N__12284),
            .PADIN(N__12283),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__12276),
            .DIN(N__12275),
            .DOUT(N__12274),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__12276),
            .PADOUT(N__12275),
            .PADIN(N__12274),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__12267),
            .DIN(N__12266),
            .DOUT(N__12265),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__12267),
            .PADOUT(N__12266),
            .PADIN(N__12265),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__12258),
            .DIN(N__12257),
            .DOUT(N__12256),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__12258),
            .PADOUT(N__12257),
            .PADIN(N__12256),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__12249),
            .DIN(N__12248),
            .DOUT(N__12247),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__12249),
            .PADOUT(N__12248),
            .PADIN(N__12247),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6728),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__12240),
            .DIN(N__12239),
            .DOUT(N__12238),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__12240),
            .PADOUT(N__12239),
            .PADIN(N__12238),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__12231),
            .DIN(N__12230),
            .DOUT(N__12229),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__12231),
            .PADOUT(N__12230),
            .PADIN(N__12229),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__12222),
            .DIN(N__12221),
            .DOUT(N__12220),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__12222),
            .PADOUT(N__12221),
            .PADIN(N__12220),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__12213),
            .DIN(N__12212),
            .DOUT(N__12211),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__12213),
            .PADOUT(N__12212),
            .PADIN(N__12211),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__12204),
            .DIN(N__12203),
            .DOUT(N__12202),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__12204),
            .PADOUT(N__12203),
            .PADIN(N__12202),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__12195),
            .DIN(N__12194),
            .DOUT(N__12193),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__12195),
            .PADOUT(N__12194),
            .PADIN(N__12193),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9719),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__12186),
            .DIN(N__12185),
            .DOUT(N__12184),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__12186),
            .PADOUT(N__12185),
            .PADIN(N__12184),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6503),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__12177),
            .DIN(N__12176),
            .DOUT(N__12175),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__12177),
            .PADOUT(N__12176),
            .PADIN(N__12175),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__12168),
            .DIN(N__12167),
            .DOUT(N__12166),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__12168),
            .PADOUT(N__12167),
            .PADIN(N__12166),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5441),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_0_iopad (
            .OE(N__12159),
            .DIN(N__12158),
            .DOUT(N__12157),
            .PACKAGEPIN(DA[0]));
    defparam DA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_0_preio (
            .PADOEN(N__12159),
            .PADOUT(N__12158),
            .PADIN(N__12157),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7442),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__12150),
            .DIN(N__12149),
            .DOUT(N__12148),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__12150),
            .PADOUT(N__12149),
            .PADIN(N__12148),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__12141),
            .DIN(N__12140),
            .DOUT(N__12139),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__12141),
            .PADOUT(N__12140),
            .PADIN(N__12139),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8849),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__12132),
            .DIN(N__12131),
            .DOUT(N__12130),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__12132),
            .PADOUT(N__12131),
            .PADIN(N__12130),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10487),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__12123),
            .DIN(N__12122),
            .DOUT(N__12121),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__12123),
            .PADOUT(N__12122),
            .PADIN(N__12121),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11618),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__12114),
            .DIN(N__12113),
            .DOUT(N__12112),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__12114),
            .PADOUT(N__12113),
            .PADIN(N__12112),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8627),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__12105),
            .DIN(N__12104),
            .DOUT(N__12103),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__12105),
            .PADOUT(N__12104),
            .PADIN(N__12103),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9383),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__12096),
            .DIN(N__12095),
            .DOUT(N__12094),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__12096),
            .PADOUT(N__12095),
            .PADIN(N__12094),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4412),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__12087),
            .DIN(N__12086),
            .DOUT(N__12085),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__12087),
            .PADOUT(N__12086),
            .PADIN(N__12085),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__12078),
            .DIN(N__12077),
            .DOUT(N__12076),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__12078),
            .PADOUT(N__12077),
            .PADIN(N__12076),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__12069),
            .DIN(N__12068),
            .DOUT(N__12067),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__12069),
            .PADOUT(N__12068),
            .PADIN(N__12067),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6014),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__12060),
            .DIN(N__12059),
            .DOUT(N__12058),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__12060),
            .PADOUT(N__12059),
            .PADIN(N__12058),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5323),
            .DIN0(),
            .DOUT0(N__5258),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__12051),
            .DIN(N__12050),
            .DOUT(N__12049),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__12051),
            .PADOUT(N__12050),
            .PADIN(N__12049),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9800),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__12042),
            .DIN(N__12041),
            .DOUT(N__12040),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__12042),
            .PADOUT(N__12041),
            .PADIN(N__12040),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4679),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__12033),
            .DIN(N__12032),
            .DOUT(N__12031),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__12033),
            .PADOUT(N__12032),
            .PADIN(N__12031),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8798),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__12024),
            .DIN(N__12023),
            .DOUT(N__12022),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__12024),
            .PADOUT(N__12023),
            .PADIN(N__12022),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__12015),
            .DIN(N__12014),
            .DOUT(N__12013),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__12015),
            .PADOUT(N__12014),
            .PADIN(N__12013),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_2_iopad (
            .OE(N__12006),
            .DIN(N__12005),
            .DOUT(N__12004),
            .PACKAGEPIN(DA[2]));
    defparam DA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_2_preio (
            .PADOEN(N__12006),
            .PADOUT(N__12005),
            .PADIN(N__12004),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8897),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11997),
            .DIN(N__11996),
            .DOUT(N__11995),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11997),
            .PADOUT(N__11996),
            .PADIN(N__11995),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11988),
            .DIN(N__11987),
            .DOUT(N__11986),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11988),
            .PADOUT(N__11987),
            .PADIN(N__11986),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__11979),
            .DIN(N__11978),
            .DOUT(N__11977),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__11979),
            .PADOUT(N__11978),
            .PADIN(N__11977),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8606),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__11970),
            .DIN(N__11969),
            .DOUT(N__11968),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__11970),
            .PADOUT(N__11969),
            .PADIN(N__11968),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6746),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__11961),
            .DIN(N__11960),
            .DOUT(N__11959),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__11961),
            .PADOUT(N__11960),
            .PADIN(N__11959),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__11952),
            .DIN(N__11951),
            .DOUT(N__11950),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__11952),
            .PADOUT(N__11951),
            .PADIN(N__11950),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8744),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__11943),
            .DIN(N__11942),
            .DOUT(N__11941),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__11943),
            .PADOUT(N__11942),
            .PADIN(N__11941),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5324),
            .DIN0(),
            .DOUT0(N__5253),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__11934),
            .DIN(N__11933),
            .DOUT(N__11932),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__11934),
            .PADOUT(N__11933),
            .PADIN(N__11932),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9950),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__11925),
            .DIN(N__11924),
            .DOUT(N__11923),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__11925),
            .PADOUT(N__11924),
            .PADIN(N__11923),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11916),
            .DIN(N__11915),
            .DOUT(N__11914),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11916),
            .PADOUT(N__11915),
            .PADIN(N__11914),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__11907),
            .DIN(N__11906),
            .DOUT(N__11905),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__11907),
            .PADOUT(N__11906),
            .PADIN(N__11905),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9101),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__11898),
            .DIN(N__11897),
            .DOUT(N__11896),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__11898),
            .PADOUT(N__11897),
            .PADIN(N__11896),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__11889),
            .DIN(N__11888),
            .DOUT(N__11887),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__11889),
            .PADOUT(N__11888),
            .PADIN(N__11887),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_1_iopad (
            .OE(N__11880),
            .DIN(N__11879),
            .DOUT(N__11878),
            .PACKAGEPIN(DA[1]));
    defparam DA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_1_preio (
            .PADOEN(N__11880),
            .PADOUT(N__11879),
            .PADIN(N__11878),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9002),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11871),
            .DIN(N__11870),
            .DOUT(N__11869),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11871),
            .PADOUT(N__11870),
            .PADIN(N__11869),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11862),
            .DIN(N__11861),
            .DOUT(N__11860),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11862),
            .PADOUT(N__11861),
            .PADIN(N__11860),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__11853),
            .DIN(N__11852),
            .DOUT(N__11851),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__11853),
            .PADOUT(N__11852),
            .PADIN(N__11851),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9062),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__11844),
            .DIN(N__11843),
            .DOUT(N__11842),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__11844),
            .PADOUT(N__11843),
            .PADIN(N__11842),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4757),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__11835),
            .DIN(N__11834),
            .DOUT(N__11833),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__11835),
            .PADOUT(N__11834),
            .PADIN(N__11833),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8837),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__11826),
            .DIN(N__11825),
            .DOUT(N__11824),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__11826),
            .PADOUT(N__11825),
            .PADIN(N__11824),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6419),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__11817),
            .DIN(N__11816),
            .DOUT(N__11815),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__11817),
            .PADOUT(N__11816),
            .PADIN(N__11815),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11808),
            .DIN(N__11807),
            .DOUT(N__11806),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11808),
            .PADOUT(N__11807),
            .PADIN(N__11806),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__11799),
            .DIN(N__11798),
            .DOUT(N__11797),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__11799),
            .PADOUT(N__11798),
            .PADIN(N__11797),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10508),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__11790),
            .DIN(N__11789),
            .DOUT(N__11788),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__11790),
            .PADOUT(N__11789),
            .PADIN(N__11788),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__11781),
            .DIN(N__11780),
            .DOUT(N__11779),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__11781),
            .PADOUT(N__11780),
            .PADIN(N__11779),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__11772),
            .DIN(N__11771),
            .DOUT(N__11770),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__11772),
            .PADOUT(N__11771),
            .PADIN(N__11770),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5156),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__11763),
            .DIN(N__11762),
            .DOUT(N__11761),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__11763),
            .PADOUT(N__11762),
            .PADIN(N__11761),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4709),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11754),
            .DIN(N__11753),
            .DOUT(N__11752),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11754),
            .PADOUT(N__11753),
            .PADIN(N__11752),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5102),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11745),
            .DIN(N__11744),
            .DOUT(N__11743),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11745),
            .PADOUT(N__11744),
            .PADIN(N__11743),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11736),
            .DIN(N__11735),
            .DOUT(N__11734),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11736),
            .PADOUT(N__11735),
            .PADIN(N__11734),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5101),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11727),
            .DIN(N__11726),
            .DOUT(N__11725),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11727),
            .PADOUT(N__11726),
            .PADIN(N__11725),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4280),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11718),
            .DIN(N__11717),
            .DOUT(N__11716),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11718),
            .PADOUT(N__11717),
            .PADIN(N__11716),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9926),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11709),
            .DIN(N__11708),
            .DOUT(N__11707),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11709),
            .PADOUT(N__11708),
            .PADIN(N__11707),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11700),
            .DIN(N__11699),
            .DOUT(N__11698),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11700),
            .PADOUT(N__11699),
            .PADIN(N__11698),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11691),
            .DIN(N__11690),
            .DOUT(N__11689),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11691),
            .PADOUT(N__11690),
            .PADIN(N__11689),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11682),
            .DIN(N__11681),
            .DOUT(N__11680),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11682),
            .PADOUT(N__11681),
            .PADIN(N__11680),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11673),
            .DIN(N__11672),
            .DOUT(N__11671),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11673),
            .PADOUT(N__11672),
            .PADIN(N__11671),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5088),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2838 (
            .O(N__11654),
            .I(N__11650));
    InMux I__2837 (
            .O(N__11653),
            .I(N__11647));
    LocalMux I__2836 (
            .O(N__11650),
            .I(N__11644));
    LocalMux I__2835 (
            .O(N__11647),
            .I(N__11641));
    Span12Mux_s9_h I__2834 (
            .O(N__11644),
            .I(N__11638));
    Span4Mux_h I__2833 (
            .O(N__11641),
            .I(N__11635));
    Span12Mux_h I__2832 (
            .O(N__11638),
            .I(N__11631));
    Span4Mux_v I__2831 (
            .O(N__11635),
            .I(N__11628));
    InMux I__2830 (
            .O(N__11634),
            .I(N__11625));
    Odrv12 I__2829 (
            .O(N__11631),
            .I(REG_CYCLEm));
    Odrv4 I__2828 (
            .O(N__11628),
            .I(REG_CYCLEm));
    LocalMux I__2827 (
            .O(N__11625),
            .I(REG_CYCLEm));
    IoInMux I__2826 (
            .O(N__11618),
            .I(N__11615));
    LocalMux I__2825 (
            .O(N__11615),
            .I(N__11612));
    Span4Mux_s2_v I__2824 (
            .O(N__11612),
            .I(N__11609));
    Span4Mux_v I__2823 (
            .O(N__11609),
            .I(N__11606));
    Odrv4 I__2822 (
            .O(N__11606),
            .I(DRDENn_c));
    InMux I__2821 (
            .O(N__11603),
            .I(N__11600));
    LocalMux I__2820 (
            .O(N__11600),
            .I(N__11597));
    Odrv12 I__2819 (
            .O(N__11597),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2818 (
            .O(N__11594),
            .I(N__11590));
    InMux I__2817 (
            .O(N__11593),
            .I(N__11586));
    LocalMux I__2816 (
            .O(N__11590),
            .I(N__11583));
    InMux I__2815 (
            .O(N__11589),
            .I(N__11580));
    LocalMux I__2814 (
            .O(N__11586),
            .I(N__11572));
    Span4Mux_v I__2813 (
            .O(N__11583),
            .I(N__11572));
    LocalMux I__2812 (
            .O(N__11580),
            .I(N__11572));
    InMux I__2811 (
            .O(N__11579),
            .I(N__11569));
    Span4Mux_h I__2810 (
            .O(N__11572),
            .I(N__11566));
    LocalMux I__2809 (
            .O(N__11569),
            .I(N__11563));
    Span4Mux_v I__2808 (
            .O(N__11566),
            .I(N__11560));
    Sp12to4 I__2807 (
            .O(N__11563),
            .I(N__11557));
    Sp12to4 I__2806 (
            .O(N__11560),
            .I(N__11552));
    Span12Mux_v I__2805 (
            .O(N__11557),
            .I(N__11552));
    Odrv12 I__2804 (
            .O(N__11552),
            .I(DRA_c_2));
    InMux I__2803 (
            .O(N__11549),
            .I(N__11543));
    InMux I__2802 (
            .O(N__11548),
            .I(N__11543));
    LocalMux I__2801 (
            .O(N__11543),
            .I(N__11540));
    Span4Mux_h I__2800 (
            .O(N__11540),
            .I(N__11537));
    Odrv4 I__2799 (
            .O(N__11537),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2798 (
            .O(N__11534),
            .I(N__11531));
    LocalMux I__2797 (
            .O(N__11531),
            .I(N__11527));
    InMux I__2796 (
            .O(N__11530),
            .I(N__11524));
    Span4Mux_h I__2795 (
            .O(N__11527),
            .I(N__11517));
    LocalMux I__2794 (
            .O(N__11524),
            .I(N__11517));
    InMux I__2793 (
            .O(N__11523),
            .I(N__11514));
    InMux I__2792 (
            .O(N__11522),
            .I(N__11511));
    Span4Mux_h I__2791 (
            .O(N__11517),
            .I(N__11504));
    LocalMux I__2790 (
            .O(N__11514),
            .I(N__11504));
    LocalMux I__2789 (
            .O(N__11511),
            .I(N__11504));
    Span4Mux_v I__2788 (
            .O(N__11504),
            .I(N__11501));
    Span4Mux_v I__2787 (
            .O(N__11501),
            .I(N__11498));
    Sp12to4 I__2786 (
            .O(N__11498),
            .I(N__11495));
    Odrv12 I__2785 (
            .O(N__11495),
            .I(DRA_c_1));
    InMux I__2784 (
            .O(N__11492),
            .I(N__11488));
    InMux I__2783 (
            .O(N__11491),
            .I(N__11485));
    LocalMux I__2782 (
            .O(N__11488),
            .I(N__11480));
    LocalMux I__2781 (
            .O(N__11485),
            .I(N__11480));
    Span4Mux_h I__2780 (
            .O(N__11480),
            .I(N__11477));
    Sp12to4 I__2779 (
            .O(N__11477),
            .I(N__11474));
    Span12Mux_v I__2778 (
            .O(N__11474),
            .I(N__11471));
    Odrv12 I__2777 (
            .O(N__11471),
            .I(DRA_c_0));
    InMux I__2776 (
            .O(N__11468),
            .I(N__11465));
    LocalMux I__2775 (
            .O(N__11465),
            .I(N__11462));
    Span4Mux_h I__2774 (
            .O(N__11462),
            .I(N__11459));
    Odrv4 I__2773 (
            .O(N__11459),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2772 (
            .O(N__11456),
            .I(N__11452));
    InMux I__2771 (
            .O(N__11455),
            .I(N__11448));
    LocalMux I__2770 (
            .O(N__11452),
            .I(N__11444));
    InMux I__2769 (
            .O(N__11451),
            .I(N__11441));
    LocalMux I__2768 (
            .O(N__11448),
            .I(N__11438));
    InMux I__2767 (
            .O(N__11447),
            .I(N__11435));
    Span12Mux_v I__2766 (
            .O(N__11444),
            .I(N__11430));
    LocalMux I__2765 (
            .O(N__11441),
            .I(N__11430));
    Span4Mux_v I__2764 (
            .O(N__11438),
            .I(N__11427));
    LocalMux I__2763 (
            .O(N__11435),
            .I(N__11424));
    Span12Mux_h I__2762 (
            .O(N__11430),
            .I(N__11421));
    Sp12to4 I__2761 (
            .O(N__11427),
            .I(N__11416));
    Span12Mux_v I__2760 (
            .O(N__11424),
            .I(N__11416));
    Odrv12 I__2759 (
            .O(N__11421),
            .I(DRA_c_8));
    Odrv12 I__2758 (
            .O(N__11416),
            .I(DRA_c_8));
    InMux I__2757 (
            .O(N__11411),
            .I(N__11408));
    LocalMux I__2756 (
            .O(N__11408),
            .I(N__11405));
    Odrv4 I__2755 (
            .O(N__11405),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2754 (
            .O(N__11402),
            .I(N__11399));
    LocalMux I__2753 (
            .O(N__11399),
            .I(N__11396));
    Span4Mux_v I__2752 (
            .O(N__11396),
            .I(N__11390));
    InMux I__2751 (
            .O(N__11395),
            .I(N__11387));
    InMux I__2750 (
            .O(N__11394),
            .I(N__11382));
    InMux I__2749 (
            .O(N__11393),
            .I(N__11382));
    Span4Mux_h I__2748 (
            .O(N__11390),
            .I(N__11379));
    LocalMux I__2747 (
            .O(N__11387),
            .I(N__11374));
    LocalMux I__2746 (
            .O(N__11382),
            .I(N__11374));
    Sp12to4 I__2745 (
            .O(N__11379),
            .I(N__11369));
    Span12Mux_h I__2744 (
            .O(N__11374),
            .I(N__11369));
    Odrv12 I__2743 (
            .O(N__11369),
            .I(DRA_c_7));
    InMux I__2742 (
            .O(N__11366),
            .I(N__11362));
    InMux I__2741 (
            .O(N__11365),
            .I(N__11359));
    LocalMux I__2740 (
            .O(N__11362),
            .I(N__11353));
    LocalMux I__2739 (
            .O(N__11359),
            .I(N__11353));
    InMux I__2738 (
            .O(N__11358),
            .I(N__11349));
    Span4Mux_v I__2737 (
            .O(N__11353),
            .I(N__11346));
    InMux I__2736 (
            .O(N__11352),
            .I(N__11343));
    LocalMux I__2735 (
            .O(N__11349),
            .I(N__11340));
    Sp12to4 I__2734 (
            .O(N__11346),
            .I(N__11337));
    LocalMux I__2733 (
            .O(N__11343),
            .I(N__11334));
    Span4Mux_v I__2732 (
            .O(N__11340),
            .I(N__11331));
    Span12Mux_h I__2731 (
            .O(N__11337),
            .I(N__11328));
    Span12Mux_v I__2730 (
            .O(N__11334),
            .I(N__11323));
    Sp12to4 I__2729 (
            .O(N__11331),
            .I(N__11323));
    Odrv12 I__2728 (
            .O(N__11328),
            .I(DRA_c_6));
    Odrv12 I__2727 (
            .O(N__11323),
            .I(DRA_c_6));
    InMux I__2726 (
            .O(N__11318),
            .I(N__11315));
    LocalMux I__2725 (
            .O(N__11315),
            .I(N__11312));
    Odrv4 I__2724 (
            .O(N__11312),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2723 (
            .O(N__11309),
            .I(N__11306));
    LocalMux I__2722 (
            .O(N__11306),
            .I(N__11303));
    Span12Mux_v I__2721 (
            .O(N__11303),
            .I(N__11300));
    Odrv12 I__2720 (
            .O(N__11300),
            .I(RAS0n_c));
    InMux I__2719 (
            .O(N__11297),
            .I(N__11294));
    LocalMux I__2718 (
            .O(N__11294),
            .I(N__11276));
    InMux I__2717 (
            .O(N__11293),
            .I(N__11269));
    InMux I__2716 (
            .O(N__11292),
            .I(N__11269));
    InMux I__2715 (
            .O(N__11291),
            .I(N__11262));
    InMux I__2714 (
            .O(N__11290),
            .I(N__11262));
    InMux I__2713 (
            .O(N__11289),
            .I(N__11262));
    InMux I__2712 (
            .O(N__11288),
            .I(N__11259));
    InMux I__2711 (
            .O(N__11287),
            .I(N__11256));
    InMux I__2710 (
            .O(N__11286),
            .I(N__11253));
    InMux I__2709 (
            .O(N__11285),
            .I(N__11250));
    InMux I__2708 (
            .O(N__11284),
            .I(N__11247));
    InMux I__2707 (
            .O(N__11283),
            .I(N__11244));
    InMux I__2706 (
            .O(N__11282),
            .I(N__11241));
    InMux I__2705 (
            .O(N__11281),
            .I(N__11238));
    InMux I__2704 (
            .O(N__11280),
            .I(N__11235));
    InMux I__2703 (
            .O(N__11279),
            .I(N__11230));
    Span4Mux_v I__2702 (
            .O(N__11276),
            .I(N__11226));
    InMux I__2701 (
            .O(N__11275),
            .I(N__11223));
    InMux I__2700 (
            .O(N__11274),
            .I(N__11220));
    LocalMux I__2699 (
            .O(N__11269),
            .I(N__11217));
    LocalMux I__2698 (
            .O(N__11262),
            .I(N__11210));
    LocalMux I__2697 (
            .O(N__11259),
            .I(N__11210));
    LocalMux I__2696 (
            .O(N__11256),
            .I(N__11210));
    LocalMux I__2695 (
            .O(N__11253),
            .I(N__11207));
    LocalMux I__2694 (
            .O(N__11250),
            .I(N__11194));
    LocalMux I__2693 (
            .O(N__11247),
            .I(N__11194));
    LocalMux I__2692 (
            .O(N__11244),
            .I(N__11194));
    LocalMux I__2691 (
            .O(N__11241),
            .I(N__11194));
    LocalMux I__2690 (
            .O(N__11238),
            .I(N__11194));
    LocalMux I__2689 (
            .O(N__11235),
            .I(N__11194));
    InMux I__2688 (
            .O(N__11234),
            .I(N__11191));
    InMux I__2687 (
            .O(N__11233),
            .I(N__11188));
    LocalMux I__2686 (
            .O(N__11230),
            .I(N__11185));
    InMux I__2685 (
            .O(N__11229),
            .I(N__11182));
    Span4Mux_h I__2684 (
            .O(N__11226),
            .I(N__11171));
    LocalMux I__2683 (
            .O(N__11223),
            .I(N__11171));
    LocalMux I__2682 (
            .O(N__11220),
            .I(N__11171));
    Span4Mux_v I__2681 (
            .O(N__11217),
            .I(N__11171));
    Span4Mux_v I__2680 (
            .O(N__11210),
            .I(N__11171));
    Span4Mux_v I__2679 (
            .O(N__11207),
            .I(N__11166));
    Span4Mux_v I__2678 (
            .O(N__11194),
            .I(N__11166));
    LocalMux I__2677 (
            .O(N__11191),
            .I(N__11161));
    LocalMux I__2676 (
            .O(N__11188),
            .I(N__11161));
    Span4Mux_h I__2675 (
            .O(N__11185),
            .I(N__11158));
    LocalMux I__2674 (
            .O(N__11182),
            .I(N__11151));
    Sp12to4 I__2673 (
            .O(N__11171),
            .I(N__11151));
    Sp12to4 I__2672 (
            .O(N__11166),
            .I(N__11151));
    Span12Mux_v I__2671 (
            .O(N__11161),
            .I(N__11148));
    Sp12to4 I__2670 (
            .O(N__11158),
            .I(N__11143));
    Span12Mux_h I__2669 (
            .O(N__11151),
            .I(N__11143));
    Span12Mux_h I__2668 (
            .O(N__11148),
            .I(N__11140));
    Span12Mux_v I__2667 (
            .O(N__11143),
            .I(N__11137));
    Odrv12 I__2666 (
            .O(N__11140),
            .I(AGNUS_REV_c));
    Odrv12 I__2665 (
            .O(N__11137),
            .I(AGNUS_REV_c));
    InMux I__2664 (
            .O(N__11132),
            .I(N__11128));
    InMux I__2663 (
            .O(N__11131),
            .I(N__11125));
    LocalMux I__2662 (
            .O(N__11128),
            .I(N__11118));
    LocalMux I__2661 (
            .O(N__11125),
            .I(N__11118));
    InMux I__2660 (
            .O(N__11124),
            .I(N__11115));
    InMux I__2659 (
            .O(N__11123),
            .I(N__11112));
    Span12Mux_v I__2658 (
            .O(N__11118),
            .I(N__11109));
    LocalMux I__2657 (
            .O(N__11115),
            .I(N__11106));
    LocalMux I__2656 (
            .O(N__11112),
            .I(N__11103));
    Span12Mux_h I__2655 (
            .O(N__11109),
            .I(N__11100));
    Span12Mux_v I__2654 (
            .O(N__11106),
            .I(N__11097));
    Span12Mux_v I__2653 (
            .O(N__11103),
            .I(N__11094));
    Span12Mux_v I__2652 (
            .O(N__11100),
            .I(N__11089));
    Span12Mux_h I__2651 (
            .O(N__11097),
            .I(N__11089));
    Span12Mux_v I__2650 (
            .O(N__11094),
            .I(N__11086));
    Odrv12 I__2649 (
            .O(N__11089),
            .I(DRA_c_9));
    Odrv12 I__2648 (
            .O(N__11086),
            .I(DRA_c_9));
    InMux I__2647 (
            .O(N__11081),
            .I(N__11078));
    LocalMux I__2646 (
            .O(N__11078),
            .I(N__11075));
    Span12Mux_v I__2645 (
            .O(N__11075),
            .I(N__11072));
    Odrv12 I__2644 (
            .O(N__11072),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    ClkMux I__2643 (
            .O(N__11069),
            .I(N__11042));
    ClkMux I__2642 (
            .O(N__11068),
            .I(N__11042));
    ClkMux I__2641 (
            .O(N__11067),
            .I(N__11042));
    ClkMux I__2640 (
            .O(N__11066),
            .I(N__11042));
    ClkMux I__2639 (
            .O(N__11065),
            .I(N__11042));
    ClkMux I__2638 (
            .O(N__11064),
            .I(N__11042));
    ClkMux I__2637 (
            .O(N__11063),
            .I(N__11042));
    ClkMux I__2636 (
            .O(N__11062),
            .I(N__11042));
    ClkMux I__2635 (
            .O(N__11061),
            .I(N__11042));
    GlobalMux I__2634 (
            .O(N__11042),
            .I(N__11039));
    gio2CtrlBuf I__2633 (
            .O(N__11039),
            .I(C3_c_g));
    CEMux I__2632 (
            .O(N__11036),
            .I(N__10988));
    CEMux I__2631 (
            .O(N__11035),
            .I(N__10988));
    CEMux I__2630 (
            .O(N__11034),
            .I(N__10988));
    CEMux I__2629 (
            .O(N__11033),
            .I(N__10988));
    CEMux I__2628 (
            .O(N__11032),
            .I(N__10988));
    CEMux I__2627 (
            .O(N__11031),
            .I(N__10988));
    CEMux I__2626 (
            .O(N__11030),
            .I(N__10988));
    CEMux I__2625 (
            .O(N__11029),
            .I(N__10988));
    CEMux I__2624 (
            .O(N__11028),
            .I(N__10988));
    CEMux I__2623 (
            .O(N__11027),
            .I(N__10988));
    CEMux I__2622 (
            .O(N__11026),
            .I(N__10988));
    CEMux I__2621 (
            .O(N__11025),
            .I(N__10988));
    CEMux I__2620 (
            .O(N__11024),
            .I(N__10988));
    CEMux I__2619 (
            .O(N__11023),
            .I(N__10988));
    CEMux I__2618 (
            .O(N__11022),
            .I(N__10988));
    CEMux I__2617 (
            .O(N__11021),
            .I(N__10988));
    GlobalMux I__2616 (
            .O(N__10988),
            .I(N__10985));
    gio2CtrlBuf I__2615 (
            .O(N__10985),
            .I(DBRn_c_i_0_g));
    InMux I__2614 (
            .O(N__10982),
            .I(N__10976));
    InMux I__2613 (
            .O(N__10981),
            .I(N__10973));
    InMux I__2612 (
            .O(N__10980),
            .I(N__10970));
    InMux I__2611 (
            .O(N__10979),
            .I(N__10967));
    LocalMux I__2610 (
            .O(N__10976),
            .I(N__10959));
    LocalMux I__2609 (
            .O(N__10973),
            .I(N__10935));
    LocalMux I__2608 (
            .O(N__10970),
            .I(N__10919));
    LocalMux I__2607 (
            .O(N__10967),
            .I(N__10914));
    SRMux I__2606 (
            .O(N__10966),
            .I(N__10820));
    SRMux I__2605 (
            .O(N__10965),
            .I(N__10820));
    SRMux I__2604 (
            .O(N__10964),
            .I(N__10820));
    SRMux I__2603 (
            .O(N__10963),
            .I(N__10820));
    SRMux I__2602 (
            .O(N__10962),
            .I(N__10820));
    Glb2LocalMux I__2601 (
            .O(N__10959),
            .I(N__10820));
    SRMux I__2600 (
            .O(N__10958),
            .I(N__10820));
    SRMux I__2599 (
            .O(N__10957),
            .I(N__10820));
    SRMux I__2598 (
            .O(N__10956),
            .I(N__10820));
    SRMux I__2597 (
            .O(N__10955),
            .I(N__10820));
    SRMux I__2596 (
            .O(N__10954),
            .I(N__10820));
    SRMux I__2595 (
            .O(N__10953),
            .I(N__10820));
    SRMux I__2594 (
            .O(N__10952),
            .I(N__10820));
    SRMux I__2593 (
            .O(N__10951),
            .I(N__10820));
    SRMux I__2592 (
            .O(N__10950),
            .I(N__10820));
    SRMux I__2591 (
            .O(N__10949),
            .I(N__10820));
    SRMux I__2590 (
            .O(N__10948),
            .I(N__10820));
    SRMux I__2589 (
            .O(N__10947),
            .I(N__10820));
    SRMux I__2588 (
            .O(N__10946),
            .I(N__10820));
    SRMux I__2587 (
            .O(N__10945),
            .I(N__10820));
    SRMux I__2586 (
            .O(N__10944),
            .I(N__10820));
    SRMux I__2585 (
            .O(N__10943),
            .I(N__10820));
    SRMux I__2584 (
            .O(N__10942),
            .I(N__10820));
    SRMux I__2583 (
            .O(N__10941),
            .I(N__10820));
    SRMux I__2582 (
            .O(N__10940),
            .I(N__10820));
    SRMux I__2581 (
            .O(N__10939),
            .I(N__10820));
    SRMux I__2580 (
            .O(N__10938),
            .I(N__10820));
    Glb2LocalMux I__2579 (
            .O(N__10935),
            .I(N__10820));
    SRMux I__2578 (
            .O(N__10934),
            .I(N__10820));
    SRMux I__2577 (
            .O(N__10933),
            .I(N__10820));
    SRMux I__2576 (
            .O(N__10932),
            .I(N__10820));
    SRMux I__2575 (
            .O(N__10931),
            .I(N__10820));
    SRMux I__2574 (
            .O(N__10930),
            .I(N__10820));
    SRMux I__2573 (
            .O(N__10929),
            .I(N__10820));
    SRMux I__2572 (
            .O(N__10928),
            .I(N__10820));
    SRMux I__2571 (
            .O(N__10927),
            .I(N__10820));
    SRMux I__2570 (
            .O(N__10926),
            .I(N__10820));
    SRMux I__2569 (
            .O(N__10925),
            .I(N__10820));
    SRMux I__2568 (
            .O(N__10924),
            .I(N__10820));
    SRMux I__2567 (
            .O(N__10923),
            .I(N__10820));
    SRMux I__2566 (
            .O(N__10922),
            .I(N__10820));
    Glb2LocalMux I__2565 (
            .O(N__10919),
            .I(N__10820));
    SRMux I__2564 (
            .O(N__10918),
            .I(N__10820));
    SRMux I__2563 (
            .O(N__10917),
            .I(N__10820));
    Glb2LocalMux I__2562 (
            .O(N__10914),
            .I(N__10820));
    SRMux I__2561 (
            .O(N__10913),
            .I(N__10820));
    GlobalMux I__2560 (
            .O(N__10820),
            .I(N__10817));
    gio2CtrlBuf I__2559 (
            .O(N__10817),
            .I(RESETn_c_i_g));
    InMux I__2558 (
            .O(N__10814),
            .I(N__10810));
    InMux I__2557 (
            .O(N__10813),
            .I(N__10807));
    LocalMux I__2556 (
            .O(N__10810),
            .I(N__10802));
    LocalMux I__2555 (
            .O(N__10807),
            .I(N__10798));
    InMux I__2554 (
            .O(N__10806),
            .I(N__10795));
    InMux I__2553 (
            .O(N__10805),
            .I(N__10792));
    Span4Mux_v I__2552 (
            .O(N__10802),
            .I(N__10789));
    InMux I__2551 (
            .O(N__10801),
            .I(N__10786));
    Span4Mux_v I__2550 (
            .O(N__10798),
            .I(N__10781));
    LocalMux I__2549 (
            .O(N__10795),
            .I(N__10781));
    LocalMux I__2548 (
            .O(N__10792),
            .I(N__10778));
    Sp12to4 I__2547 (
            .O(N__10789),
            .I(N__10775));
    LocalMux I__2546 (
            .O(N__10786),
            .I(N__10772));
    Span4Mux_v I__2545 (
            .O(N__10781),
            .I(N__10769));
    Span4Mux_v I__2544 (
            .O(N__10778),
            .I(N__10766));
    Span12Mux_h I__2543 (
            .O(N__10775),
            .I(N__10761));
    Span12Mux_v I__2542 (
            .O(N__10772),
            .I(N__10761));
    Sp12to4 I__2541 (
            .O(N__10769),
            .I(N__10756));
    Sp12to4 I__2540 (
            .O(N__10766),
            .I(N__10756));
    Span12Mux_h I__2539 (
            .O(N__10761),
            .I(N__10753));
    Span12Mux_h I__2538 (
            .O(N__10756),
            .I(N__10750));
    Odrv12 I__2537 (
            .O(N__10753),
            .I(RnW_c));
    Odrv12 I__2536 (
            .O(N__10750),
            .I(RnW_c));
    CascadeMux I__2535 (
            .O(N__10745),
            .I(N__10742));
    InMux I__2534 (
            .O(N__10742),
            .I(N__10739));
    LocalMux I__2533 (
            .O(N__10739),
            .I(N__10735));
    InMux I__2532 (
            .O(N__10738),
            .I(N__10732));
    Span12Mux_s10_v I__2531 (
            .O(N__10735),
            .I(N__10729));
    LocalMux I__2530 (
            .O(N__10732),
            .I(N__10726));
    Span12Mux_h I__2529 (
            .O(N__10729),
            .I(N__10717));
    Span12Mux_v I__2528 (
            .O(N__10726),
            .I(N__10714));
    InMux I__2527 (
            .O(N__10725),
            .I(N__10711));
    InMux I__2526 (
            .O(N__10724),
            .I(N__10708));
    InMux I__2525 (
            .O(N__10723),
            .I(N__10705));
    InMux I__2524 (
            .O(N__10722),
            .I(N__10700));
    InMux I__2523 (
            .O(N__10721),
            .I(N__10700));
    InMux I__2522 (
            .O(N__10720),
            .I(N__10697));
    Odrv12 I__2521 (
            .O(N__10717),
            .I(WRITE_CYCLEm));
    Odrv12 I__2520 (
            .O(N__10714),
            .I(WRITE_CYCLEm));
    LocalMux I__2519 (
            .O(N__10711),
            .I(WRITE_CYCLEm));
    LocalMux I__2518 (
            .O(N__10708),
            .I(WRITE_CYCLEm));
    LocalMux I__2517 (
            .O(N__10705),
            .I(WRITE_CYCLEm));
    LocalMux I__2516 (
            .O(N__10700),
            .I(WRITE_CYCLEm));
    LocalMux I__2515 (
            .O(N__10697),
            .I(WRITE_CYCLEm));
    IoInMux I__2514 (
            .O(N__10682),
            .I(N__10679));
    LocalMux I__2513 (
            .O(N__10679),
            .I(N__10676));
    Span4Mux_s3_h I__2512 (
            .O(N__10676),
            .I(N__10673));
    Span4Mux_v I__2511 (
            .O(N__10673),
            .I(N__10670));
    Odrv4 I__2510 (
            .O(N__10670),
            .I(DRDDIR_c));
    InMux I__2509 (
            .O(N__10667),
            .I(N__10662));
    InMux I__2508 (
            .O(N__10666),
            .I(N__10656));
    InMux I__2507 (
            .O(N__10665),
            .I(N__10656));
    LocalMux I__2506 (
            .O(N__10662),
            .I(N__10653));
    InMux I__2505 (
            .O(N__10661),
            .I(N__10650));
    LocalMux I__2504 (
            .O(N__10656),
            .I(N__10647));
    Span4Mux_v I__2503 (
            .O(N__10653),
            .I(N__10644));
    LocalMux I__2502 (
            .O(N__10650),
            .I(N__10641));
    Span4Mux_v I__2501 (
            .O(N__10647),
            .I(N__10638));
    Sp12to4 I__2500 (
            .O(N__10644),
            .I(N__10633));
    Sp12to4 I__2499 (
            .O(N__10641),
            .I(N__10630));
    Sp12to4 I__2498 (
            .O(N__10638),
            .I(N__10627));
    InMux I__2497 (
            .O(N__10637),
            .I(N__10622));
    InMux I__2496 (
            .O(N__10636),
            .I(N__10622));
    Span12Mux_h I__2495 (
            .O(N__10633),
            .I(N__10619));
    Span12Mux_v I__2494 (
            .O(N__10630),
            .I(N__10616));
    Span12Mux_h I__2493 (
            .O(N__10627),
            .I(N__10611));
    LocalMux I__2492 (
            .O(N__10622),
            .I(N__10611));
    Span12Mux_v I__2491 (
            .O(N__10619),
            .I(N__10608));
    Span12Mux_h I__2490 (
            .O(N__10616),
            .I(N__10603));
    Span12Mux_v I__2489 (
            .O(N__10611),
            .I(N__10603));
    Odrv12 I__2488 (
            .O(N__10608),
            .I(CASLn_c));
    Odrv12 I__2487 (
            .O(N__10603),
            .I(CASLn_c));
    CascadeMux I__2486 (
            .O(N__10598),
            .I(N__10595));
    InMux I__2485 (
            .O(N__10595),
            .I(N__10592));
    LocalMux I__2484 (
            .O(N__10592),
            .I(N__10589));
    Span4Mux_v I__2483 (
            .O(N__10589),
            .I(N__10585));
    InMux I__2482 (
            .O(N__10588),
            .I(N__10581));
    Span4Mux_v I__2481 (
            .O(N__10585),
            .I(N__10577));
    InMux I__2480 (
            .O(N__10584),
            .I(N__10574));
    LocalMux I__2479 (
            .O(N__10581),
            .I(N__10570));
    InMux I__2478 (
            .O(N__10580),
            .I(N__10567));
    Span4Mux_v I__2477 (
            .O(N__10577),
            .I(N__10562));
    LocalMux I__2476 (
            .O(N__10574),
            .I(N__10562));
    CascadeMux I__2475 (
            .O(N__10573),
            .I(N__10559));
    Sp12to4 I__2474 (
            .O(N__10570),
            .I(N__10555));
    LocalMux I__2473 (
            .O(N__10567),
            .I(N__10552));
    Span4Mux_v I__2472 (
            .O(N__10562),
            .I(N__10549));
    InMux I__2471 (
            .O(N__10559),
            .I(N__10544));
    InMux I__2470 (
            .O(N__10558),
            .I(N__10544));
    Span12Mux_v I__2469 (
            .O(N__10555),
            .I(N__10541));
    Span12Mux_h I__2468 (
            .O(N__10552),
            .I(N__10538));
    Sp12to4 I__2467 (
            .O(N__10549),
            .I(N__10535));
    LocalMux I__2466 (
            .O(N__10544),
            .I(N__10532));
    Span12Mux_h I__2465 (
            .O(N__10541),
            .I(N__10529));
    Span12Mux_v I__2464 (
            .O(N__10538),
            .I(N__10524));
    Span12Mux_h I__2463 (
            .O(N__10535),
            .I(N__10524));
    Span4Mux_v I__2462 (
            .O(N__10532),
            .I(N__10521));
    Odrv12 I__2461 (
            .O(N__10529),
            .I(CASUn_c));
    Odrv12 I__2460 (
            .O(N__10524),
            .I(CASUn_c));
    Odrv4 I__2459 (
            .O(N__10521),
            .I(CASUn_c));
    InMux I__2458 (
            .O(N__10514),
            .I(N__10511));
    LocalMux I__2457 (
            .O(N__10511),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__2456 (
            .O(N__10508),
            .I(N__10505));
    LocalMux I__2455 (
            .O(N__10505),
            .I(N__10502));
    Span12Mux_s4_h I__2454 (
            .O(N__10502),
            .I(N__10499));
    Span12Mux_v I__2453 (
            .O(N__10499),
            .I(N__10496));
    Odrv12 I__2452 (
            .O(N__10496),
            .I(CMA_c_6));
    InMux I__2451 (
            .O(N__10493),
            .I(N__10490));
    LocalMux I__2450 (
            .O(N__10490),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__2449 (
            .O(N__10487),
            .I(N__10484));
    LocalMux I__2448 (
            .O(N__10484),
            .I(N__10481));
    IoSpan4Mux I__2447 (
            .O(N__10481),
            .I(N__10478));
    Span4Mux_s0_h I__2446 (
            .O(N__10478),
            .I(N__10475));
    Sp12to4 I__2445 (
            .O(N__10475),
            .I(N__10472));
    Span12Mux_v I__2444 (
            .O(N__10472),
            .I(N__10469));
    Odrv12 I__2443 (
            .O(N__10469),
            .I(CMA_c_4));
    InMux I__2442 (
            .O(N__10466),
            .I(N__10457));
    InMux I__2441 (
            .O(N__10465),
            .I(N__10457));
    InMux I__2440 (
            .O(N__10464),
            .I(N__10457));
    LocalMux I__2439 (
            .O(N__10457),
            .I(N__10451));
    InMux I__2438 (
            .O(N__10456),
            .I(N__10444));
    InMux I__2437 (
            .O(N__10455),
            .I(N__10444));
    InMux I__2436 (
            .O(N__10454),
            .I(N__10444));
    Odrv4 I__2435 (
            .O(N__10451),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ));
    LocalMux I__2434 (
            .O(N__10444),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ));
    CascadeMux I__2433 (
            .O(N__10439),
            .I(N__10432));
    CascadeMux I__2432 (
            .O(N__10438),
            .I(N__10429));
    CascadeMux I__2431 (
            .O(N__10437),
            .I(N__10426));
    CascadeMux I__2430 (
            .O(N__10436),
            .I(N__10422));
    CascadeMux I__2429 (
            .O(N__10435),
            .I(N__10419));
    InMux I__2428 (
            .O(N__10432),
            .I(N__10412));
    InMux I__2427 (
            .O(N__10429),
            .I(N__10412));
    InMux I__2426 (
            .O(N__10426),
            .I(N__10412));
    InMux I__2425 (
            .O(N__10425),
            .I(N__10408));
    InMux I__2424 (
            .O(N__10422),
            .I(N__10403));
    InMux I__2423 (
            .O(N__10419),
            .I(N__10403));
    LocalMux I__2422 (
            .O(N__10412),
            .I(N__10400));
    CascadeMux I__2421 (
            .O(N__10411),
            .I(N__10395));
    LocalMux I__2420 (
            .O(N__10408),
            .I(N__10390));
    LocalMux I__2419 (
            .O(N__10403),
            .I(N__10390));
    Span4Mux_h I__2418 (
            .O(N__10400),
            .I(N__10387));
    InMux I__2417 (
            .O(N__10399),
            .I(N__10384));
    InMux I__2416 (
            .O(N__10398),
            .I(N__10379));
    InMux I__2415 (
            .O(N__10395),
            .I(N__10379));
    Odrv12 I__2414 (
            .O(N__10390),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__2413 (
            .O(N__10387),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__2412 (
            .O(N__10384),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__2411 (
            .O(N__10379),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    InMux I__2410 (
            .O(N__10370),
            .I(N__10367));
    LocalMux I__2409 (
            .O(N__10367),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__2408 (
            .O(N__10364),
            .I(N__10361));
    LocalMux I__2407 (
            .O(N__10361),
            .I(N__10358));
    IoSpan4Mux I__2406 (
            .O(N__10358),
            .I(N__10355));
    Span4Mux_s2_h I__2405 (
            .O(N__10355),
            .I(N__10352));
    Sp12to4 I__2404 (
            .O(N__10352),
            .I(N__10349));
    Span12Mux_v I__2403 (
            .O(N__10349),
            .I(N__10346));
    Odrv12 I__2402 (
            .O(N__10346),
            .I(CMA_c_7));
    InMux I__2401 (
            .O(N__10343),
            .I(N__10340));
    LocalMux I__2400 (
            .O(N__10340),
            .I(N__10301));
    ClkMux I__2399 (
            .O(N__10339),
            .I(N__10202));
    ClkMux I__2398 (
            .O(N__10338),
            .I(N__10202));
    ClkMux I__2397 (
            .O(N__10337),
            .I(N__10202));
    ClkMux I__2396 (
            .O(N__10336),
            .I(N__10202));
    ClkMux I__2395 (
            .O(N__10335),
            .I(N__10202));
    ClkMux I__2394 (
            .O(N__10334),
            .I(N__10202));
    ClkMux I__2393 (
            .O(N__10333),
            .I(N__10202));
    ClkMux I__2392 (
            .O(N__10332),
            .I(N__10202));
    ClkMux I__2391 (
            .O(N__10331),
            .I(N__10202));
    ClkMux I__2390 (
            .O(N__10330),
            .I(N__10202));
    ClkMux I__2389 (
            .O(N__10329),
            .I(N__10202));
    ClkMux I__2388 (
            .O(N__10328),
            .I(N__10202));
    ClkMux I__2387 (
            .O(N__10327),
            .I(N__10202));
    ClkMux I__2386 (
            .O(N__10326),
            .I(N__10202));
    ClkMux I__2385 (
            .O(N__10325),
            .I(N__10202));
    ClkMux I__2384 (
            .O(N__10324),
            .I(N__10202));
    ClkMux I__2383 (
            .O(N__10323),
            .I(N__10202));
    ClkMux I__2382 (
            .O(N__10322),
            .I(N__10202));
    ClkMux I__2381 (
            .O(N__10321),
            .I(N__10202));
    ClkMux I__2380 (
            .O(N__10320),
            .I(N__10202));
    ClkMux I__2379 (
            .O(N__10319),
            .I(N__10202));
    ClkMux I__2378 (
            .O(N__10318),
            .I(N__10202));
    ClkMux I__2377 (
            .O(N__10317),
            .I(N__10202));
    ClkMux I__2376 (
            .O(N__10316),
            .I(N__10202));
    ClkMux I__2375 (
            .O(N__10315),
            .I(N__10202));
    ClkMux I__2374 (
            .O(N__10314),
            .I(N__10202));
    ClkMux I__2373 (
            .O(N__10313),
            .I(N__10202));
    ClkMux I__2372 (
            .O(N__10312),
            .I(N__10202));
    ClkMux I__2371 (
            .O(N__10311),
            .I(N__10202));
    ClkMux I__2370 (
            .O(N__10310),
            .I(N__10202));
    ClkMux I__2369 (
            .O(N__10309),
            .I(N__10202));
    ClkMux I__2368 (
            .O(N__10308),
            .I(N__10202));
    ClkMux I__2367 (
            .O(N__10307),
            .I(N__10202));
    ClkMux I__2366 (
            .O(N__10306),
            .I(N__10202));
    ClkMux I__2365 (
            .O(N__10305),
            .I(N__10202));
    ClkMux I__2364 (
            .O(N__10304),
            .I(N__10202));
    Glb2LocalMux I__2363 (
            .O(N__10301),
            .I(N__10202));
    ClkMux I__2362 (
            .O(N__10300),
            .I(N__10202));
    ClkMux I__2361 (
            .O(N__10299),
            .I(N__10202));
    ClkMux I__2360 (
            .O(N__10298),
            .I(N__10202));
    ClkMux I__2359 (
            .O(N__10297),
            .I(N__10202));
    ClkMux I__2358 (
            .O(N__10296),
            .I(N__10202));
    ClkMux I__2357 (
            .O(N__10295),
            .I(N__10202));
    ClkMux I__2356 (
            .O(N__10294),
            .I(N__10202));
    ClkMux I__2355 (
            .O(N__10293),
            .I(N__10202));
    GlobalMux I__2354 (
            .O(N__10202),
            .I(CLK80_PLL));
    CEMux I__2353 (
            .O(N__10199),
            .I(N__10194));
    CEMux I__2352 (
            .O(N__10198),
            .I(N__10191));
    CEMux I__2351 (
            .O(N__10197),
            .I(N__10187));
    LocalMux I__2350 (
            .O(N__10194),
            .I(N__10182));
    LocalMux I__2349 (
            .O(N__10191),
            .I(N__10182));
    CEMux I__2348 (
            .O(N__10190),
            .I(N__10179));
    LocalMux I__2347 (
            .O(N__10187),
            .I(N__10174));
    Span4Mux_v I__2346 (
            .O(N__10182),
            .I(N__10171));
    LocalMux I__2345 (
            .O(N__10179),
            .I(N__10168));
    CEMux I__2344 (
            .O(N__10178),
            .I(N__10165));
    CEMux I__2343 (
            .O(N__10177),
            .I(N__10162));
    Span4Mux_h I__2342 (
            .O(N__10174),
            .I(N__10159));
    Span4Mux_v I__2341 (
            .O(N__10171),
            .I(N__10152));
    Span4Mux_h I__2340 (
            .O(N__10168),
            .I(N__10152));
    LocalMux I__2339 (
            .O(N__10165),
            .I(N__10152));
    LocalMux I__2338 (
            .O(N__10162),
            .I(N__10149));
    Span4Mux_v I__2337 (
            .O(N__10159),
            .I(N__10146));
    Span4Mux_h I__2336 (
            .O(N__10152),
            .I(N__10143));
    Span4Mux_h I__2335 (
            .O(N__10149),
            .I(N__10140));
    Odrv4 I__2334 (
            .O(N__10146),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__2333 (
            .O(N__10143),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__2332 (
            .O(N__10140),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__2331 (
            .O(N__10133),
            .I(N__10127));
    InMux I__2330 (
            .O(N__10132),
            .I(N__10124));
    InMux I__2329 (
            .O(N__10131),
            .I(N__10121));
    InMux I__2328 (
            .O(N__10130),
            .I(N__10118));
    LocalMux I__2327 (
            .O(N__10127),
            .I(N__10111));
    LocalMux I__2326 (
            .O(N__10124),
            .I(N__10111));
    LocalMux I__2325 (
            .O(N__10121),
            .I(N__10111));
    LocalMux I__2324 (
            .O(N__10118),
            .I(N__10108));
    Span4Mux_v I__2323 (
            .O(N__10111),
            .I(N__10105));
    Span4Mux_v I__2322 (
            .O(N__10108),
            .I(N__10102));
    Sp12to4 I__2321 (
            .O(N__10105),
            .I(N__10099));
    Sp12to4 I__2320 (
            .O(N__10102),
            .I(N__10096));
    Span12Mux_h I__2319 (
            .O(N__10099),
            .I(N__10093));
    Odrv12 I__2318 (
            .O(N__10096),
            .I(DRA_c_5));
    Odrv12 I__2317 (
            .O(N__10093),
            .I(DRA_c_5));
    InMux I__2316 (
            .O(N__10088),
            .I(N__10085));
    LocalMux I__2315 (
            .O(N__10085),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2314 (
            .O(N__10082),
            .I(N__10074));
    InMux I__2313 (
            .O(N__10081),
            .I(N__10074));
    InMux I__2312 (
            .O(N__10080),
            .I(N__10071));
    InMux I__2311 (
            .O(N__10079),
            .I(N__10068));
    LocalMux I__2310 (
            .O(N__10074),
            .I(N__10065));
    LocalMux I__2309 (
            .O(N__10071),
            .I(N__10060));
    LocalMux I__2308 (
            .O(N__10068),
            .I(N__10060));
    Span4Mux_v I__2307 (
            .O(N__10065),
            .I(N__10057));
    Span12Mux_v I__2306 (
            .O(N__10060),
            .I(N__10052));
    Sp12to4 I__2305 (
            .O(N__10057),
            .I(N__10052));
    Span12Mux_h I__2304 (
            .O(N__10052),
            .I(N__10049));
    Odrv12 I__2303 (
            .O(N__10049),
            .I(DRA_c_4));
    InMux I__2302 (
            .O(N__10046),
            .I(N__10038));
    InMux I__2301 (
            .O(N__10045),
            .I(N__10038));
    InMux I__2300 (
            .O(N__10044),
            .I(N__10035));
    InMux I__2299 (
            .O(N__10043),
            .I(N__10032));
    LocalMux I__2298 (
            .O(N__10038),
            .I(N__10027));
    LocalMux I__2297 (
            .O(N__10035),
            .I(N__10027));
    LocalMux I__2296 (
            .O(N__10032),
            .I(N__10024));
    Span4Mux_v I__2295 (
            .O(N__10027),
            .I(N__10021));
    Span4Mux_v I__2294 (
            .O(N__10024),
            .I(N__10018));
    Sp12to4 I__2293 (
            .O(N__10021),
            .I(N__10015));
    Sp12to4 I__2292 (
            .O(N__10018),
            .I(N__10012));
    Span12Mux_h I__2291 (
            .O(N__10015),
            .I(N__10009));
    Odrv12 I__2290 (
            .O(N__10012),
            .I(DRA_c_3));
    Odrv12 I__2289 (
            .O(N__10009),
            .I(DRA_c_3));
    CascadeMux I__2288 (
            .O(N__10004),
            .I(N__10001));
    InMux I__2287 (
            .O(N__10001),
            .I(N__9998));
    LocalMux I__2286 (
            .O(N__9998),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2285 (
            .O(N__9995),
            .I(N__9992));
    LocalMux I__2284 (
            .O(N__9992),
            .I(N__9989));
    Span4Mux_h I__2283 (
            .O(N__9989),
            .I(N__9986));
    Odrv4 I__2282 (
            .O(N__9986),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__2281 (
            .O(N__9983),
            .I(N__9980));
    LocalMux I__2280 (
            .O(N__9980),
            .I(N__9977));
    Span4Mux_v I__2279 (
            .O(N__9977),
            .I(N__9974));
    Span4Mux_h I__2278 (
            .O(N__9974),
            .I(N__9971));
    Odrv4 I__2277 (
            .O(N__9971),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    CascadeMux I__2276 (
            .O(N__9968),
            .I(N__9965));
    InMux I__2275 (
            .O(N__9965),
            .I(N__9962));
    LocalMux I__2274 (
            .O(N__9962),
            .I(N__9959));
    Odrv12 I__2273 (
            .O(N__9959),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2272 (
            .O(N__9956),
            .I(N__9953));
    LocalMux I__2271 (
            .O(N__9953),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__2270 (
            .O(N__9950),
            .I(N__9947));
    LocalMux I__2269 (
            .O(N__9947),
            .I(N__9944));
    IoSpan4Mux I__2268 (
            .O(N__9944),
            .I(N__9941));
    Sp12to4 I__2267 (
            .O(N__9941),
            .I(N__9938));
    Span12Mux_s9_v I__2266 (
            .O(N__9938),
            .I(N__9935));
    Odrv12 I__2265 (
            .O(N__9935),
            .I(CMA_c_2));
    InMux I__2264 (
            .O(N__9932),
            .I(N__9929));
    LocalMux I__2263 (
            .O(N__9929),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__2262 (
            .O(N__9926),
            .I(N__9923));
    LocalMux I__2261 (
            .O(N__9923),
            .I(N__9920));
    Span4Mux_s1_h I__2260 (
            .O(N__9920),
            .I(N__9917));
    Sp12to4 I__2259 (
            .O(N__9917),
            .I(N__9914));
    Span12Mux_v I__2258 (
            .O(N__9914),
            .I(N__9911));
    Span12Mux_h I__2257 (
            .O(N__9911),
            .I(N__9908));
    Odrv12 I__2256 (
            .O(N__9908),
            .I(CMA_c_3));
    CascadeMux I__2255 (
            .O(N__9905),
            .I(N__9902));
    InMux I__2254 (
            .O(N__9902),
            .I(N__9899));
    LocalMux I__2253 (
            .O(N__9899),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2252 (
            .O(N__9896),
            .I(N__9893));
    LocalMux I__2251 (
            .O(N__9893),
            .I(N__9890));
    Span4Mux_h I__2250 (
            .O(N__9890),
            .I(N__9887));
    Odrv4 I__2249 (
            .O(N__9887),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__2248 (
            .O(N__9884),
            .I(N__9881));
    LocalMux I__2247 (
            .O(N__9881),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__2246 (
            .O(N__9878),
            .I(N__9875));
    LocalMux I__2245 (
            .O(N__9875),
            .I(N__9872));
    Odrv4 I__2244 (
            .O(N__9872),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__2243 (
            .O(N__9869),
            .I(N__9865));
    InMux I__2242 (
            .O(N__9868),
            .I(N__9860));
    LocalMux I__2241 (
            .O(N__9865),
            .I(N__9857));
    InMux I__2240 (
            .O(N__9864),
            .I(N__9853));
    CascadeMux I__2239 (
            .O(N__9863),
            .I(N__9850));
    LocalMux I__2238 (
            .O(N__9860),
            .I(N__9847));
    Sp12to4 I__2237 (
            .O(N__9857),
            .I(N__9844));
    InMux I__2236 (
            .O(N__9856),
            .I(N__9840));
    LocalMux I__2235 (
            .O(N__9853),
            .I(N__9836));
    InMux I__2234 (
            .O(N__9850),
            .I(N__9833));
    Span12Mux_h I__2233 (
            .O(N__9847),
            .I(N__9830));
    Span12Mux_v I__2232 (
            .O(N__9844),
            .I(N__9827));
    InMux I__2231 (
            .O(N__9843),
            .I(N__9824));
    LocalMux I__2230 (
            .O(N__9840),
            .I(N__9821));
    InMux I__2229 (
            .O(N__9839),
            .I(N__9818));
    Span4Mux_h I__2228 (
            .O(N__9836),
            .I(N__9815));
    LocalMux I__2227 (
            .O(N__9833),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv12 I__2226 (
            .O(N__9830),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv12 I__2225 (
            .O(N__9827),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__2224 (
            .O(N__9824),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__2223 (
            .O(N__9821),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__2222 (
            .O(N__9818),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__2221 (
            .O(N__9815),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__2220 (
            .O(N__9800),
            .I(N__9797));
    LocalMux I__2219 (
            .O(N__9797),
            .I(N__9794));
    Span4Mux_s3_h I__2218 (
            .O(N__9794),
            .I(N__9791));
    Span4Mux_v I__2217 (
            .O(N__9791),
            .I(N__9788));
    Span4Mux_h I__2216 (
            .O(N__9788),
            .I(N__9785));
    Span4Mux_h I__2215 (
            .O(N__9785),
            .I(N__9782));
    Odrv4 I__2214 (
            .O(N__9782),
            .I(WEn_c));
    InMux I__2213 (
            .O(N__9779),
            .I(N__9776));
    LocalMux I__2212 (
            .O(N__9776),
            .I(N__9772));
    InMux I__2211 (
            .O(N__9775),
            .I(N__9769));
    Span4Mux_v I__2210 (
            .O(N__9772),
            .I(N__9762));
    LocalMux I__2209 (
            .O(N__9769),
            .I(N__9762));
    InMux I__2208 (
            .O(N__9768),
            .I(N__9759));
    InMux I__2207 (
            .O(N__9767),
            .I(N__9753));
    Span4Mux_h I__2206 (
            .O(N__9762),
            .I(N__9750));
    LocalMux I__2205 (
            .O(N__9759),
            .I(N__9747));
    InMux I__2204 (
            .O(N__9758),
            .I(N__9744));
    InMux I__2203 (
            .O(N__9757),
            .I(N__9741));
    InMux I__2202 (
            .O(N__9756),
            .I(N__9738));
    LocalMux I__2201 (
            .O(N__9753),
            .I(N__9735));
    Span4Mux_v I__2200 (
            .O(N__9750),
            .I(N__9730));
    Span4Mux_h I__2199 (
            .O(N__9747),
            .I(N__9730));
    LocalMux I__2198 (
            .O(N__9744),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__2197 (
            .O(N__9741),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__2196 (
            .O(N__9738),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2195 (
            .O(N__9735),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2194 (
            .O(N__9730),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__2193 (
            .O(N__9719),
            .I(N__9716));
    LocalMux I__2192 (
            .O(N__9716),
            .I(N__9713));
    Span12Mux_s9_v I__2191 (
            .O(N__9713),
            .I(N__9710));
    Odrv12 I__2190 (
            .O(N__9710),
            .I(RASn_c));
    InMux I__2189 (
            .O(N__9707),
            .I(N__9700));
    InMux I__2188 (
            .O(N__9706),
            .I(N__9695));
    CascadeMux I__2187 (
            .O(N__9705),
            .I(N__9692));
    CascadeMux I__2186 (
            .O(N__9704),
            .I(N__9687));
    CascadeMux I__2185 (
            .O(N__9703),
            .I(N__9683));
    LocalMux I__2184 (
            .O(N__9700),
            .I(N__9680));
    InMux I__2183 (
            .O(N__9699),
            .I(N__9677));
    CascadeMux I__2182 (
            .O(N__9698),
            .I(N__9674));
    LocalMux I__2181 (
            .O(N__9695),
            .I(N__9671));
    InMux I__2180 (
            .O(N__9692),
            .I(N__9664));
    InMux I__2179 (
            .O(N__9691),
            .I(N__9664));
    CascadeMux I__2178 (
            .O(N__9690),
            .I(N__9661));
    InMux I__2177 (
            .O(N__9687),
            .I(N__9652));
    InMux I__2176 (
            .O(N__9686),
            .I(N__9652));
    InMux I__2175 (
            .O(N__9683),
            .I(N__9652));
    Span4Mux_v I__2174 (
            .O(N__9680),
            .I(N__9647));
    LocalMux I__2173 (
            .O(N__9677),
            .I(N__9647));
    InMux I__2172 (
            .O(N__9674),
            .I(N__9644));
    Span4Mux_v I__2171 (
            .O(N__9671),
            .I(N__9638));
    InMux I__2170 (
            .O(N__9670),
            .I(N__9633));
    InMux I__2169 (
            .O(N__9669),
            .I(N__9633));
    LocalMux I__2168 (
            .O(N__9664),
            .I(N__9630));
    InMux I__2167 (
            .O(N__9661),
            .I(N__9617));
    InMux I__2166 (
            .O(N__9660),
            .I(N__9617));
    InMux I__2165 (
            .O(N__9659),
            .I(N__9617));
    LocalMux I__2164 (
            .O(N__9652),
            .I(N__9612));
    Span4Mux_v I__2163 (
            .O(N__9647),
            .I(N__9612));
    LocalMux I__2162 (
            .O(N__9644),
            .I(N__9609));
    InMux I__2161 (
            .O(N__9643),
            .I(N__9602));
    InMux I__2160 (
            .O(N__9642),
            .I(N__9602));
    InMux I__2159 (
            .O(N__9641),
            .I(N__9602));
    Span4Mux_v I__2158 (
            .O(N__9638),
            .I(N__9597));
    LocalMux I__2157 (
            .O(N__9633),
            .I(N__9597));
    Span4Mux_h I__2156 (
            .O(N__9630),
            .I(N__9594));
    InMux I__2155 (
            .O(N__9629),
            .I(N__9589));
    InMux I__2154 (
            .O(N__9628),
            .I(N__9589));
    InMux I__2153 (
            .O(N__9627),
            .I(N__9582));
    InMux I__2152 (
            .O(N__9626),
            .I(N__9582));
    InMux I__2151 (
            .O(N__9625),
            .I(N__9582));
    InMux I__2150 (
            .O(N__9624),
            .I(N__9579));
    LocalMux I__2149 (
            .O(N__9617),
            .I(N__9576));
    Span4Mux_h I__2148 (
            .O(N__9612),
            .I(N__9571));
    Span4Mux_h I__2147 (
            .O(N__9609),
            .I(N__9571));
    LocalMux I__2146 (
            .O(N__9602),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2145 (
            .O(N__9597),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2144 (
            .O(N__9594),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2143 (
            .O(N__9589),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2142 (
            .O(N__9582),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2141 (
            .O(N__9579),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__2140 (
            .O(N__9576),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2139 (
            .O(N__9571),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__2138 (
            .O(N__9554),
            .I(N__9551));
    LocalMux I__2137 (
            .O(N__9551),
            .I(N__9548));
    Span12Mux_s10_v I__2136 (
            .O(N__9548),
            .I(N__9545));
    Odrv12 I__2135 (
            .O(N__9545),
            .I(CASn_c));
    CascadeMux I__2134 (
            .O(N__9542),
            .I(N__9538));
    InMux I__2133 (
            .O(N__9541),
            .I(N__9535));
    InMux I__2132 (
            .O(N__9538),
            .I(N__9532));
    LocalMux I__2131 (
            .O(N__9535),
            .I(N__9529));
    LocalMux I__2130 (
            .O(N__9532),
            .I(N__9526));
    Span4Mux_v I__2129 (
            .O(N__9529),
            .I(N__9523));
    Odrv12 I__2128 (
            .O(N__9526),
            .I(DBRn_c_i));
    Odrv4 I__2127 (
            .O(N__9523),
            .I(DBRn_c_i));
    InMux I__2126 (
            .O(N__9518),
            .I(N__9515));
    LocalMux I__2125 (
            .O(N__9515),
            .I(N__9511));
    InMux I__2124 (
            .O(N__9514),
            .I(N__9508));
    Span4Mux_h I__2123 (
            .O(N__9511),
            .I(N__9505));
    LocalMux I__2122 (
            .O(N__9508),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    Odrv4 I__2121 (
            .O(N__9505),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    InMux I__2120 (
            .O(N__9500),
            .I(N__9496));
    CascadeMux I__2119 (
            .O(N__9499),
            .I(N__9493));
    LocalMux I__2118 (
            .O(N__9496),
            .I(N__9490));
    InMux I__2117 (
            .O(N__9493),
            .I(N__9487));
    Span4Mux_v I__2116 (
            .O(N__9490),
            .I(N__9480));
    LocalMux I__2115 (
            .O(N__9487),
            .I(N__9480));
    CascadeMux I__2114 (
            .O(N__9486),
            .I(N__9477));
    InMux I__2113 (
            .O(N__9485),
            .I(N__9474));
    Span4Mux_h I__2112 (
            .O(N__9480),
            .I(N__9471));
    InMux I__2111 (
            .O(N__9477),
            .I(N__9468));
    LocalMux I__2110 (
            .O(N__9474),
            .I(N__9465));
    Span4Mux_v I__2109 (
            .O(N__9471),
            .I(N__9458));
    LocalMux I__2108 (
            .O(N__9468),
            .I(N__9458));
    Span4Mux_h I__2107 (
            .O(N__9465),
            .I(N__9458));
    Odrv4 I__2106 (
            .O(N__9458),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__2105 (
            .O(N__9455),
            .I(N__9452));
    LocalMux I__2104 (
            .O(N__9452),
            .I(N__9449));
    Span4Mux_s3_v I__2103 (
            .O(N__9449),
            .I(N__9446));
    Span4Mux_v I__2102 (
            .O(N__9446),
            .I(N__9443));
    Span4Mux_h I__2101 (
            .O(N__9443),
            .I(N__9440));
    Odrv4 I__2100 (
            .O(N__9440),
            .I(CRCSn_c));
    InMux I__2099 (
            .O(N__9437),
            .I(N__9433));
    InMux I__2098 (
            .O(N__9436),
            .I(N__9430));
    LocalMux I__2097 (
            .O(N__9433),
            .I(N__9424));
    LocalMux I__2096 (
            .O(N__9430),
            .I(N__9424));
    CascadeMux I__2095 (
            .O(N__9429),
            .I(N__9421));
    Span4Mux_h I__2094 (
            .O(N__9424),
            .I(N__9417));
    InMux I__2093 (
            .O(N__9421),
            .I(N__9412));
    InMux I__2092 (
            .O(N__9420),
            .I(N__9412));
    Span4Mux_v I__2091 (
            .O(N__9417),
            .I(N__9409));
    LocalMux I__2090 (
            .O(N__9412),
            .I(N__9406));
    Odrv4 I__2089 (
            .O(N__9409),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    Odrv12 I__2088 (
            .O(N__9406),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    InMux I__2087 (
            .O(N__9401),
            .I(N__9398));
    LocalMux I__2086 (
            .O(N__9398),
            .I(N__9395));
    Sp12to4 I__2085 (
            .O(N__9395),
            .I(N__9392));
    Span12Mux_v I__2084 (
            .O(N__9392),
            .I(N__9389));
    Span12Mux_h I__2083 (
            .O(N__9389),
            .I(N__9386));
    Odrv12 I__2082 (
            .O(N__9386),
            .I(A_c_19));
    IoInMux I__2081 (
            .O(N__9383),
            .I(N__9380));
    LocalMux I__2080 (
            .O(N__9380),
            .I(N__9377));
    IoSpan4Mux I__2079 (
            .O(N__9377),
            .I(N__9374));
    Span4Mux_s2_h I__2078 (
            .O(N__9374),
            .I(N__9371));
    Span4Mux_v I__2077 (
            .O(N__9371),
            .I(N__9368));
    Sp12to4 I__2076 (
            .O(N__9368),
            .I(N__9365));
    Odrv12 I__2075 (
            .O(N__9365),
            .I(CMA_c_9));
    InMux I__2074 (
            .O(N__9362),
            .I(N__9359));
    LocalMux I__2073 (
            .O(N__9359),
            .I(N__9356));
    Odrv4 I__2072 (
            .O(N__9356),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    InMux I__2071 (
            .O(N__9353),
            .I(N__9350));
    LocalMux I__2070 (
            .O(N__9350),
            .I(N__9347));
    Odrv4 I__2069 (
            .O(N__9347),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    CascadeMux I__2068 (
            .O(N__9344),
            .I(N__9334));
    CascadeMux I__2067 (
            .O(N__9343),
            .I(N__9328));
    CascadeMux I__2066 (
            .O(N__9342),
            .I(N__9325));
    CascadeMux I__2065 (
            .O(N__9341),
            .I(N__9321));
    CascadeMux I__2064 (
            .O(N__9340),
            .I(N__9318));
    CascadeMux I__2063 (
            .O(N__9339),
            .I(N__9315));
    CascadeMux I__2062 (
            .O(N__9338),
            .I(N__9310));
    InMux I__2061 (
            .O(N__9337),
            .I(N__9300));
    InMux I__2060 (
            .O(N__9334),
            .I(N__9296));
    InMux I__2059 (
            .O(N__9333),
            .I(N__9293));
    InMux I__2058 (
            .O(N__9332),
            .I(N__9288));
    InMux I__2057 (
            .O(N__9331),
            .I(N__9288));
    InMux I__2056 (
            .O(N__9328),
            .I(N__9285));
    InMux I__2055 (
            .O(N__9325),
            .I(N__9274));
    InMux I__2054 (
            .O(N__9324),
            .I(N__9274));
    InMux I__2053 (
            .O(N__9321),
            .I(N__9274));
    InMux I__2052 (
            .O(N__9318),
            .I(N__9274));
    InMux I__2051 (
            .O(N__9315),
            .I(N__9274));
    InMux I__2050 (
            .O(N__9314),
            .I(N__9271));
    InMux I__2049 (
            .O(N__9313),
            .I(N__9268));
    InMux I__2048 (
            .O(N__9310),
            .I(N__9265));
    InMux I__2047 (
            .O(N__9309),
            .I(N__9258));
    InMux I__2046 (
            .O(N__9308),
            .I(N__9258));
    InMux I__2045 (
            .O(N__9307),
            .I(N__9258));
    InMux I__2044 (
            .O(N__9306),
            .I(N__9251));
    InMux I__2043 (
            .O(N__9305),
            .I(N__9251));
    InMux I__2042 (
            .O(N__9304),
            .I(N__9251));
    InMux I__2041 (
            .O(N__9303),
            .I(N__9246));
    LocalMux I__2040 (
            .O(N__9300),
            .I(N__9243));
    InMux I__2039 (
            .O(N__9299),
            .I(N__9240));
    LocalMux I__2038 (
            .O(N__9296),
            .I(N__9237));
    LocalMux I__2037 (
            .O(N__9293),
            .I(N__9234));
    LocalMux I__2036 (
            .O(N__9288),
            .I(N__9225));
    LocalMux I__2035 (
            .O(N__9285),
            .I(N__9225));
    LocalMux I__2034 (
            .O(N__9274),
            .I(N__9225));
    LocalMux I__2033 (
            .O(N__9271),
            .I(N__9225));
    LocalMux I__2032 (
            .O(N__9268),
            .I(N__9222));
    LocalMux I__2031 (
            .O(N__9265),
            .I(N__9219));
    LocalMux I__2030 (
            .O(N__9258),
            .I(N__9214));
    LocalMux I__2029 (
            .O(N__9251),
            .I(N__9214));
    InMux I__2028 (
            .O(N__9250),
            .I(N__9211));
    InMux I__2027 (
            .O(N__9249),
            .I(N__9208));
    LocalMux I__2026 (
            .O(N__9246),
            .I(N__9205));
    Span4Mux_v I__2025 (
            .O(N__9243),
            .I(N__9194));
    LocalMux I__2024 (
            .O(N__9240),
            .I(N__9194));
    Span4Mux_v I__2023 (
            .O(N__9237),
            .I(N__9194));
    Span4Mux_h I__2022 (
            .O(N__9234),
            .I(N__9194));
    Span4Mux_v I__2021 (
            .O(N__9225),
            .I(N__9194));
    Span4Mux_v I__2020 (
            .O(N__9222),
            .I(N__9187));
    Span4Mux_h I__2019 (
            .O(N__9219),
            .I(N__9187));
    Span4Mux_h I__2018 (
            .O(N__9214),
            .I(N__9187));
    LocalMux I__2017 (
            .O(N__9211),
            .I(N__9184));
    LocalMux I__2016 (
            .O(N__9208),
            .I(CPU_CYCLEm));
    Odrv4 I__2015 (
            .O(N__9205),
            .I(CPU_CYCLEm));
    Odrv4 I__2014 (
            .O(N__9194),
            .I(CPU_CYCLEm));
    Odrv4 I__2013 (
            .O(N__9187),
            .I(CPU_CYCLEm));
    Odrv12 I__2012 (
            .O(N__9184),
            .I(CPU_CYCLEm));
    InMux I__2011 (
            .O(N__9173),
            .I(N__9170));
    LocalMux I__2010 (
            .O(N__9170),
            .I(N__9167));
    Odrv4 I__2009 (
            .O(N__9167),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__2008 (
            .O(N__9164),
            .I(N__9161));
    LocalMux I__2007 (
            .O(N__9161),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__2006 (
            .O(N__9158),
            .I(N__9155));
    LocalMux I__2005 (
            .O(N__9155),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2004 (
            .O(N__9152),
            .I(N__9149));
    LocalMux I__2003 (
            .O(N__9149),
            .I(N__9146));
    Odrv4 I__2002 (
            .O(N__9146),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    IoInMux I__2001 (
            .O(N__9143),
            .I(N__9140));
    LocalMux I__2000 (
            .O(N__9140),
            .I(N__9137));
    Span4Mux_s1_v I__1999 (
            .O(N__9137),
            .I(N__9134));
    Sp12to4 I__1998 (
            .O(N__9134),
            .I(N__9131));
    Span12Mux_h I__1997 (
            .O(N__9131),
            .I(N__9128));
    Span12Mux_v I__1996 (
            .O(N__9128),
            .I(N__9125));
    Odrv12 I__1995 (
            .O(N__9125),
            .I(CMA_c_0));
    InMux I__1994 (
            .O(N__9122),
            .I(N__9119));
    LocalMux I__1993 (
            .O(N__9119),
            .I(N__9116));
    Span4Mux_v I__1992 (
            .O(N__9116),
            .I(N__9113));
    Span4Mux_v I__1991 (
            .O(N__9113),
            .I(N__9110));
    Sp12to4 I__1990 (
            .O(N__9110),
            .I(N__9107));
    Span12Mux_h I__1989 (
            .O(N__9107),
            .I(N__9104));
    Odrv12 I__1988 (
            .O(N__9104),
            .I(A_c_17));
    IoInMux I__1987 (
            .O(N__9101),
            .I(N__9098));
    LocalMux I__1986 (
            .O(N__9098),
            .I(N__9095));
    IoSpan4Mux I__1985 (
            .O(N__9095),
            .I(N__9092));
    IoSpan4Mux I__1984 (
            .O(N__9092),
            .I(N__9089));
    Sp12to4 I__1983 (
            .O(N__9089),
            .I(N__9086));
    Span12Mux_s9_h I__1982 (
            .O(N__9086),
            .I(N__9083));
    Odrv12 I__1981 (
            .O(N__9083),
            .I(CMA_c_8));
    InMux I__1980 (
            .O(N__9080),
            .I(N__9077));
    LocalMux I__1979 (
            .O(N__9077),
            .I(N__9074));
    Odrv4 I__1978 (
            .O(N__9074),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    CascadeMux I__1977 (
            .O(N__9071),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_ ));
    InMux I__1976 (
            .O(N__9068),
            .I(N__9065));
    LocalMux I__1975 (
            .O(N__9065),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    IoInMux I__1974 (
            .O(N__9062),
            .I(N__9059));
    LocalMux I__1973 (
            .O(N__9059),
            .I(N__9056));
    Span12Mux_s2_h I__1972 (
            .O(N__9056),
            .I(N__9053));
    Span12Mux_h I__1971 (
            .O(N__9053),
            .I(N__9050));
    Span12Mux_v I__1970 (
            .O(N__9050),
            .I(N__9047));
    Odrv12 I__1969 (
            .O(N__9047),
            .I(CMA_c_5));
    InMux I__1968 (
            .O(N__9044),
            .I(N__9038));
    InMux I__1967 (
            .O(N__9043),
            .I(N__9038));
    LocalMux I__1966 (
            .O(N__9038),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1965 (
            .O(N__9035),
            .I(N__9032));
    LocalMux I__1964 (
            .O(N__9032),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__1963 (
            .O(N__9029),
            .I(N__9026));
    LocalMux I__1962 (
            .O(N__9026),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    InMux I__1961 (
            .O(N__9023),
            .I(N__9020));
    LocalMux I__1960 (
            .O(N__9020),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    CascadeMux I__1959 (
            .O(N__9017),
            .I(\U712_CHIP_RAM.N_11_cascade_ ));
    InMux I__1958 (
            .O(N__9014),
            .I(N__9011));
    LocalMux I__1957 (
            .O(N__9011),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    InMux I__1956 (
            .O(N__9008),
            .I(N__9005));
    LocalMux I__1955 (
            .O(N__9005),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ));
    IoInMux I__1954 (
            .O(N__9002),
            .I(N__8999));
    LocalMux I__1953 (
            .O(N__8999),
            .I(N__8996));
    IoSpan4Mux I__1952 (
            .O(N__8996),
            .I(N__8993));
    Span4Mux_s2_v I__1951 (
            .O(N__8993),
            .I(N__8988));
    InMux I__1950 (
            .O(N__8992),
            .I(N__8983));
    InMux I__1949 (
            .O(N__8991),
            .I(N__8983));
    Sp12to4 I__1948 (
            .O(N__8988),
            .I(N__8980));
    LocalMux I__1947 (
            .O(N__8983),
            .I(N__8977));
    Span12Mux_s8_v I__1946 (
            .O(N__8980),
            .I(N__8972));
    Sp12to4 I__1945 (
            .O(N__8977),
            .I(N__8972));
    Span12Mux_v I__1944 (
            .O(N__8972),
            .I(N__8969));
    Span12Mux_h I__1943 (
            .O(N__8969),
            .I(N__8966));
    Odrv12 I__1942 (
            .O(N__8966),
            .I(A_c_10));
    InMux I__1941 (
            .O(N__8963),
            .I(N__8960));
    LocalMux I__1940 (
            .O(N__8960),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    InMux I__1939 (
            .O(N__8957),
            .I(N__8954));
    LocalMux I__1938 (
            .O(N__8954),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    InMux I__1937 (
            .O(N__8951),
            .I(N__8948));
    LocalMux I__1936 (
            .O(N__8948),
            .I(N__8945));
    Span4Mux_v I__1935 (
            .O(N__8945),
            .I(N__8942));
    Sp12to4 I__1934 (
            .O(N__8942),
            .I(N__8939));
    Span12Mux_h I__1933 (
            .O(N__8939),
            .I(N__8936));
    Odrv12 I__1932 (
            .O(N__8936),
            .I(A_c_5));
    InMux I__1931 (
            .O(N__8933),
            .I(N__8930));
    LocalMux I__1930 (
            .O(N__8930),
            .I(N__8927));
    Sp12to4 I__1929 (
            .O(N__8927),
            .I(N__8924));
    Span12Mux_v I__1928 (
            .O(N__8924),
            .I(N__8921));
    Span12Mux_h I__1927 (
            .O(N__8921),
            .I(N__8918));
    Odrv12 I__1926 (
            .O(N__8918),
            .I(A_c_12));
    InMux I__1925 (
            .O(N__8915),
            .I(N__8912));
    LocalMux I__1924 (
            .O(N__8912),
            .I(N__8909));
    Span4Mux_v I__1923 (
            .O(N__8909),
            .I(N__8906));
    Sp12to4 I__1922 (
            .O(N__8906),
            .I(N__8903));
    Span12Mux_h I__1921 (
            .O(N__8903),
            .I(N__8900));
    Odrv12 I__1920 (
            .O(N__8900),
            .I(A_c_4));
    IoInMux I__1919 (
            .O(N__8897),
            .I(N__8894));
    LocalMux I__1918 (
            .O(N__8894),
            .I(N__8891));
    IoSpan4Mux I__1917 (
            .O(N__8891),
            .I(N__8887));
    InMux I__1916 (
            .O(N__8890),
            .I(N__8884));
    Span4Mux_s2_v I__1915 (
            .O(N__8887),
            .I(N__8881));
    LocalMux I__1914 (
            .O(N__8884),
            .I(N__8878));
    Sp12to4 I__1913 (
            .O(N__8881),
            .I(N__8875));
    Span4Mux_v I__1912 (
            .O(N__8878),
            .I(N__8872));
    Span12Mux_s8_v I__1911 (
            .O(N__8875),
            .I(N__8869));
    Span4Mux_v I__1910 (
            .O(N__8872),
            .I(N__8866));
    Span12Mux_h I__1909 (
            .O(N__8869),
            .I(N__8863));
    Sp12to4 I__1908 (
            .O(N__8866),
            .I(N__8860));
    Span12Mux_v I__1907 (
            .O(N__8863),
            .I(N__8857));
    Span12Mux_h I__1906 (
            .O(N__8860),
            .I(N__8854));
    Odrv12 I__1905 (
            .O(N__8857),
            .I(A_c_11));
    Odrv12 I__1904 (
            .O(N__8854),
            .I(A_c_11));
    IoInMux I__1903 (
            .O(N__8849),
            .I(N__8846));
    LocalMux I__1902 (
            .O(N__8846),
            .I(N__8843));
    Span12Mux_s11_v I__1901 (
            .O(N__8843),
            .I(N__8840));
    Odrv12 I__1900 (
            .O(N__8840),
            .I(CMA_c_10));
    IoInMux I__1899 (
            .O(N__8837),
            .I(N__8834));
    LocalMux I__1898 (
            .O(N__8834),
            .I(N__8831));
    Span4Mux_s3_v I__1897 (
            .O(N__8831),
            .I(N__8827));
    InMux I__1896 (
            .O(N__8830),
            .I(N__8824));
    Span4Mux_v I__1895 (
            .O(N__8827),
            .I(N__8821));
    LocalMux I__1894 (
            .O(N__8824),
            .I(N__8818));
    Sp12to4 I__1893 (
            .O(N__8821),
            .I(N__8815));
    Span4Mux_v I__1892 (
            .O(N__8818),
            .I(N__8812));
    Span12Mux_h I__1891 (
            .O(N__8815),
            .I(N__8809));
    Span4Mux_v I__1890 (
            .O(N__8812),
            .I(N__8806));
    Odrv12 I__1889 (
            .O(N__8809),
            .I(UMBEn_c));
    Odrv4 I__1888 (
            .O(N__8806),
            .I(UMBEn_c));
    CascadeMux I__1887 (
            .O(N__8801),
            .I(\U712_BYTE_ENABLE.un3_CUMBEnZ0Z_1_cascade_ ));
    IoInMux I__1886 (
            .O(N__8798),
            .I(N__8795));
    LocalMux I__1885 (
            .O(N__8795),
            .I(N__8792));
    Span12Mux_s3_h I__1884 (
            .O(N__8792),
            .I(N__8789));
    Span12Mux_h I__1883 (
            .O(N__8789),
            .I(N__8786));
    Span12Mux_v I__1882 (
            .O(N__8786),
            .I(N__8783));
    Odrv12 I__1881 (
            .O(N__8783),
            .I(CUMBEn_c));
    InMux I__1880 (
            .O(N__8780),
            .I(N__8776));
    IoInMux I__1879 (
            .O(N__8779),
            .I(N__8773));
    LocalMux I__1878 (
            .O(N__8776),
            .I(N__8770));
    LocalMux I__1877 (
            .O(N__8773),
            .I(N__8767));
    Span4Mux_v I__1876 (
            .O(N__8770),
            .I(N__8764));
    Span12Mux_s9_v I__1875 (
            .O(N__8767),
            .I(N__8761));
    Span4Mux_v I__1874 (
            .O(N__8764),
            .I(N__8758));
    Odrv12 I__1873 (
            .O(N__8761),
            .I(UUBEn_c));
    Odrv4 I__1872 (
            .O(N__8758),
            .I(UUBEn_c));
    CascadeMux I__1871 (
            .O(N__8753),
            .I(N__8750));
    InMux I__1870 (
            .O(N__8750),
            .I(N__8747));
    LocalMux I__1869 (
            .O(N__8747),
            .I(\U712_BYTE_ENABLE.un3_CUMBEnZ0Z_1 ));
    IoInMux I__1868 (
            .O(N__8744),
            .I(N__8741));
    LocalMux I__1867 (
            .O(N__8741),
            .I(N__8738));
    Span4Mux_s3_h I__1866 (
            .O(N__8738),
            .I(N__8735));
    Sp12to4 I__1865 (
            .O(N__8735),
            .I(N__8732));
    Span12Mux_v I__1864 (
            .O(N__8732),
            .I(N__8729));
    Span12Mux_h I__1863 (
            .O(N__8729),
            .I(N__8726));
    Odrv12 I__1862 (
            .O(N__8726),
            .I(CUUBEn_c));
    IoInMux I__1861 (
            .O(N__8723),
            .I(N__8720));
    LocalMux I__1860 (
            .O(N__8720),
            .I(N__8715));
    InMux I__1859 (
            .O(N__8719),
            .I(N__8710));
    InMux I__1858 (
            .O(N__8718),
            .I(N__8710));
    Span12Mux_s2_v I__1857 (
            .O(N__8715),
            .I(N__8707));
    LocalMux I__1856 (
            .O(N__8710),
            .I(N__8704));
    Span12Mux_v I__1855 (
            .O(N__8707),
            .I(N__8700));
    Span4Mux_v I__1854 (
            .O(N__8704),
            .I(N__8697));
    InMux I__1853 (
            .O(N__8703),
            .I(N__8694));
    Odrv12 I__1852 (
            .O(N__8700),
            .I(DBENn_c));
    Odrv4 I__1851 (
            .O(N__8697),
            .I(DBENn_c));
    LocalMux I__1850 (
            .O(N__8694),
            .I(DBENn_c));
    InMux I__1849 (
            .O(N__8687),
            .I(N__8683));
    InMux I__1848 (
            .O(N__8686),
            .I(N__8680));
    LocalMux I__1847 (
            .O(N__8683),
            .I(N__8675));
    LocalMux I__1846 (
            .O(N__8680),
            .I(N__8672));
    InMux I__1845 (
            .O(N__8679),
            .I(N__8667));
    InMux I__1844 (
            .O(N__8678),
            .I(N__8667));
    Span4Mux_v I__1843 (
            .O(N__8675),
            .I(N__8664));
    Span4Mux_h I__1842 (
            .O(N__8672),
            .I(N__8661));
    LocalMux I__1841 (
            .O(N__8667),
            .I(DMA_CYCLEm));
    Odrv4 I__1840 (
            .O(N__8664),
            .I(DMA_CYCLEm));
    Odrv4 I__1839 (
            .O(N__8661),
            .I(DMA_CYCLEm));
    InMux I__1838 (
            .O(N__8654),
            .I(N__8651));
    LocalMux I__1837 (
            .O(N__8651),
            .I(N__8648));
    Odrv4 I__1836 (
            .O(N__8648),
            .I(\U712_BYTE_ENABLE.un3_CLLBEnZ0Z_0 ));
    InMux I__1835 (
            .O(N__8645),
            .I(N__8642));
    LocalMux I__1834 (
            .O(N__8642),
            .I(N__8639));
    Span4Mux_v I__1833 (
            .O(N__8639),
            .I(N__8636));
    Span4Mux_v I__1832 (
            .O(N__8636),
            .I(N__8633));
    Odrv4 I__1831 (
            .O(N__8633),
            .I(\U712_BYTE_ENABLE.N_56 ));
    CascadeMux I__1830 (
            .O(N__8630),
            .I(\U712_BYTE_ENABLE.un3_CLLBEnZ0Z_0_cascade_ ));
    IoInMux I__1829 (
            .O(N__8627),
            .I(N__8624));
    LocalMux I__1828 (
            .O(N__8624),
            .I(N__8621));
    IoSpan4Mux I__1827 (
            .O(N__8621),
            .I(N__8618));
    Span4Mux_s2_v I__1826 (
            .O(N__8618),
            .I(N__8615));
    Sp12to4 I__1825 (
            .O(N__8615),
            .I(N__8612));
    Span12Mux_v I__1824 (
            .O(N__8612),
            .I(N__8609));
    Odrv12 I__1823 (
            .O(N__8609),
            .I(CLLBEn_c));
    IoInMux I__1822 (
            .O(N__8606),
            .I(N__8603));
    LocalMux I__1821 (
            .O(N__8603),
            .I(N__8600));
    IoSpan4Mux I__1820 (
            .O(N__8600),
            .I(N__8597));
    Span4Mux_s2_v I__1819 (
            .O(N__8597),
            .I(N__8594));
    Sp12to4 I__1818 (
            .O(N__8594),
            .I(N__8591));
    Span12Mux_s11_v I__1817 (
            .O(N__8591),
            .I(N__8588));
    Odrv12 I__1816 (
            .O(N__8588),
            .I(CMA_c_1));
    InMux I__1815 (
            .O(N__8585),
            .I(N__8582));
    LocalMux I__1814 (
            .O(N__8582),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    InMux I__1813 (
            .O(N__8579),
            .I(N__8576));
    LocalMux I__1812 (
            .O(N__8576),
            .I(N__8573));
    Span4Mux_v I__1811 (
            .O(N__8573),
            .I(N__8570));
    Span4Mux_v I__1810 (
            .O(N__8570),
            .I(N__8567));
    Sp12to4 I__1809 (
            .O(N__8567),
            .I(N__8564));
    Span12Mux_h I__1808 (
            .O(N__8564),
            .I(N__8561));
    Odrv12 I__1807 (
            .O(N__8561),
            .I(A_c_3));
    InMux I__1806 (
            .O(N__8558),
            .I(N__8555));
    LocalMux I__1805 (
            .O(N__8555),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER17_1_0 ));
    InMux I__1804 (
            .O(N__8552),
            .I(N__8548));
    InMux I__1803 (
            .O(N__8551),
            .I(N__8545));
    LocalMux I__1802 (
            .O(N__8548),
            .I(N__8540));
    LocalMux I__1801 (
            .O(N__8545),
            .I(N__8540));
    Odrv4 I__1800 (
            .O(N__8540),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa ));
    CascadeMux I__1799 (
            .O(N__8537),
            .I(\U712_CHIP_RAM.N_38_cascade_ ));
    InMux I__1798 (
            .O(N__8534),
            .I(N__8531));
    LocalMux I__1797 (
            .O(N__8531),
            .I(\U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa ));
    InMux I__1796 (
            .O(N__8528),
            .I(N__8525));
    LocalMux I__1795 (
            .O(N__8525),
            .I(N__8522));
    Span4Mux_h I__1794 (
            .O(N__8522),
            .I(N__8519));
    Odrv4 I__1793 (
            .O(N__8519),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_i_1_1 ));
    CascadeMux I__1792 (
            .O(N__8516),
            .I(N__8512));
    InMux I__1791 (
            .O(N__8515),
            .I(N__8509));
    InMux I__1790 (
            .O(N__8512),
            .I(N__8506));
    LocalMux I__1789 (
            .O(N__8509),
            .I(\U712_CHIP_RAM.N_151 ));
    LocalMux I__1788 (
            .O(N__8506),
            .I(\U712_CHIP_RAM.N_151 ));
    InMux I__1787 (
            .O(N__8501),
            .I(N__8495));
    InMux I__1786 (
            .O(N__8500),
            .I(N__8495));
    LocalMux I__1785 (
            .O(N__8495),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER19_0 ));
    CEMux I__1784 (
            .O(N__8492),
            .I(N__8489));
    LocalMux I__1783 (
            .O(N__8489),
            .I(N__8486));
    Span4Mux_v I__1782 (
            .O(N__8486),
            .I(N__8483));
    Span4Mux_h I__1781 (
            .O(N__8483),
            .I(N__8480));
    Odrv4 I__1780 (
            .O(N__8480),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_i ));
    InMux I__1779 (
            .O(N__8477),
            .I(N__8468));
    InMux I__1778 (
            .O(N__8476),
            .I(N__8460));
    InMux I__1777 (
            .O(N__8475),
            .I(N__8460));
    CascadeMux I__1776 (
            .O(N__8474),
            .I(N__8454));
    InMux I__1775 (
            .O(N__8473),
            .I(N__8449));
    InMux I__1774 (
            .O(N__8472),
            .I(N__8449));
    InMux I__1773 (
            .O(N__8471),
            .I(N__8445));
    LocalMux I__1772 (
            .O(N__8468),
            .I(N__8442));
    InMux I__1771 (
            .O(N__8467),
            .I(N__8439));
    InMux I__1770 (
            .O(N__8466),
            .I(N__8436));
    InMux I__1769 (
            .O(N__8465),
            .I(N__8433));
    LocalMux I__1768 (
            .O(N__8460),
            .I(N__8430));
    InMux I__1767 (
            .O(N__8459),
            .I(N__8425));
    InMux I__1766 (
            .O(N__8458),
            .I(N__8425));
    InMux I__1765 (
            .O(N__8457),
            .I(N__8420));
    InMux I__1764 (
            .O(N__8454),
            .I(N__8420));
    LocalMux I__1763 (
            .O(N__8449),
            .I(N__8417));
    InMux I__1762 (
            .O(N__8448),
            .I(N__8414));
    LocalMux I__1761 (
            .O(N__8445),
            .I(\U712_CHIP_RAM.N_331_3 ));
    Odrv4 I__1760 (
            .O(N__8442),
            .I(\U712_CHIP_RAM.N_331_3 ));
    LocalMux I__1759 (
            .O(N__8439),
            .I(\U712_CHIP_RAM.N_331_3 ));
    LocalMux I__1758 (
            .O(N__8436),
            .I(\U712_CHIP_RAM.N_331_3 ));
    LocalMux I__1757 (
            .O(N__8433),
            .I(\U712_CHIP_RAM.N_331_3 ));
    Odrv4 I__1756 (
            .O(N__8430),
            .I(\U712_CHIP_RAM.N_331_3 ));
    LocalMux I__1755 (
            .O(N__8425),
            .I(\U712_CHIP_RAM.N_331_3 ));
    LocalMux I__1754 (
            .O(N__8420),
            .I(\U712_CHIP_RAM.N_331_3 ));
    Odrv4 I__1753 (
            .O(N__8417),
            .I(\U712_CHIP_RAM.N_331_3 ));
    LocalMux I__1752 (
            .O(N__8414),
            .I(\U712_CHIP_RAM.N_331_3 ));
    InMux I__1751 (
            .O(N__8393),
            .I(N__8390));
    LocalMux I__1750 (
            .O(N__8390),
            .I(N__8387));
    Span4Mux_h I__1749 (
            .O(N__8387),
            .I(N__8384));
    Odrv4 I__1748 (
            .O(N__8384),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_29_i_a2_i_1 ));
    CascadeMux I__1747 (
            .O(N__8381),
            .I(\U712_CHIP_RAM.N_61_cascade_ ));
    InMux I__1746 (
            .O(N__8378),
            .I(N__8372));
    InMux I__1745 (
            .O(N__8377),
            .I(N__8372));
    LocalMux I__1744 (
            .O(N__8372),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1 ));
    InMux I__1743 (
            .O(N__8369),
            .I(N__8366));
    LocalMux I__1742 (
            .O(N__8366),
            .I(\U712_CHIP_RAM.N_218 ));
    InMux I__1741 (
            .O(N__8363),
            .I(N__8357));
    InMux I__1740 (
            .O(N__8362),
            .I(N__8357));
    LocalMux I__1739 (
            .O(N__8357),
            .I(N__8353));
    InMux I__1738 (
            .O(N__8356),
            .I(N__8350));
    Span4Mux_h I__1737 (
            .O(N__8353),
            .I(N__8345));
    LocalMux I__1736 (
            .O(N__8350),
            .I(N__8345));
    Odrv4 I__1735 (
            .O(N__8345),
            .I(\U712_CHIP_RAM.N_154 ));
    InMux I__1734 (
            .O(N__8342),
            .I(N__8339));
    LocalMux I__1733 (
            .O(N__8339),
            .I(N__8334));
    InMux I__1732 (
            .O(N__8338),
            .I(N__8331));
    InMux I__1731 (
            .O(N__8337),
            .I(N__8323));
    Span4Mux_v I__1730 (
            .O(N__8334),
            .I(N__8315));
    LocalMux I__1729 (
            .O(N__8331),
            .I(N__8312));
    InMux I__1728 (
            .O(N__8330),
            .I(N__8307));
    InMux I__1727 (
            .O(N__8329),
            .I(N__8307));
    InMux I__1726 (
            .O(N__8328),
            .I(N__8304));
    CascadeMux I__1725 (
            .O(N__8327),
            .I(N__8298));
    InMux I__1724 (
            .O(N__8326),
            .I(N__8294));
    LocalMux I__1723 (
            .O(N__8323),
            .I(N__8291));
    InMux I__1722 (
            .O(N__8322),
            .I(N__8286));
    InMux I__1721 (
            .O(N__8321),
            .I(N__8286));
    InMux I__1720 (
            .O(N__8320),
            .I(N__8279));
    InMux I__1719 (
            .O(N__8319),
            .I(N__8279));
    InMux I__1718 (
            .O(N__8318),
            .I(N__8279));
    Span4Mux_h I__1717 (
            .O(N__8315),
            .I(N__8272));
    Span4Mux_v I__1716 (
            .O(N__8312),
            .I(N__8272));
    LocalMux I__1715 (
            .O(N__8307),
            .I(N__8272));
    LocalMux I__1714 (
            .O(N__8304),
            .I(N__8269));
    InMux I__1713 (
            .O(N__8303),
            .I(N__8266));
    InMux I__1712 (
            .O(N__8302),
            .I(N__8257));
    InMux I__1711 (
            .O(N__8301),
            .I(N__8257));
    InMux I__1710 (
            .O(N__8298),
            .I(N__8257));
    InMux I__1709 (
            .O(N__8297),
            .I(N__8257));
    LocalMux I__1708 (
            .O(N__8294),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1707 (
            .O(N__8291),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1706 (
            .O(N__8286),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1705 (
            .O(N__8279),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1704 (
            .O(N__8272),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1703 (
            .O(N__8269),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1702 (
            .O(N__8266),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1701 (
            .O(N__8257),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__1700 (
            .O(N__8240),
            .I(N__8235));
    InMux I__1699 (
            .O(N__8239),
            .I(N__8231));
    CascadeMux I__1698 (
            .O(N__8238),
            .I(N__8228));
    LocalMux I__1697 (
            .O(N__8235),
            .I(N__8221));
    CascadeMux I__1696 (
            .O(N__8234),
            .I(N__8216));
    LocalMux I__1695 (
            .O(N__8231),
            .I(N__8209));
    InMux I__1694 (
            .O(N__8228),
            .I(N__8204));
    InMux I__1693 (
            .O(N__8227),
            .I(N__8204));
    InMux I__1692 (
            .O(N__8226),
            .I(N__8201));
    InMux I__1691 (
            .O(N__8225),
            .I(N__8193));
    InMux I__1690 (
            .O(N__8224),
            .I(N__8190));
    Span4Mux_v I__1689 (
            .O(N__8221),
            .I(N__8187));
    InMux I__1688 (
            .O(N__8220),
            .I(N__8184));
    InMux I__1687 (
            .O(N__8219),
            .I(N__8181));
    InMux I__1686 (
            .O(N__8216),
            .I(N__8176));
    InMux I__1685 (
            .O(N__8215),
            .I(N__8176));
    InMux I__1684 (
            .O(N__8214),
            .I(N__8169));
    InMux I__1683 (
            .O(N__8213),
            .I(N__8169));
    InMux I__1682 (
            .O(N__8212),
            .I(N__8169));
    Span4Mux_h I__1681 (
            .O(N__8209),
            .I(N__8162));
    LocalMux I__1680 (
            .O(N__8204),
            .I(N__8162));
    LocalMux I__1679 (
            .O(N__8201),
            .I(N__8162));
    InMux I__1678 (
            .O(N__8200),
            .I(N__8159));
    InMux I__1677 (
            .O(N__8199),
            .I(N__8154));
    InMux I__1676 (
            .O(N__8198),
            .I(N__8154));
    InMux I__1675 (
            .O(N__8197),
            .I(N__8149));
    InMux I__1674 (
            .O(N__8196),
            .I(N__8149));
    LocalMux I__1673 (
            .O(N__8193),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1672 (
            .O(N__8190),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1671 (
            .O(N__8187),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1670 (
            .O(N__8184),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1669 (
            .O(N__8181),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1668 (
            .O(N__8176),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1667 (
            .O(N__8169),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1666 (
            .O(N__8162),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1665 (
            .O(N__8159),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1664 (
            .O(N__8154),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1663 (
            .O(N__8149),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    CascadeMux I__1662 (
            .O(N__8126),
            .I(N__8122));
    CascadeMux I__1661 (
            .O(N__8125),
            .I(N__8118));
    InMux I__1660 (
            .O(N__8122),
            .I(N__8114));
    CascadeMux I__1659 (
            .O(N__8121),
            .I(N__8109));
    InMux I__1658 (
            .O(N__8118),
            .I(N__8103));
    InMux I__1657 (
            .O(N__8117),
            .I(N__8103));
    LocalMux I__1656 (
            .O(N__8114),
            .I(N__8100));
    InMux I__1655 (
            .O(N__8113),
            .I(N__8093));
    InMux I__1654 (
            .O(N__8112),
            .I(N__8093));
    InMux I__1653 (
            .O(N__8109),
            .I(N__8093));
    InMux I__1652 (
            .O(N__8108),
            .I(N__8084));
    LocalMux I__1651 (
            .O(N__8103),
            .I(N__8081));
    Span4Mux_v I__1650 (
            .O(N__8100),
            .I(N__8076));
    LocalMux I__1649 (
            .O(N__8093),
            .I(N__8076));
    InMux I__1648 (
            .O(N__8092),
            .I(N__8073));
    InMux I__1647 (
            .O(N__8091),
            .I(N__8070));
    InMux I__1646 (
            .O(N__8090),
            .I(N__8063));
    InMux I__1645 (
            .O(N__8089),
            .I(N__8063));
    InMux I__1644 (
            .O(N__8088),
            .I(N__8063));
    InMux I__1643 (
            .O(N__8087),
            .I(N__8060));
    LocalMux I__1642 (
            .O(N__8084),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1641 (
            .O(N__8081),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1640 (
            .O(N__8076),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1639 (
            .O(N__8073),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1638 (
            .O(N__8070),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1637 (
            .O(N__8063),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1636 (
            .O(N__8060),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    CascadeMux I__1635 (
            .O(N__8045),
            .I(N__8039));
    CascadeMux I__1634 (
            .O(N__8044),
            .I(N__8036));
    CascadeMux I__1633 (
            .O(N__8043),
            .I(N__8031));
    InMux I__1632 (
            .O(N__8042),
            .I(N__8022));
    InMux I__1631 (
            .O(N__8039),
            .I(N__8019));
    InMux I__1630 (
            .O(N__8036),
            .I(N__8016));
    CascadeMux I__1629 (
            .O(N__8035),
            .I(N__8012));
    InMux I__1628 (
            .O(N__8034),
            .I(N__8006));
    InMux I__1627 (
            .O(N__8031),
            .I(N__8001));
    InMux I__1626 (
            .O(N__8030),
            .I(N__8001));
    InMux I__1625 (
            .O(N__8029),
            .I(N__7998));
    InMux I__1624 (
            .O(N__8028),
            .I(N__7995));
    InMux I__1623 (
            .O(N__8027),
            .I(N__7988));
    InMux I__1622 (
            .O(N__8026),
            .I(N__7988));
    InMux I__1621 (
            .O(N__8025),
            .I(N__7988));
    LocalMux I__1620 (
            .O(N__8022),
            .I(N__7981));
    LocalMux I__1619 (
            .O(N__8019),
            .I(N__7981));
    LocalMux I__1618 (
            .O(N__8016),
            .I(N__7981));
    InMux I__1617 (
            .O(N__8015),
            .I(N__7978));
    InMux I__1616 (
            .O(N__8012),
            .I(N__7974));
    InMux I__1615 (
            .O(N__8011),
            .I(N__7970));
    CascadeMux I__1614 (
            .O(N__8010),
            .I(N__7965));
    InMux I__1613 (
            .O(N__8009),
            .I(N__7962));
    LocalMux I__1612 (
            .O(N__8006),
            .I(N__7959));
    LocalMux I__1611 (
            .O(N__8001),
            .I(N__7956));
    LocalMux I__1610 (
            .O(N__7998),
            .I(N__7945));
    LocalMux I__1609 (
            .O(N__7995),
            .I(N__7945));
    LocalMux I__1608 (
            .O(N__7988),
            .I(N__7945));
    Span4Mux_v I__1607 (
            .O(N__7981),
            .I(N__7945));
    LocalMux I__1606 (
            .O(N__7978),
            .I(N__7945));
    InMux I__1605 (
            .O(N__7977),
            .I(N__7939));
    LocalMux I__1604 (
            .O(N__7974),
            .I(N__7936));
    InMux I__1603 (
            .O(N__7973),
            .I(N__7933));
    LocalMux I__1602 (
            .O(N__7970),
            .I(N__7930));
    InMux I__1601 (
            .O(N__7969),
            .I(N__7927));
    InMux I__1600 (
            .O(N__7968),
            .I(N__7922));
    InMux I__1599 (
            .O(N__7965),
            .I(N__7922));
    LocalMux I__1598 (
            .O(N__7962),
            .I(N__7919));
    Span4Mux_v I__1597 (
            .O(N__7959),
            .I(N__7912));
    Span4Mux_h I__1596 (
            .O(N__7956),
            .I(N__7912));
    Span4Mux_v I__1595 (
            .O(N__7945),
            .I(N__7912));
    InMux I__1594 (
            .O(N__7944),
            .I(N__7905));
    InMux I__1593 (
            .O(N__7943),
            .I(N__7905));
    InMux I__1592 (
            .O(N__7942),
            .I(N__7905));
    LocalMux I__1591 (
            .O(N__7939),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1590 (
            .O(N__7936),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1589 (
            .O(N__7933),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1588 (
            .O(N__7930),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1587 (
            .O(N__7927),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1586 (
            .O(N__7922),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv12 I__1585 (
            .O(N__7919),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1584 (
            .O(N__7912),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1583 (
            .O(N__7905),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1582 (
            .O(N__7886),
            .I(N__7883));
    LocalMux I__1581 (
            .O(N__7883),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_29_i_a2_i_1_0 ));
    InMux I__1580 (
            .O(N__7880),
            .I(N__7873));
    InMux I__1579 (
            .O(N__7879),
            .I(N__7870));
    InMux I__1578 (
            .O(N__7878),
            .I(N__7863));
    InMux I__1577 (
            .O(N__7877),
            .I(N__7863));
    InMux I__1576 (
            .O(N__7876),
            .I(N__7863));
    LocalMux I__1575 (
            .O(N__7873),
            .I(N__7860));
    LocalMux I__1574 (
            .O(N__7870),
            .I(N__7855));
    LocalMux I__1573 (
            .O(N__7863),
            .I(N__7855));
    Span4Mux_v I__1572 (
            .O(N__7860),
            .I(N__7840));
    Span4Mux_h I__1571 (
            .O(N__7855),
            .I(N__7840));
    InMux I__1570 (
            .O(N__7854),
            .I(N__7837));
    InMux I__1569 (
            .O(N__7853),
            .I(N__7834));
    InMux I__1568 (
            .O(N__7852),
            .I(N__7829));
    InMux I__1567 (
            .O(N__7851),
            .I(N__7829));
    InMux I__1566 (
            .O(N__7850),
            .I(N__7826));
    InMux I__1565 (
            .O(N__7849),
            .I(N__7821));
    InMux I__1564 (
            .O(N__7848),
            .I(N__7821));
    InMux I__1563 (
            .O(N__7847),
            .I(N__7813));
    InMux I__1562 (
            .O(N__7846),
            .I(N__7813));
    InMux I__1561 (
            .O(N__7845),
            .I(N__7813));
    Span4Mux_h I__1560 (
            .O(N__7840),
            .I(N__7807));
    LocalMux I__1559 (
            .O(N__7837),
            .I(N__7807));
    LocalMux I__1558 (
            .O(N__7834),
            .I(N__7798));
    LocalMux I__1557 (
            .O(N__7829),
            .I(N__7798));
    LocalMux I__1556 (
            .O(N__7826),
            .I(N__7793));
    LocalMux I__1555 (
            .O(N__7821),
            .I(N__7793));
    CascadeMux I__1554 (
            .O(N__7820),
            .I(N__7787));
    LocalMux I__1553 (
            .O(N__7813),
            .I(N__7779));
    InMux I__1552 (
            .O(N__7812),
            .I(N__7776));
    Span4Mux_v I__1551 (
            .O(N__7807),
            .I(N__7773));
    InMux I__1550 (
            .O(N__7806),
            .I(N__7766));
    InMux I__1549 (
            .O(N__7805),
            .I(N__7766));
    InMux I__1548 (
            .O(N__7804),
            .I(N__7766));
    InMux I__1547 (
            .O(N__7803),
            .I(N__7763));
    Span4Mux_v I__1546 (
            .O(N__7798),
            .I(N__7756));
    Span4Mux_v I__1545 (
            .O(N__7793),
            .I(N__7756));
    InMux I__1544 (
            .O(N__7792),
            .I(N__7751));
    InMux I__1543 (
            .O(N__7791),
            .I(N__7751));
    InMux I__1542 (
            .O(N__7790),
            .I(N__7746));
    InMux I__1541 (
            .O(N__7787),
            .I(N__7746));
    InMux I__1540 (
            .O(N__7786),
            .I(N__7739));
    InMux I__1539 (
            .O(N__7785),
            .I(N__7739));
    InMux I__1538 (
            .O(N__7784),
            .I(N__7739));
    InMux I__1537 (
            .O(N__7783),
            .I(N__7734));
    InMux I__1536 (
            .O(N__7782),
            .I(N__7734));
    Span4Mux_v I__1535 (
            .O(N__7779),
            .I(N__7731));
    LocalMux I__1534 (
            .O(N__7776),
            .I(N__7722));
    Sp12to4 I__1533 (
            .O(N__7773),
            .I(N__7722));
    LocalMux I__1532 (
            .O(N__7766),
            .I(N__7722));
    LocalMux I__1531 (
            .O(N__7763),
            .I(N__7722));
    InMux I__1530 (
            .O(N__7762),
            .I(N__7717));
    InMux I__1529 (
            .O(N__7761),
            .I(N__7717));
    Sp12to4 I__1528 (
            .O(N__7756),
            .I(N__7706));
    LocalMux I__1527 (
            .O(N__7751),
            .I(N__7706));
    LocalMux I__1526 (
            .O(N__7746),
            .I(N__7706));
    LocalMux I__1525 (
            .O(N__7739),
            .I(N__7706));
    LocalMux I__1524 (
            .O(N__7734),
            .I(N__7706));
    Sp12to4 I__1523 (
            .O(N__7731),
            .I(N__7699));
    Span12Mux_v I__1522 (
            .O(N__7722),
            .I(N__7699));
    LocalMux I__1521 (
            .O(N__7717),
            .I(N__7699));
    Span12Mux_h I__1520 (
            .O(N__7706),
            .I(N__7696));
    Span12Mux_h I__1519 (
            .O(N__7699),
            .I(N__7693));
    Odrv12 I__1518 (
            .O(N__7696),
            .I(RESETn_c));
    Odrv12 I__1517 (
            .O(N__7693),
            .I(RESETn_c));
    IoInMux I__1516 (
            .O(N__7688),
            .I(N__7685));
    LocalMux I__1515 (
            .O(N__7685),
            .I(N__7682));
    Span12Mux_s9_v I__1514 (
            .O(N__7682),
            .I(N__7679));
    Odrv12 I__1513 (
            .O(N__7679),
            .I(RESETn_c_i));
    InMux I__1512 (
            .O(N__7676),
            .I(N__7673));
    LocalMux I__1511 (
            .O(N__7673),
            .I(N__7670));
    Span4Mux_h I__1510 (
            .O(N__7670),
            .I(N__7667));
    Sp12to4 I__1509 (
            .O(N__7667),
            .I(N__7664));
    Odrv12 I__1508 (
            .O(N__7664),
            .I(\U712_CHIP_RAM.un3_CPU_CYCLE_START ));
    CascadeMux I__1507 (
            .O(N__7661),
            .I(N__7658));
    InMux I__1506 (
            .O(N__7658),
            .I(N__7653));
    InMux I__1505 (
            .O(N__7657),
            .I(N__7650));
    InMux I__1504 (
            .O(N__7656),
            .I(N__7647));
    LocalMux I__1503 (
            .O(N__7653),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__1502 (
            .O(N__7650),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__1501 (
            .O(N__7647),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__1500 (
            .O(N__7640),
            .I(N__7637));
    InMux I__1499 (
            .O(N__7637),
            .I(N__7633));
    InMux I__1498 (
            .O(N__7636),
            .I(N__7630));
    LocalMux I__1497 (
            .O(N__7633),
            .I(N__7627));
    LocalMux I__1496 (
            .O(N__7630),
            .I(N__7624));
    Odrv4 I__1495 (
            .O(N__7627),
            .I(\U712_CHIP_RAM.N_177 ));
    Odrv4 I__1494 (
            .O(N__7624),
            .I(\U712_CHIP_RAM.N_177 ));
    InMux I__1493 (
            .O(N__7619),
            .I(N__7611));
    InMux I__1492 (
            .O(N__7618),
            .I(N__7608));
    InMux I__1491 (
            .O(N__7617),
            .I(N__7605));
    InMux I__1490 (
            .O(N__7616),
            .I(N__7602));
    InMux I__1489 (
            .O(N__7615),
            .I(N__7597));
    InMux I__1488 (
            .O(N__7614),
            .I(N__7597));
    LocalMux I__1487 (
            .O(N__7611),
            .I(N__7594));
    LocalMux I__1486 (
            .O(N__7608),
            .I(\U712_CHIP_RAM.N_172 ));
    LocalMux I__1485 (
            .O(N__7605),
            .I(\U712_CHIP_RAM.N_172 ));
    LocalMux I__1484 (
            .O(N__7602),
            .I(\U712_CHIP_RAM.N_172 ));
    LocalMux I__1483 (
            .O(N__7597),
            .I(\U712_CHIP_RAM.N_172 ));
    Odrv4 I__1482 (
            .O(N__7594),
            .I(\U712_CHIP_RAM.N_172 ));
    CascadeMux I__1481 (
            .O(N__7583),
            .I(N__7580));
    InMux I__1480 (
            .O(N__7580),
            .I(N__7576));
    InMux I__1479 (
            .O(N__7579),
            .I(N__7573));
    LocalMux I__1478 (
            .O(N__7576),
            .I(N__7570));
    LocalMux I__1477 (
            .O(N__7573),
            .I(\U712_CHIP_RAM.SDRAM_CMD_1_sqmuxa_1_0 ));
    Odrv12 I__1476 (
            .O(N__7570),
            .I(\U712_CHIP_RAM.SDRAM_CMD_1_sqmuxa_1_0 ));
    InMux I__1475 (
            .O(N__7565),
            .I(N__7561));
    InMux I__1474 (
            .O(N__7564),
            .I(N__7555));
    LocalMux I__1473 (
            .O(N__7561),
            .I(N__7551));
    InMux I__1472 (
            .O(N__7560),
            .I(N__7548));
    CascadeMux I__1471 (
            .O(N__7559),
            .I(N__7538));
    InMux I__1470 (
            .O(N__7558),
            .I(N__7534));
    LocalMux I__1469 (
            .O(N__7555),
            .I(N__7531));
    InMux I__1468 (
            .O(N__7554),
            .I(N__7528));
    Span4Mux_h I__1467 (
            .O(N__7551),
            .I(N__7525));
    LocalMux I__1466 (
            .O(N__7548),
            .I(N__7522));
    InMux I__1465 (
            .O(N__7547),
            .I(N__7517));
    InMux I__1464 (
            .O(N__7546),
            .I(N__7517));
    InMux I__1463 (
            .O(N__7545),
            .I(N__7508));
    InMux I__1462 (
            .O(N__7544),
            .I(N__7508));
    InMux I__1461 (
            .O(N__7543),
            .I(N__7508));
    InMux I__1460 (
            .O(N__7542),
            .I(N__7508));
    InMux I__1459 (
            .O(N__7541),
            .I(N__7505));
    InMux I__1458 (
            .O(N__7538),
            .I(N__7500));
    InMux I__1457 (
            .O(N__7537),
            .I(N__7500));
    LocalMux I__1456 (
            .O(N__7534),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1455 (
            .O(N__7531),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1454 (
            .O(N__7528),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1453 (
            .O(N__7525),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1452 (
            .O(N__7522),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1451 (
            .O(N__7517),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1450 (
            .O(N__7508),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1449 (
            .O(N__7505),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1448 (
            .O(N__7500),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1447 (
            .O(N__7481),
            .I(N__7475));
    InMux I__1446 (
            .O(N__7480),
            .I(N__7475));
    LocalMux I__1445 (
            .O(N__7475),
            .I(\U712_CHIP_RAM.N_186 ));
    CascadeMux I__1444 (
            .O(N__7472),
            .I(N__7469));
    InMux I__1443 (
            .O(N__7469),
            .I(N__7466));
    LocalMux I__1442 (
            .O(N__7466),
            .I(N__7463));
    Odrv4 I__1441 (
            .O(N__7463),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER34 ));
    CascadeMux I__1440 (
            .O(N__7460),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER34_cascade_ ));
    InMux I__1439 (
            .O(N__7457),
            .I(N__7454));
    LocalMux I__1438 (
            .O(N__7454),
            .I(N__7451));
    Span12Mux_v I__1437 (
            .O(N__7451),
            .I(N__7448));
    Span12Mux_h I__1436 (
            .O(N__7448),
            .I(N__7445));
    Odrv12 I__1435 (
            .O(N__7445),
            .I(A_c_2));
    IoInMux I__1434 (
            .O(N__7442),
            .I(N__7439));
    LocalMux I__1433 (
            .O(N__7439),
            .I(N__7435));
    InMux I__1432 (
            .O(N__7438),
            .I(N__7432));
    Span12Mux_s4_v I__1431 (
            .O(N__7435),
            .I(N__7427));
    LocalMux I__1430 (
            .O(N__7432),
            .I(N__7427));
    Span12Mux_v I__1429 (
            .O(N__7427),
            .I(N__7424));
    Span12Mux_h I__1428 (
            .O(N__7424),
            .I(N__7421));
    Odrv12 I__1427 (
            .O(N__7421),
            .I(A_c_9));
    InMux I__1426 (
            .O(N__7418),
            .I(N__7415));
    LocalMux I__1425 (
            .O(N__7415),
            .I(N__7412));
    Odrv12 I__1424 (
            .O(N__7412),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER16_2 ));
    InMux I__1423 (
            .O(N__7409),
            .I(N__7405));
    InMux I__1422 (
            .O(N__7408),
            .I(N__7402));
    LocalMux I__1421 (
            .O(N__7405),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER17_0 ));
    LocalMux I__1420 (
            .O(N__7402),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER17_0 ));
    CascadeMux I__1419 (
            .O(N__7397),
            .I(N__7391));
    InMux I__1418 (
            .O(N__7396),
            .I(N__7388));
    CascadeMux I__1417 (
            .O(N__7395),
            .I(N__7384));
    InMux I__1416 (
            .O(N__7394),
            .I(N__7381));
    InMux I__1415 (
            .O(N__7391),
            .I(N__7376));
    LocalMux I__1414 (
            .O(N__7388),
            .I(N__7371));
    InMux I__1413 (
            .O(N__7387),
            .I(N__7368));
    InMux I__1412 (
            .O(N__7384),
            .I(N__7365));
    LocalMux I__1411 (
            .O(N__7381),
            .I(N__7362));
    InMux I__1410 (
            .O(N__7380),
            .I(N__7359));
    InMux I__1409 (
            .O(N__7379),
            .I(N__7356));
    LocalMux I__1408 (
            .O(N__7376),
            .I(N__7353));
    InMux I__1407 (
            .O(N__7375),
            .I(N__7348));
    InMux I__1406 (
            .O(N__7374),
            .I(N__7348));
    Span4Mux_v I__1405 (
            .O(N__7371),
            .I(N__7343));
    LocalMux I__1404 (
            .O(N__7368),
            .I(N__7343));
    LocalMux I__1403 (
            .O(N__7365),
            .I(N__7334));
    Span4Mux_h I__1402 (
            .O(N__7362),
            .I(N__7334));
    LocalMux I__1401 (
            .O(N__7359),
            .I(N__7334));
    LocalMux I__1400 (
            .O(N__7356),
            .I(N__7334));
    Odrv12 I__1399 (
            .O(N__7353),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    LocalMux I__1398 (
            .O(N__7348),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__1397 (
            .O(N__7343),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    Odrv4 I__1396 (
            .O(N__7334),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15 ));
    CascadeMux I__1395 (
            .O(N__7325),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER17_0_cascade_ ));
    InMux I__1394 (
            .O(N__7322),
            .I(N__7318));
    InMux I__1393 (
            .O(N__7321),
            .I(N__7315));
    LocalMux I__1392 (
            .O(N__7318),
            .I(\U712_CHIP_RAM.N_33 ));
    LocalMux I__1391 (
            .O(N__7315),
            .I(\U712_CHIP_RAM.N_33 ));
    CascadeMux I__1390 (
            .O(N__7310),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER19_0_cascade_ ));
    CascadeMux I__1389 (
            .O(N__7307),
            .I(N__7304));
    InMux I__1388 (
            .O(N__7304),
            .I(N__7301));
    LocalMux I__1387 (
            .O(N__7301),
            .I(N__7296));
    InMux I__1386 (
            .O(N__7300),
            .I(N__7293));
    InMux I__1385 (
            .O(N__7299),
            .I(N__7290));
    Odrv12 I__1384 (
            .O(N__7296),
            .I(\U712_CHIP_RAM.CPU_CYCLE_DISABLEZ0 ));
    LocalMux I__1383 (
            .O(N__7293),
            .I(\U712_CHIP_RAM.CPU_CYCLE_DISABLEZ0 ));
    LocalMux I__1382 (
            .O(N__7290),
            .I(\U712_CHIP_RAM.CPU_CYCLE_DISABLEZ0 ));
    InMux I__1381 (
            .O(N__7283),
            .I(N__7280));
    LocalMux I__1380 (
            .O(N__7280),
            .I(N__7277));
    Span12Mux_h I__1379 (
            .O(N__7277),
            .I(N__7274));
    Odrv12 I__1378 (
            .O(N__7274),
            .I(\U712_CHIP_RAM.N_95 ));
    CascadeMux I__1377 (
            .O(N__7271),
            .I(N__7264));
    InMux I__1376 (
            .O(N__7270),
            .I(N__7261));
    InMux I__1375 (
            .O(N__7269),
            .I(N__7258));
    InMux I__1374 (
            .O(N__7268),
            .I(N__7252));
    InMux I__1373 (
            .O(N__7267),
            .I(N__7252));
    InMux I__1372 (
            .O(N__7264),
            .I(N__7249));
    LocalMux I__1371 (
            .O(N__7261),
            .I(N__7244));
    LocalMux I__1370 (
            .O(N__7258),
            .I(N__7241));
    InMux I__1369 (
            .O(N__7257),
            .I(N__7238));
    LocalMux I__1368 (
            .O(N__7252),
            .I(N__7233));
    LocalMux I__1367 (
            .O(N__7249),
            .I(N__7233));
    InMux I__1366 (
            .O(N__7248),
            .I(N__7230));
    InMux I__1365 (
            .O(N__7247),
            .I(N__7227));
    Span4Mux_v I__1364 (
            .O(N__7244),
            .I(N__7220));
    Span4Mux_v I__1363 (
            .O(N__7241),
            .I(N__7220));
    LocalMux I__1362 (
            .O(N__7238),
            .I(N__7220));
    Span4Mux_v I__1361 (
            .O(N__7233),
            .I(N__7217));
    LocalMux I__1360 (
            .O(N__7230),
            .I(\U712_CHIP_RAM.N_119 ));
    LocalMux I__1359 (
            .O(N__7227),
            .I(\U712_CHIP_RAM.N_119 ));
    Odrv4 I__1358 (
            .O(N__7220),
            .I(\U712_CHIP_RAM.N_119 ));
    Odrv4 I__1357 (
            .O(N__7217),
            .I(\U712_CHIP_RAM.N_119 ));
    InMux I__1356 (
            .O(N__7208),
            .I(N__7205));
    LocalMux I__1355 (
            .O(N__7205),
            .I(N__7201));
    InMux I__1354 (
            .O(N__7204),
            .I(N__7198));
    Span4Mux_h I__1353 (
            .O(N__7201),
            .I(N__7193));
    LocalMux I__1352 (
            .O(N__7198),
            .I(N__7190));
    InMux I__1351 (
            .O(N__7197),
            .I(N__7187));
    InMux I__1350 (
            .O(N__7196),
            .I(N__7184));
    Odrv4 I__1349 (
            .O(N__7193),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__1348 (
            .O(N__7190),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1347 (
            .O(N__7187),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1346 (
            .O(N__7184),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    CascadeMux I__1345 (
            .O(N__7175),
            .I(\U712_CHIP_RAM.N_95_cascade_ ));
    InMux I__1344 (
            .O(N__7172),
            .I(N__7169));
    LocalMux I__1343 (
            .O(N__7169),
            .I(N__7166));
    Span4Mux_h I__1342 (
            .O(N__7166),
            .I(N__7163));
    Odrv4 I__1341 (
            .O(N__7163),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_3_sqmuxa_1 ));
    CascadeMux I__1340 (
            .O(N__7160),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_3_sqmuxa_1_cascade_ ));
    CascadeMux I__1339 (
            .O(N__7157),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_cascade_ ));
    InMux I__1338 (
            .O(N__7154),
            .I(N__7151));
    LocalMux I__1337 (
            .O(N__7151),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_7 ));
    InMux I__1336 (
            .O(N__7148),
            .I(N__7142));
    InMux I__1335 (
            .O(N__7147),
            .I(N__7139));
    InMux I__1334 (
            .O(N__7146),
            .I(N__7136));
    InMux I__1333 (
            .O(N__7145),
            .I(N__7133));
    LocalMux I__1332 (
            .O(N__7142),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER38_1_0 ));
    LocalMux I__1331 (
            .O(N__7139),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER38_1_0 ));
    LocalMux I__1330 (
            .O(N__7136),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER38_1_0 ));
    LocalMux I__1329 (
            .O(N__7133),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER38_1_0 ));
    InMux I__1328 (
            .O(N__7124),
            .I(N__7121));
    LocalMux I__1327 (
            .O(N__7121),
            .I(N__7115));
    InMux I__1326 (
            .O(N__7120),
            .I(N__7110));
    InMux I__1325 (
            .O(N__7119),
            .I(N__7110));
    InMux I__1324 (
            .O(N__7118),
            .I(N__7107));
    Odrv4 I__1323 (
            .O(N__7115),
            .I(\U712_CHIP_RAM.N_94 ));
    LocalMux I__1322 (
            .O(N__7110),
            .I(\U712_CHIP_RAM.N_94 ));
    LocalMux I__1321 (
            .O(N__7107),
            .I(\U712_CHIP_RAM.N_94 ));
    CascadeMux I__1320 (
            .O(N__7100),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_cascade_ ));
    InMux I__1319 (
            .O(N__7097),
            .I(N__7094));
    LocalMux I__1318 (
            .O(N__7094),
            .I(\U712_CHIP_RAM.CPU_TACK_7_0 ));
    InMux I__1317 (
            .O(N__7091),
            .I(N__7085));
    InMux I__1316 (
            .O(N__7090),
            .I(N__7085));
    LocalMux I__1315 (
            .O(N__7085),
            .I(N__7081));
    InMux I__1314 (
            .O(N__7084),
            .I(N__7077));
    Span4Mux_h I__1313 (
            .O(N__7081),
            .I(N__7074));
    InMux I__1312 (
            .O(N__7080),
            .I(N__7071));
    LocalMux I__1311 (
            .O(N__7077),
            .I(CPU_TACKm));
    Odrv4 I__1310 (
            .O(N__7074),
            .I(CPU_TACKm));
    LocalMux I__1309 (
            .O(N__7071),
            .I(CPU_TACKm));
    InMux I__1308 (
            .O(N__7064),
            .I(N__7061));
    LocalMux I__1307 (
            .O(N__7061),
            .I(N__7058));
    Span12Mux_h I__1306 (
            .O(N__7058),
            .I(N__7055));
    Odrv12 I__1305 (
            .O(N__7055),
            .I(A_c_7));
    InMux I__1304 (
            .O(N__7052),
            .I(N__7049));
    LocalMux I__1303 (
            .O(N__7049),
            .I(N__7046));
    Span12Mux_h I__1302 (
            .O(N__7046),
            .I(N__7043));
    Span12Mux_v I__1301 (
            .O(N__7043),
            .I(N__7040));
    Odrv12 I__1300 (
            .O(N__7040),
            .I(A_c_14));
    InMux I__1299 (
            .O(N__7037),
            .I(N__7034));
    LocalMux I__1298 (
            .O(N__7034),
            .I(\U712_CHIP_RAM.N_173 ));
    IoInMux I__1297 (
            .O(N__7031),
            .I(N__7028));
    LocalMux I__1296 (
            .O(N__7028),
            .I(N__7025));
    Span4Mux_s2_v I__1295 (
            .O(N__7025),
            .I(N__7022));
    Span4Mux_h I__1294 (
            .O(N__7022),
            .I(N__7019));
    Span4Mux_v I__1293 (
            .O(N__7019),
            .I(N__7016));
    Odrv4 I__1292 (
            .O(N__7016),
            .I(N_56_i));
    InMux I__1291 (
            .O(N__7013),
            .I(N__7003));
    InMux I__1290 (
            .O(N__7012),
            .I(N__7003));
    InMux I__1289 (
            .O(N__7011),
            .I(N__6999));
    InMux I__1288 (
            .O(N__7010),
            .I(N__6992));
    InMux I__1287 (
            .O(N__7009),
            .I(N__6992));
    InMux I__1286 (
            .O(N__7008),
            .I(N__6992));
    LocalMux I__1285 (
            .O(N__7003),
            .I(N__6989));
    CascadeMux I__1284 (
            .O(N__7002),
            .I(N__6986));
    LocalMux I__1283 (
            .O(N__6999),
            .I(N__6983));
    LocalMux I__1282 (
            .O(N__6992),
            .I(N__6978));
    Span4Mux_v I__1281 (
            .O(N__6989),
            .I(N__6978));
    InMux I__1280 (
            .O(N__6986),
            .I(N__6975));
    Span4Mux_v I__1279 (
            .O(N__6983),
            .I(N__6972));
    Span4Mux_h I__1278 (
            .O(N__6978),
            .I(N__6966));
    LocalMux I__1277 (
            .O(N__6975),
            .I(N__6966));
    Span4Mux_v I__1276 (
            .O(N__6972),
            .I(N__6963));
    InMux I__1275 (
            .O(N__6971),
            .I(N__6960));
    Span4Mux_h I__1274 (
            .O(N__6966),
            .I(N__6957));
    Span4Mux_h I__1273 (
            .O(N__6963),
            .I(N__6954));
    LocalMux I__1272 (
            .O(N__6960),
            .I(N__6951));
    Sp12to4 I__1271 (
            .O(N__6957),
            .I(N__6948));
    Sp12to4 I__1270 (
            .O(N__6954),
            .I(N__6943));
    Span12Mux_v I__1269 (
            .O(N__6951),
            .I(N__6943));
    Span12Mux_v I__1268 (
            .O(N__6948),
            .I(N__6940));
    Odrv12 I__1267 (
            .O(N__6943),
            .I(SIZ_c_0));
    Odrv12 I__1266 (
            .O(N__6940),
            .I(SIZ_c_0));
    InMux I__1265 (
            .O(N__6935),
            .I(N__6923));
    InMux I__1264 (
            .O(N__6934),
            .I(N__6923));
    InMux I__1263 (
            .O(N__6933),
            .I(N__6923));
    InMux I__1262 (
            .O(N__6932),
            .I(N__6920));
    InMux I__1261 (
            .O(N__6931),
            .I(N__6915));
    InMux I__1260 (
            .O(N__6930),
            .I(N__6915));
    LocalMux I__1259 (
            .O(N__6923),
            .I(N__6908));
    LocalMux I__1258 (
            .O(N__6920),
            .I(N__6908));
    LocalMux I__1257 (
            .O(N__6915),
            .I(N__6908));
    Span4Mux_v I__1256 (
            .O(N__6908),
            .I(N__6905));
    Sp12to4 I__1255 (
            .O(N__6905),
            .I(N__6902));
    Span12Mux_h I__1254 (
            .O(N__6902),
            .I(N__6899));
    Odrv12 I__1253 (
            .O(N__6899),
            .I(A_c_1));
    CascadeMux I__1252 (
            .O(N__6896),
            .I(N__6891));
    CascadeMux I__1251 (
            .O(N__6895),
            .I(N__6888));
    CascadeMux I__1250 (
            .O(N__6894),
            .I(N__6885));
    InMux I__1249 (
            .O(N__6891),
            .I(N__6880));
    InMux I__1248 (
            .O(N__6888),
            .I(N__6880));
    InMux I__1247 (
            .O(N__6885),
            .I(N__6877));
    LocalMux I__1246 (
            .O(N__6880),
            .I(N__6870));
    LocalMux I__1245 (
            .O(N__6877),
            .I(N__6870));
    CascadeMux I__1244 (
            .O(N__6876),
            .I(N__6867));
    CascadeMux I__1243 (
            .O(N__6875),
            .I(N__6864));
    Span4Mux_v I__1242 (
            .O(N__6870),
            .I(N__6859));
    InMux I__1241 (
            .O(N__6867),
            .I(N__6852));
    InMux I__1240 (
            .O(N__6864),
            .I(N__6852));
    InMux I__1239 (
            .O(N__6863),
            .I(N__6852));
    InMux I__1238 (
            .O(N__6862),
            .I(N__6849));
    Span4Mux_h I__1237 (
            .O(N__6859),
            .I(N__6845));
    LocalMux I__1236 (
            .O(N__6852),
            .I(N__6842));
    LocalMux I__1235 (
            .O(N__6849),
            .I(N__6839));
    InMux I__1234 (
            .O(N__6848),
            .I(N__6836));
    Sp12to4 I__1233 (
            .O(N__6845),
            .I(N__6827));
    Span12Mux_h I__1232 (
            .O(N__6842),
            .I(N__6827));
    Sp12to4 I__1231 (
            .O(N__6839),
            .I(N__6827));
    LocalMux I__1230 (
            .O(N__6836),
            .I(N__6827));
    Odrv12 I__1229 (
            .O(N__6827),
            .I(A_c_0));
    CascadeMux I__1228 (
            .O(N__6824),
            .I(N__6819));
    InMux I__1227 (
            .O(N__6823),
            .I(N__6808));
    InMux I__1226 (
            .O(N__6822),
            .I(N__6808));
    InMux I__1225 (
            .O(N__6819),
            .I(N__6808));
    CascadeMux I__1224 (
            .O(N__6818),
            .I(N__6805));
    InMux I__1223 (
            .O(N__6817),
            .I(N__6802));
    InMux I__1222 (
            .O(N__6816),
            .I(N__6797));
    InMux I__1221 (
            .O(N__6815),
            .I(N__6797));
    LocalMux I__1220 (
            .O(N__6808),
            .I(N__6794));
    InMux I__1219 (
            .O(N__6805),
            .I(N__6791));
    LocalMux I__1218 (
            .O(N__6802),
            .I(N__6786));
    LocalMux I__1217 (
            .O(N__6797),
            .I(N__6786));
    Span4Mux_h I__1216 (
            .O(N__6794),
            .I(N__6781));
    LocalMux I__1215 (
            .O(N__6791),
            .I(N__6781));
    Span4Mux_v I__1214 (
            .O(N__6786),
            .I(N__6778));
    Span4Mux_h I__1213 (
            .O(N__6781),
            .I(N__6775));
    Span4Mux_v I__1212 (
            .O(N__6778),
            .I(N__6771));
    Span4Mux_v I__1211 (
            .O(N__6775),
            .I(N__6768));
    InMux I__1210 (
            .O(N__6774),
            .I(N__6765));
    Span4Mux_h I__1209 (
            .O(N__6771),
            .I(N__6762));
    Span4Mux_v I__1208 (
            .O(N__6768),
            .I(N__6759));
    LocalMux I__1207 (
            .O(N__6765),
            .I(N__6756));
    Sp12to4 I__1206 (
            .O(N__6762),
            .I(N__6749));
    Sp12to4 I__1205 (
            .O(N__6759),
            .I(N__6749));
    Span12Mux_v I__1204 (
            .O(N__6756),
            .I(N__6749));
    Odrv12 I__1203 (
            .O(N__6749),
            .I(SIZ_c_1));
    IoInMux I__1202 (
            .O(N__6746),
            .I(N__6743));
    LocalMux I__1201 (
            .O(N__6743),
            .I(N__6740));
    Span4Mux_s1_v I__1200 (
            .O(N__6740),
            .I(N__6737));
    Span4Mux_h I__1199 (
            .O(N__6737),
            .I(N__6734));
    Span4Mux_v I__1198 (
            .O(N__6734),
            .I(N__6731));
    Odrv4 I__1197 (
            .O(N__6731),
            .I(N_58_i));
    IoInMux I__1196 (
            .O(N__6728),
            .I(N__6725));
    LocalMux I__1195 (
            .O(N__6725),
            .I(N__6722));
    IoSpan4Mux I__1194 (
            .O(N__6722),
            .I(N__6719));
    IoSpan4Mux I__1193 (
            .O(N__6719),
            .I(N__6716));
    Span4Mux_s3_v I__1192 (
            .O(N__6716),
            .I(N__6713));
    Odrv4 I__1191 (
            .O(N__6713),
            .I(DMA_LATCH_EN_c));
    CEMux I__1190 (
            .O(N__6710),
            .I(N__6707));
    LocalMux I__1189 (
            .O(N__6707),
            .I(N__6704));
    Odrv4 I__1188 (
            .O(N__6704),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0_0 ));
    InMux I__1187 (
            .O(N__6701),
            .I(N__6698));
    LocalMux I__1186 (
            .O(N__6698),
            .I(N__6695));
    Span4Mux_v I__1185 (
            .O(N__6695),
            .I(N__6692));
    Sp12to4 I__1184 (
            .O(N__6692),
            .I(N__6689));
    Span12Mux_h I__1183 (
            .O(N__6689),
            .I(N__6686));
    Odrv12 I__1182 (
            .O(N__6686),
            .I(A_c_8));
    InMux I__1181 (
            .O(N__6683),
            .I(N__6680));
    LocalMux I__1180 (
            .O(N__6680),
            .I(N__6677));
    Span12Mux_v I__1179 (
            .O(N__6677),
            .I(N__6674));
    Span12Mux_h I__1178 (
            .O(N__6674),
            .I(N__6671));
    Odrv12 I__1177 (
            .O(N__6671),
            .I(A_c_15));
    InMux I__1176 (
            .O(N__6668),
            .I(N__6665));
    LocalMux I__1175 (
            .O(N__6665),
            .I(N__6662));
    Span4Mux_v I__1174 (
            .O(N__6662),
            .I(N__6659));
    Sp12to4 I__1173 (
            .O(N__6659),
            .I(N__6656));
    Span12Mux_h I__1172 (
            .O(N__6656),
            .I(N__6653));
    Span12Mux_v I__1171 (
            .O(N__6653),
            .I(N__6650));
    Odrv12 I__1170 (
            .O(N__6650),
            .I(A_c_16));
    InMux I__1169 (
            .O(N__6647),
            .I(N__6644));
    LocalMux I__1168 (
            .O(N__6644),
            .I(N__6641));
    Span12Mux_h I__1167 (
            .O(N__6641),
            .I(N__6638));
    Span12Mux_v I__1166 (
            .O(N__6638),
            .I(N__6635));
    Odrv12 I__1165 (
            .O(N__6635),
            .I(A_c_18));
    InMux I__1164 (
            .O(N__6632),
            .I(N__6629));
    LocalMux I__1163 (
            .O(N__6629),
            .I(N__6626));
    Span12Mux_v I__1162 (
            .O(N__6626),
            .I(N__6623));
    Span12Mux_h I__1161 (
            .O(N__6623),
            .I(N__6620));
    Odrv12 I__1160 (
            .O(N__6620),
            .I(A_c_13));
    InMux I__1159 (
            .O(N__6617),
            .I(N__6614));
    LocalMux I__1158 (
            .O(N__6614),
            .I(N__6611));
    Span4Mux_v I__1157 (
            .O(N__6611),
            .I(N__6608));
    Sp12to4 I__1156 (
            .O(N__6608),
            .I(N__6605));
    Span12Mux_h I__1155 (
            .O(N__6605),
            .I(N__6602));
    Odrv12 I__1154 (
            .O(N__6602),
            .I(A_c_6));
    InMux I__1153 (
            .O(N__6599),
            .I(N__6595));
    InMux I__1152 (
            .O(N__6598),
            .I(N__6592));
    LocalMux I__1151 (
            .O(N__6595),
            .I(\U712_CHIP_RAM.CLK_EN_5_0 ));
    LocalMux I__1150 (
            .O(N__6592),
            .I(\U712_CHIP_RAM.CLK_EN_5_0 ));
    CascadeMux I__1149 (
            .O(N__6587),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1_cascade_ ));
    InMux I__1148 (
            .O(N__6584),
            .I(N__6577));
    InMux I__1147 (
            .O(N__6583),
            .I(N__6577));
    InMux I__1146 (
            .O(N__6582),
            .I(N__6574));
    LocalMux I__1145 (
            .O(N__6577),
            .I(N__6571));
    LocalMux I__1144 (
            .O(N__6574),
            .I(\U712_CHIP_RAM.N_187 ));
    Odrv4 I__1143 (
            .O(N__6571),
            .I(\U712_CHIP_RAM.N_187 ));
    InMux I__1142 (
            .O(N__6566),
            .I(N__6563));
    LocalMux I__1141 (
            .O(N__6563),
            .I(N__6560));
    Odrv12 I__1140 (
            .O(N__6560),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0 ));
    InMux I__1139 (
            .O(N__6557),
            .I(N__6553));
    InMux I__1138 (
            .O(N__6556),
            .I(N__6550));
    LocalMux I__1137 (
            .O(N__6553),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0 ));
    LocalMux I__1136 (
            .O(N__6550),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0 ));
    CascadeMux I__1135 (
            .O(N__6545),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1_1_cascade_ ));
    InMux I__1134 (
            .O(N__6542),
            .I(N__6539));
    LocalMux I__1133 (
            .O(N__6539),
            .I(\U712_CHIP_RAM.N_155 ));
    CascadeMux I__1132 (
            .O(N__6536),
            .I(N__6533));
    InMux I__1131 (
            .O(N__6533),
            .I(N__6530));
    LocalMux I__1130 (
            .O(N__6530),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1 ));
    CascadeMux I__1129 (
            .O(N__6527),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ));
    InMux I__1128 (
            .O(N__6524),
            .I(N__6521));
    LocalMux I__1127 (
            .O(N__6521),
            .I(N__6518));
    Odrv12 I__1126 (
            .O(N__6518),
            .I(\U712_BYTE_ENABLE.N_58 ));
    CascadeMux I__1125 (
            .O(N__6515),
            .I(N__6512));
    InMux I__1124 (
            .O(N__6512),
            .I(N__6509));
    LocalMux I__1123 (
            .O(N__6509),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_7_2 ));
    CascadeMux I__1122 (
            .O(N__6506),
            .I(\U712_CHIP_RAM.BANK0_7_0_cascade_ ));
    IoInMux I__1121 (
            .O(N__6503),
            .I(N__6500));
    LocalMux I__1120 (
            .O(N__6500),
            .I(N__6497));
    IoSpan4Mux I__1119 (
            .O(N__6497),
            .I(N__6494));
    Sp12to4 I__1118 (
            .O(N__6494),
            .I(N__6491));
    Span12Mux_s7_v I__1117 (
            .O(N__6491),
            .I(N__6487));
    InMux I__1116 (
            .O(N__6490),
            .I(N__6484));
    Odrv12 I__1115 (
            .O(N__6487),
            .I(BANK0_c));
    LocalMux I__1114 (
            .O(N__6484),
            .I(BANK0_c));
    InMux I__1113 (
            .O(N__6479),
            .I(N__6476));
    LocalMux I__1112 (
            .O(N__6476),
            .I(N__6473));
    Span4Mux_v I__1111 (
            .O(N__6473),
            .I(N__6470));
    Sp12to4 I__1110 (
            .O(N__6470),
            .I(N__6467));
    Span12Mux_h I__1109 (
            .O(N__6467),
            .I(N__6464));
    Odrv12 I__1108 (
            .O(N__6464),
            .I(A_c_20));
    InMux I__1107 (
            .O(N__6461),
            .I(N__6458));
    LocalMux I__1106 (
            .O(N__6458),
            .I(\U712_CHIP_RAM.A_m_20 ));
    CascadeMux I__1105 (
            .O(N__6455),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ));
    InMux I__1104 (
            .O(N__6452),
            .I(N__6449));
    LocalMux I__1103 (
            .O(N__6449),
            .I(N__6445));
    InMux I__1102 (
            .O(N__6448),
            .I(N__6442));
    Odrv12 I__1101 (
            .O(N__6445),
            .I(\U712_CHIP_RAM.A_m_2_20 ));
    LocalMux I__1100 (
            .O(N__6442),
            .I(\U712_CHIP_RAM.A_m_2_20 ));
    CascadeMux I__1099 (
            .O(N__6437),
            .I(\U712_CHIP_RAM.N_94_cascade_ ));
    CascadeMux I__1098 (
            .O(N__6434),
            .I(\U712_CHIP_RAM.N_108_cascade_ ));
    CascadeMux I__1097 (
            .O(N__6431),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_a3_0_cascade_ ));
    InMux I__1096 (
            .O(N__6428),
            .I(N__6425));
    LocalMux I__1095 (
            .O(N__6425),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_0 ));
    CascadeMux I__1094 (
            .O(N__6422),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_0_cascade_ ));
    IoInMux I__1093 (
            .O(N__6419),
            .I(N__6416));
    LocalMux I__1092 (
            .O(N__6416),
            .I(N__6413));
    Span12Mux_s10_h I__1091 (
            .O(N__6413),
            .I(N__6410));
    Span12Mux_v I__1090 (
            .O(N__6410),
            .I(N__6406));
    InMux I__1089 (
            .O(N__6409),
            .I(N__6403));
    Odrv12 I__1088 (
            .O(N__6406),
            .I(CLK_EN_c));
    LocalMux I__1087 (
            .O(N__6403),
            .I(CLK_EN_c));
    InMux I__1086 (
            .O(N__6398),
            .I(N__6395));
    LocalMux I__1085 (
            .O(N__6395),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_0_0 ));
    InMux I__1084 (
            .O(N__6392),
            .I(N__6387));
    InMux I__1083 (
            .O(N__6391),
            .I(N__6384));
    InMux I__1082 (
            .O(N__6390),
            .I(N__6381));
    LocalMux I__1081 (
            .O(N__6387),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__1080 (
            .O(N__6384),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__1079 (
            .O(N__6381),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__1078 (
            .O(N__6374),
            .I(N__6369));
    InMux I__1077 (
            .O(N__6373),
            .I(N__6366));
    InMux I__1076 (
            .O(N__6372),
            .I(N__6363));
    LocalMux I__1075 (
            .O(N__6369),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__1074 (
            .O(N__6366),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__1073 (
            .O(N__6363),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__1072 (
            .O(N__6356),
            .I(N__6351));
    CascadeMux I__1071 (
            .O(N__6355),
            .I(N__6348));
    InMux I__1070 (
            .O(N__6354),
            .I(N__6345));
    InMux I__1069 (
            .O(N__6351),
            .I(N__6342));
    InMux I__1068 (
            .O(N__6348),
            .I(N__6339));
    LocalMux I__1067 (
            .O(N__6345),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1066 (
            .O(N__6342),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1065 (
            .O(N__6339),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__1064 (
            .O(N__6332),
            .I(N__6327));
    InMux I__1063 (
            .O(N__6331),
            .I(N__6324));
    InMux I__1062 (
            .O(N__6330),
            .I(N__6321));
    LocalMux I__1061 (
            .O(N__6327),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1060 (
            .O(N__6324),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1059 (
            .O(N__6321),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    CascadeMux I__1058 (
            .O(N__6314),
            .I(\U712_CHIP_RAM.N_331_3_cascade_ ));
    CascadeMux I__1057 (
            .O(N__6311),
            .I(N__6307));
    InMux I__1056 (
            .O(N__6310),
            .I(N__6301));
    InMux I__1055 (
            .O(N__6307),
            .I(N__6301));
    InMux I__1054 (
            .O(N__6306),
            .I(N__6298));
    LocalMux I__1053 (
            .O(N__6301),
            .I(N__6295));
    LocalMux I__1052 (
            .O(N__6298),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER37_0_a3_1_0 ));
    Odrv4 I__1051 (
            .O(N__6295),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER37_0_a3_1_0 ));
    CascadeMux I__1050 (
            .O(N__6290),
            .I(\U712_CHIP_RAM.LATCH_CLK_0_sqmuxa_cascade_ ));
    CascadeMux I__1049 (
            .O(N__6287),
            .I(N__6284));
    InMux I__1048 (
            .O(N__6284),
            .I(N__6277));
    InMux I__1047 (
            .O(N__6283),
            .I(N__6277));
    InMux I__1046 (
            .O(N__6282),
            .I(N__6274));
    LocalMux I__1045 (
            .O(N__6277),
            .I(N__6270));
    LocalMux I__1044 (
            .O(N__6274),
            .I(N__6267));
    InMux I__1043 (
            .O(N__6273),
            .I(N__6264));
    Span4Mux_v I__1042 (
            .O(N__6270),
            .I(N__6259));
    Span4Mux_h I__1041 (
            .O(N__6267),
            .I(N__6259));
    LocalMux I__1040 (
            .O(N__6264),
            .I(REG_TACK));
    Odrv4 I__1039 (
            .O(N__6259),
            .I(REG_TACK));
    InMux I__1038 (
            .O(N__6254),
            .I(N__6251));
    LocalMux I__1037 (
            .O(N__6251),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    InMux I__1036 (
            .O(N__6248),
            .I(N__6245));
    LocalMux I__1035 (
            .O(N__6245),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0 ));
    CascadeMux I__1034 (
            .O(N__6242),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0_cascade_ ));
    InMux I__1033 (
            .O(N__6239),
            .I(N__6236));
    LocalMux I__1032 (
            .O(N__6236),
            .I(N__6232));
    InMux I__1031 (
            .O(N__6235),
            .I(N__6229));
    Span4Mux_v I__1030 (
            .O(N__6232),
            .I(N__6226));
    LocalMux I__1029 (
            .O(N__6229),
            .I(N__6223));
    Span4Mux_h I__1028 (
            .O(N__6226),
            .I(N__6220));
    Span12Mux_h I__1027 (
            .O(N__6223),
            .I(N__6215));
    Sp12to4 I__1026 (
            .O(N__6220),
            .I(N__6215));
    Span12Mux_v I__1025 (
            .O(N__6215),
            .I(N__6212));
    Odrv12 I__1024 (
            .O(N__6212),
            .I(AWEn_c));
    InMux I__1023 (
            .O(N__6209),
            .I(N__6206));
    LocalMux I__1022 (
            .O(N__6206),
            .I(N__6202));
    InMux I__1021 (
            .O(N__6205),
            .I(N__6199));
    Span4Mux_h I__1020 (
            .O(N__6202),
            .I(N__6193));
    LocalMux I__1019 (
            .O(N__6199),
            .I(N__6190));
    InMux I__1018 (
            .O(N__6198),
            .I(N__6183));
    InMux I__1017 (
            .O(N__6197),
            .I(N__6183));
    InMux I__1016 (
            .O(N__6196),
            .I(N__6183));
    Span4Mux_h I__1015 (
            .O(N__6193),
            .I(N__6180));
    Span4Mux_v I__1014 (
            .O(N__6190),
            .I(N__6175));
    LocalMux I__1013 (
            .O(N__6183),
            .I(N__6175));
    Odrv4 I__1012 (
            .O(N__6180),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1011 (
            .O(N__6175),
            .I(DBR_SYNCZ0Z_1));
    InMux I__1010 (
            .O(N__6170),
            .I(N__6167));
    LocalMux I__1009 (
            .O(N__6167),
            .I(N__6164));
    Odrv4 I__1008 (
            .O(N__6164),
            .I(\U712_CHIP_RAM.N_152 ));
    CascadeMux I__1007 (
            .O(N__6161),
            .I(N__6158));
    InMux I__1006 (
            .O(N__6158),
            .I(N__6154));
    CascadeMux I__1005 (
            .O(N__6157),
            .I(N__6148));
    LocalMux I__1004 (
            .O(N__6154),
            .I(N__6145));
    InMux I__1003 (
            .O(N__6153),
            .I(N__6142));
    InMux I__1002 (
            .O(N__6152),
            .I(N__6139));
    InMux I__1001 (
            .O(N__6151),
            .I(N__6136));
    InMux I__1000 (
            .O(N__6148),
            .I(N__6133));
    Span4Mux_v I__999 (
            .O(N__6145),
            .I(N__6128));
    LocalMux I__998 (
            .O(N__6142),
            .I(N__6128));
    LocalMux I__997 (
            .O(N__6139),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__996 (
            .O(N__6136),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__995 (
            .O(N__6133),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    Odrv4 I__994 (
            .O(N__6128),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__993 (
            .O(N__6119),
            .I(N__6114));
    InMux I__992 (
            .O(N__6118),
            .I(N__6109));
    InMux I__991 (
            .O(N__6117),
            .I(N__6109));
    LocalMux I__990 (
            .O(N__6114),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__989 (
            .O(N__6109),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    CascadeMux I__988 (
            .O(N__6104),
            .I(N__6101));
    InMux I__987 (
            .O(N__6101),
            .I(N__6095));
    InMux I__986 (
            .O(N__6100),
            .I(N__6095));
    LocalMux I__985 (
            .O(N__6095),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    InMux I__984 (
            .O(N__6092),
            .I(N__6089));
    LocalMux I__983 (
            .O(N__6089),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0 ));
    InMux I__982 (
            .O(N__6086),
            .I(N__6082));
    InMux I__981 (
            .O(N__6085),
            .I(N__6079));
    LocalMux I__980 (
            .O(N__6082),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__979 (
            .O(N__6079),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__978 (
            .O(N__6074),
            .I(N__6069));
    InMux I__977 (
            .O(N__6073),
            .I(N__6066));
    InMux I__976 (
            .O(N__6072),
            .I(N__6062));
    InMux I__975 (
            .O(N__6069),
            .I(N__6059));
    LocalMux I__974 (
            .O(N__6066),
            .I(N__6056));
    InMux I__973 (
            .O(N__6065),
            .I(N__6053));
    LocalMux I__972 (
            .O(N__6062),
            .I(N__6048));
    LocalMux I__971 (
            .O(N__6059),
            .I(N__6048));
    Span4Mux_h I__970 (
            .O(N__6056),
            .I(N__6045));
    LocalMux I__969 (
            .O(N__6053),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    Odrv4 I__968 (
            .O(N__6048),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    Odrv4 I__967 (
            .O(N__6045),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__966 (
            .O(N__6038),
            .I(N__6029));
    InMux I__965 (
            .O(N__6037),
            .I(N__6029));
    InMux I__964 (
            .O(N__6036),
            .I(N__6029));
    LocalMux I__963 (
            .O(N__6029),
            .I(N__6026));
    Odrv4 I__962 (
            .O(N__6026),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    SRMux I__961 (
            .O(N__6023),
            .I(N__6020));
    LocalMux I__960 (
            .O(N__6020),
            .I(N__6017));
    Odrv4 I__959 (
            .O(N__6017),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    IoInMux I__958 (
            .O(N__6014),
            .I(N__6011));
    LocalMux I__957 (
            .O(N__6011),
            .I(N__6008));
    IoSpan4Mux I__956 (
            .O(N__6008),
            .I(N__6005));
    Span4Mux_s3_h I__955 (
            .O(N__6005),
            .I(N__6002));
    Sp12to4 I__954 (
            .O(N__6002),
            .I(N__5999));
    Span12Mux_h I__953 (
            .O(N__5999),
            .I(N__5996));
    Odrv12 I__952 (
            .O(N__5996),
            .I(CLMBEn_c));
    InMux I__951 (
            .O(N__5993),
            .I(N__5990));
    LocalMux I__950 (
            .O(N__5990),
            .I(N__5987));
    Span4Mux_h I__949 (
            .O(N__5987),
            .I(N__5984));
    Odrv4 I__948 (
            .O(N__5984),
            .I(\U712_CHIP_RAM.LATCH_CLK_0_sqmuxa ));
    InMux I__947 (
            .O(N__5981),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__946 (
            .O(N__5978),
            .I(N__5975));
    LocalMux I__945 (
            .O(N__5975),
            .I(N__5972));
    Odrv4 I__944 (
            .O(N__5972),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__943 (
            .O(N__5969),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__942 (
            .O(N__5966),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__941 (
            .O(N__5963),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__940 (
            .O(N__5960),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__939 (
            .O(N__5957),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__938 (
            .O(N__5954),
            .I(N__5941));
    InMux I__937 (
            .O(N__5953),
            .I(N__5941));
    InMux I__936 (
            .O(N__5952),
            .I(N__5941));
    InMux I__935 (
            .O(N__5951),
            .I(N__5938));
    InMux I__934 (
            .O(N__5950),
            .I(N__5931));
    InMux I__933 (
            .O(N__5949),
            .I(N__5931));
    InMux I__932 (
            .O(N__5948),
            .I(N__5931));
    LocalMux I__931 (
            .O(N__5941),
            .I(\U712_CHIP_RAM.N_64 ));
    LocalMux I__930 (
            .O(N__5938),
            .I(\U712_CHIP_RAM.N_64 ));
    LocalMux I__929 (
            .O(N__5931),
            .I(\U712_CHIP_RAM.N_64 ));
    InMux I__928 (
            .O(N__5924),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    CEMux I__927 (
            .O(N__5921),
            .I(N__5917));
    CEMux I__926 (
            .O(N__5920),
            .I(N__5914));
    LocalMux I__925 (
            .O(N__5917),
            .I(N__5911));
    LocalMux I__924 (
            .O(N__5914),
            .I(N__5908));
    Odrv4 I__923 (
            .O(N__5911),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv12 I__922 (
            .O(N__5908),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    CascadeMux I__921 (
            .O(N__5903),
            .I(N__5898));
    InMux I__920 (
            .O(N__5902),
            .I(N__5895));
    InMux I__919 (
            .O(N__5901),
            .I(N__5892));
    InMux I__918 (
            .O(N__5898),
            .I(N__5889));
    LocalMux I__917 (
            .O(N__5895),
            .I(N__5885));
    LocalMux I__916 (
            .O(N__5892),
            .I(N__5880));
    LocalMux I__915 (
            .O(N__5889),
            .I(N__5880));
    InMux I__914 (
            .O(N__5888),
            .I(N__5877));
    Span4Mux_v I__913 (
            .O(N__5885),
            .I(N__5874));
    Span4Mux_v I__912 (
            .O(N__5880),
            .I(N__5871));
    LocalMux I__911 (
            .O(N__5877),
            .I(N__5868));
    Span4Mux_v I__910 (
            .O(N__5874),
            .I(N__5865));
    Span4Mux_v I__909 (
            .O(N__5871),
            .I(N__5862));
    Span4Mux_h I__908 (
            .O(N__5868),
            .I(N__5859));
    Sp12to4 I__907 (
            .O(N__5865),
            .I(N__5856));
    Sp12to4 I__906 (
            .O(N__5862),
            .I(N__5853));
    Sp12to4 I__905 (
            .O(N__5859),
            .I(N__5850));
    Span12Mux_h I__904 (
            .O(N__5856),
            .I(N__5843));
    Span12Mux_h I__903 (
            .O(N__5853),
            .I(N__5843));
    Span12Mux_v I__902 (
            .O(N__5850),
            .I(N__5843));
    Odrv12 I__901 (
            .O(N__5843),
            .I(CLK40_PLL_i));
    CascadeMux I__900 (
            .O(N__5840),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER33_1_0_cascade_ ));
    CascadeMux I__899 (
            .O(N__5837),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_2_cascade_ ));
    CascadeMux I__898 (
            .O(N__5834),
            .I(\U712_CHIP_RAM.N_64_cascade_ ));
    IoInMux I__897 (
            .O(N__5831),
            .I(N__5828));
    LocalMux I__896 (
            .O(N__5828),
            .I(N__5824));
    InMux I__895 (
            .O(N__5827),
            .I(N__5821));
    Span12Mux_s7_v I__894 (
            .O(N__5824),
            .I(N__5818));
    LocalMux I__893 (
            .O(N__5821),
            .I(N__5815));
    Odrv12 I__892 (
            .O(N__5818),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__891 (
            .O(N__5815),
            .I(CONSTANT_ONE_NET));
    InMux I__890 (
            .O(N__5810),
            .I(N__5807));
    LocalMux I__889 (
            .O(N__5807),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0 ));
    InMux I__888 (
            .O(N__5804),
            .I(N__5799));
    InMux I__887 (
            .O(N__5803),
            .I(N__5794));
    InMux I__886 (
            .O(N__5802),
            .I(N__5794));
    LocalMux I__885 (
            .O(N__5799),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER18 ));
    LocalMux I__884 (
            .O(N__5794),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER18 ));
    InMux I__883 (
            .O(N__5789),
            .I(N__5786));
    LocalMux I__882 (
            .O(N__5786),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_1 ));
    InMux I__881 (
            .O(N__5783),
            .I(N__5780));
    LocalMux I__880 (
            .O(N__5780),
            .I(\U712_CHIP_RAM.LATCH_CLK_6 ));
    InMux I__879 (
            .O(N__5777),
            .I(N__5773));
    InMux I__878 (
            .O(N__5776),
            .I(N__5770));
    LocalMux I__877 (
            .O(N__5773),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__876 (
            .O(N__5770),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__875 (
            .O(N__5765),
            .I(N__5761));
    InMux I__874 (
            .O(N__5764),
            .I(N__5758));
    LocalMux I__873 (
            .O(N__5761),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__872 (
            .O(N__5758),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__871 (
            .O(N__5753),
            .I(N__5749));
    InMux I__870 (
            .O(N__5752),
            .I(N__5746));
    LocalMux I__869 (
            .O(N__5749),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__868 (
            .O(N__5746),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__867 (
            .O(N__5741),
            .I(N__5737));
    InMux I__866 (
            .O(N__5740),
            .I(N__5734));
    LocalMux I__865 (
            .O(N__5737),
            .I(\U712_CHIP_RAM.N_9 ));
    LocalMux I__864 (
            .O(N__5734),
            .I(\U712_CHIP_RAM.N_9 ));
    InMux I__863 (
            .O(N__5729),
            .I(N__5723));
    InMux I__862 (
            .O(N__5728),
            .I(N__5720));
    InMux I__861 (
            .O(N__5727),
            .I(N__5717));
    InMux I__860 (
            .O(N__5726),
            .I(N__5714));
    LocalMux I__859 (
            .O(N__5723),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__858 (
            .O(N__5720),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__857 (
            .O(N__5717),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__856 (
            .O(N__5714),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__855 (
            .O(N__5705),
            .I(N__5701));
    InMux I__854 (
            .O(N__5704),
            .I(N__5698));
    LocalMux I__853 (
            .O(N__5701),
            .I(N__5695));
    LocalMux I__852 (
            .O(N__5698),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    Odrv4 I__851 (
            .O(N__5695),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__850 (
            .O(N__5690),
            .I(N__5687));
    LocalMux I__849 (
            .O(N__5687),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ));
    InMux I__848 (
            .O(N__5684),
            .I(N__5681));
    LocalMux I__847 (
            .O(N__5681),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    CascadeMux I__846 (
            .O(N__5678),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER18_cascade_ ));
    CascadeMux I__845 (
            .O(N__5675),
            .I(N__5672));
    InMux I__844 (
            .O(N__5672),
            .I(N__5666));
    InMux I__843 (
            .O(N__5671),
            .I(N__5661));
    InMux I__842 (
            .O(N__5670),
            .I(N__5661));
    InMux I__841 (
            .O(N__5669),
            .I(N__5658));
    LocalMux I__840 (
            .O(N__5666),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__839 (
            .O(N__5661),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__838 (
            .O(N__5658),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__837 (
            .O(N__5651),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__836 (
            .O(N__5648),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__835 (
            .O(N__5645),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__834 (
            .O(N__5642),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__833 (
            .O(N__5639),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__832 (
            .O(N__5636),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__831 (
            .O(N__5633),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__830 (
            .O(N__5630),
            .I(N__5603));
    ClkMux I__829 (
            .O(N__5629),
            .I(N__5603));
    ClkMux I__828 (
            .O(N__5628),
            .I(N__5603));
    ClkMux I__827 (
            .O(N__5627),
            .I(N__5603));
    ClkMux I__826 (
            .O(N__5626),
            .I(N__5603));
    ClkMux I__825 (
            .O(N__5625),
            .I(N__5603));
    ClkMux I__824 (
            .O(N__5624),
            .I(N__5603));
    ClkMux I__823 (
            .O(N__5623),
            .I(N__5603));
    ClkMux I__822 (
            .O(N__5622),
            .I(N__5603));
    GlobalMux I__821 (
            .O(N__5603),
            .I(N__5600));
    gio2CtrlBuf I__820 (
            .O(N__5600),
            .I(C1_c_g));
    InMux I__819 (
            .O(N__5597),
            .I(N__5593));
    InMux I__818 (
            .O(N__5596),
            .I(N__5590));
    LocalMux I__817 (
            .O(N__5593),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__816 (
            .O(N__5590),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    InMux I__815 (
            .O(N__5585),
            .I(N__5581));
    InMux I__814 (
            .O(N__5584),
            .I(N__5578));
    LocalMux I__813 (
            .O(N__5581),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    LocalMux I__812 (
            .O(N__5578),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    CascadeMux I__811 (
            .O(N__5573),
            .I(N__5569));
    InMux I__810 (
            .O(N__5572),
            .I(N__5566));
    InMux I__809 (
            .O(N__5569),
            .I(N__5563));
    LocalMux I__808 (
            .O(N__5566),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__807 (
            .O(N__5563),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__806 (
            .O(N__5558),
            .I(N__5554));
    InMux I__805 (
            .O(N__5557),
            .I(N__5551));
    LocalMux I__804 (
            .O(N__5554),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    LocalMux I__803 (
            .O(N__5551),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__802 (
            .O(N__5546),
            .I(N__5543));
    LocalMux I__801 (
            .O(N__5543),
            .I(\U712_CHIP_RAM.DMA_CYCLE_START_2_0 ));
    InMux I__800 (
            .O(N__5540),
            .I(N__5537));
    LocalMux I__799 (
            .O(N__5537),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_3 ));
    CascadeMux I__798 (
            .O(N__5534),
            .I(N__5527));
    CascadeMux I__797 (
            .O(N__5533),
            .I(N__5518));
    InMux I__796 (
            .O(N__5532),
            .I(N__5514));
    InMux I__795 (
            .O(N__5531),
            .I(N__5509));
    InMux I__794 (
            .O(N__5530),
            .I(N__5506));
    InMux I__793 (
            .O(N__5527),
            .I(N__5501));
    InMux I__792 (
            .O(N__5526),
            .I(N__5501));
    InMux I__791 (
            .O(N__5525),
            .I(N__5496));
    InMux I__790 (
            .O(N__5524),
            .I(N__5496));
    InMux I__789 (
            .O(N__5523),
            .I(N__5489));
    InMux I__788 (
            .O(N__5522),
            .I(N__5489));
    InMux I__787 (
            .O(N__5521),
            .I(N__5489));
    InMux I__786 (
            .O(N__5518),
            .I(N__5485));
    InMux I__785 (
            .O(N__5517),
            .I(N__5482));
    LocalMux I__784 (
            .O(N__5514),
            .I(N__5479));
    InMux I__783 (
            .O(N__5513),
            .I(N__5474));
    InMux I__782 (
            .O(N__5512),
            .I(N__5474));
    LocalMux I__781 (
            .O(N__5509),
            .I(N__5471));
    LocalMux I__780 (
            .O(N__5506),
            .I(N__5466));
    LocalMux I__779 (
            .O(N__5501),
            .I(N__5466));
    LocalMux I__778 (
            .O(N__5496),
            .I(N__5461));
    LocalMux I__777 (
            .O(N__5489),
            .I(N__5461));
    InMux I__776 (
            .O(N__5488),
            .I(N__5458));
    LocalMux I__775 (
            .O(N__5485),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__774 (
            .O(N__5482),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__773 (
            .O(N__5479),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__772 (
            .O(N__5474),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__771 (
            .O(N__5471),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv12 I__770 (
            .O(N__5466),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__769 (
            .O(N__5461),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__768 (
            .O(N__5458),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    IoInMux I__767 (
            .O(N__5441),
            .I(N__5438));
    LocalMux I__766 (
            .O(N__5438),
            .I(N__5435));
    Span4Mux_s2_v I__765 (
            .O(N__5435),
            .I(N__5432));
    Span4Mux_h I__764 (
            .O(N__5432),
            .I(N__5429));
    Span4Mux_h I__763 (
            .O(N__5429),
            .I(N__5426));
    Sp12to4 I__762 (
            .O(N__5426),
            .I(N__5423));
    Span12Mux_s10_v I__761 (
            .O(N__5423),
            .I(N__5420));
    Odrv12 I__760 (
            .O(N__5420),
            .I(ASn_c));
    CEMux I__759 (
            .O(N__5417),
            .I(N__5414));
    LocalMux I__758 (
            .O(N__5414),
            .I(N__5411));
    Span4Mux_v I__757 (
            .O(N__5411),
            .I(N__5408));
    Odrv4 I__756 (
            .O(N__5408),
            .I(\U712_REG_SM.N_163_0 ));
    InMux I__755 (
            .O(N__5405),
            .I(N__5402));
    LocalMux I__754 (
            .O(N__5402),
            .I(N__5398));
    InMux I__753 (
            .O(N__5401),
            .I(N__5395));
    Span4Mux_v I__752 (
            .O(N__5398),
            .I(N__5392));
    LocalMux I__751 (
            .O(N__5395),
            .I(N__5389));
    Span4Mux_v I__750 (
            .O(N__5392),
            .I(N__5384));
    Span4Mux_h I__749 (
            .O(N__5389),
            .I(N__5384));
    Span4Mux_v I__748 (
            .O(N__5384),
            .I(N__5381));
    IoSpan4Mux I__747 (
            .O(N__5381),
            .I(N__5378));
    Odrv4 I__746 (
            .O(N__5378),
            .I(TSn_c));
    InMux I__745 (
            .O(N__5375),
            .I(N__5372));
    LocalMux I__744 (
            .O(N__5372),
            .I(N__5368));
    IoInMux I__743 (
            .O(N__5371),
            .I(N__5365));
    Span4Mux_h I__742 (
            .O(N__5368),
            .I(N__5362));
    LocalMux I__741 (
            .O(N__5365),
            .I(N__5359));
    Span4Mux_v I__740 (
            .O(N__5362),
            .I(N__5356));
    IoSpan4Mux I__739 (
            .O(N__5359),
            .I(N__5353));
    Odrv4 I__738 (
            .O(N__5356),
            .I(RAMENn_c));
    Odrv4 I__737 (
            .O(N__5353),
            .I(RAMENn_c));
    IoInMux I__736 (
            .O(N__5348),
            .I(N__5345));
    LocalMux I__735 (
            .O(N__5345),
            .I(N__5342));
    Span4Mux_s3_v I__734 (
            .O(N__5342),
            .I(N__5339));
    Span4Mux_v I__733 (
            .O(N__5339),
            .I(N__5336));
    Span4Mux_v I__732 (
            .O(N__5336),
            .I(N__5333));
    Odrv4 I__731 (
            .O(N__5333),
            .I(VBENn_c));
    InMux I__730 (
            .O(N__5330),
            .I(N__5327));
    LocalMux I__729 (
            .O(N__5327),
            .I(\U712_CYCLE_TERM.N_47_0 ));
    IoInMux I__728 (
            .O(N__5324),
            .I(N__5320));
    IoInMux I__727 (
            .O(N__5323),
            .I(N__5316));
    LocalMux I__726 (
            .O(N__5320),
            .I(N__5313));
    IoInMux I__725 (
            .O(N__5319),
            .I(N__5310));
    LocalMux I__724 (
            .O(N__5316),
            .I(N__5307));
    IoSpan4Mux I__723 (
            .O(N__5313),
            .I(N__5304));
    LocalMux I__722 (
            .O(N__5310),
            .I(N__5301));
    IoSpan4Mux I__721 (
            .O(N__5307),
            .I(N__5298));
    IoSpan4Mux I__720 (
            .O(N__5304),
            .I(N__5295));
    IoSpan4Mux I__719 (
            .O(N__5301),
            .I(N__5292));
    Sp12to4 I__718 (
            .O(N__5298),
            .I(N__5289));
    Span4Mux_s2_h I__717 (
            .O(N__5295),
            .I(N__5286));
    IoSpan4Mux I__716 (
            .O(N__5292),
            .I(N__5283));
    Span12Mux_s9_v I__715 (
            .O(N__5289),
            .I(N__5280));
    Sp12to4 I__714 (
            .O(N__5286),
            .I(N__5277));
    Sp12to4 I__713 (
            .O(N__5283),
            .I(N__5274));
    Span12Mux_h I__712 (
            .O(N__5280),
            .I(N__5266));
    Span12Mux_h I__711 (
            .O(N__5277),
            .I(N__5266));
    Span12Mux_s9_v I__710 (
            .O(N__5274),
            .I(N__5266));
    InMux I__709 (
            .O(N__5273),
            .I(N__5263));
    Odrv12 I__708 (
            .O(N__5266),
            .I(TACK_EN));
    LocalMux I__707 (
            .O(N__5263),
            .I(TACK_EN));
    IoInMux I__706 (
            .O(N__5258),
            .I(N__5254));
    IoInMux I__705 (
            .O(N__5257),
            .I(N__5250));
    LocalMux I__704 (
            .O(N__5254),
            .I(N__5247));
    IoInMux I__703 (
            .O(N__5253),
            .I(N__5244));
    LocalMux I__702 (
            .O(N__5250),
            .I(N__5241));
    Span4Mux_s1_v I__701 (
            .O(N__5247),
            .I(N__5238));
    LocalMux I__700 (
            .O(N__5244),
            .I(N__5235));
    IoSpan4Mux I__699 (
            .O(N__5241),
            .I(N__5232));
    Sp12to4 I__698 (
            .O(N__5238),
            .I(N__5229));
    Span4Mux_s2_h I__697 (
            .O(N__5235),
            .I(N__5226));
    Span4Mux_s0_v I__696 (
            .O(N__5232),
            .I(N__5223));
    Span12Mux_h I__695 (
            .O(N__5229),
            .I(N__5220));
    Sp12to4 I__694 (
            .O(N__5226),
            .I(N__5217));
    Sp12to4 I__693 (
            .O(N__5223),
            .I(N__5214));
    Span12Mux_v I__692 (
            .O(N__5220),
            .I(N__5206));
    Span12Mux_v I__691 (
            .O(N__5217),
            .I(N__5206));
    Span12Mux_v I__690 (
            .O(N__5214),
            .I(N__5206));
    InMux I__689 (
            .O(N__5213),
            .I(N__5203));
    Odrv12 I__688 (
            .O(N__5206),
            .I(TACK_OUTn));
    LocalMux I__687 (
            .O(N__5203),
            .I(TACK_OUTn));
    InMux I__686 (
            .O(N__5198),
            .I(bfn_10_9_0_));
    InMux I__685 (
            .O(N__5195),
            .I(N__5191));
    InMux I__684 (
            .O(N__5194),
            .I(N__5188));
    LocalMux I__683 (
            .O(N__5191),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_5 ));
    LocalMux I__682 (
            .O(N__5188),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_5 ));
    InMux I__681 (
            .O(N__5183),
            .I(N__5179));
    InMux I__680 (
            .O(N__5182),
            .I(N__5176));
    LocalMux I__679 (
            .O(N__5179),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_6 ));
    LocalMux I__678 (
            .O(N__5176),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_6 ));
    InMux I__677 (
            .O(N__5171),
            .I(N__5167));
    InMux I__676 (
            .O(N__5170),
            .I(N__5164));
    LocalMux I__675 (
            .O(N__5167),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_7 ));
    LocalMux I__674 (
            .O(N__5164),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_7 ));
    CascadeMux I__673 (
            .O(N__5159),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0_cascade_ ));
    IoInMux I__672 (
            .O(N__5156),
            .I(N__5153));
    LocalMux I__671 (
            .O(N__5153),
            .I(N__5150));
    IoSpan4Mux I__670 (
            .O(N__5150),
            .I(N__5147));
    IoSpan4Mux I__669 (
            .O(N__5147),
            .I(N__5144));
    Span4Mux_s3_v I__668 (
            .O(N__5144),
            .I(N__5141));
    Sp12to4 I__667 (
            .O(N__5141),
            .I(N__5137));
    InMux I__666 (
            .O(N__5140),
            .I(N__5134));
    Odrv12 I__665 (
            .O(N__5137),
            .I(LATCH_CLK_c));
    LocalMux I__664 (
            .O(N__5134),
            .I(LATCH_CLK_c));
    CascadeMux I__663 (
            .O(N__5129),
            .I(\U712_CHIP_RAM.N_144_cascade_ ));
    InMux I__662 (
            .O(N__5126),
            .I(N__5123));
    LocalMux I__661 (
            .O(N__5123),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_4 ));
    InMux I__660 (
            .O(N__5120),
            .I(N__5115));
    InMux I__659 (
            .O(N__5119),
            .I(N__5112));
    InMux I__658 (
            .O(N__5118),
            .I(N__5109));
    LocalMux I__657 (
            .O(N__5115),
            .I(\U712_REG_SM.N_163 ));
    LocalMux I__656 (
            .O(N__5112),
            .I(\U712_REG_SM.N_163 ));
    LocalMux I__655 (
            .O(N__5109),
            .I(\U712_REG_SM.N_163 ));
    IoInMux I__654 (
            .O(N__5102),
            .I(N__5098));
    IoInMux I__653 (
            .O(N__5101),
            .I(N__5095));
    LocalMux I__652 (
            .O(N__5098),
            .I(N__5092));
    LocalMux I__651 (
            .O(N__5095),
            .I(N__5089));
    IoSpan4Mux I__650 (
            .O(N__5092),
            .I(N__5085));
    Span4Mux_s2_v I__649 (
            .O(N__5089),
            .I(N__5082));
    IoInMux I__648 (
            .O(N__5088),
            .I(N__5079));
    Sp12to4 I__647 (
            .O(N__5085),
            .I(N__5076));
    Span4Mux_h I__646 (
            .O(N__5082),
            .I(N__5073));
    LocalMux I__645 (
            .O(N__5079),
            .I(N__5070));
    Span12Mux_s7_h I__644 (
            .O(N__5076),
            .I(N__5065));
    Sp12to4 I__643 (
            .O(N__5073),
            .I(N__5065));
    Span4Mux_s2_h I__642 (
            .O(N__5070),
            .I(N__5062));
    Span12Mux_v I__641 (
            .O(N__5065),
            .I(N__5059));
    Sp12to4 I__640 (
            .O(N__5062),
            .I(N__5056));
    Span12Mux_h I__639 (
            .O(N__5059),
            .I(N__5053));
    Span12Mux_v I__638 (
            .O(N__5056),
            .I(N__5050));
    Odrv12 I__637 (
            .O(N__5053),
            .I(CLK40_PLL_i_i));
    Odrv12 I__636 (
            .O(N__5050),
            .I(CLK40_PLL_i_i));
    CascadeMux I__635 (
            .O(N__5045),
            .I(\U712_CYCLE_TERM.N_51_cascade_ ));
    InMux I__634 (
            .O(N__5042),
            .I(N__5039));
    LocalMux I__633 (
            .O(N__5039),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    SRMux I__632 (
            .O(N__5036),
            .I(N__5033));
    LocalMux I__631 (
            .O(N__5033),
            .I(N__5029));
    SRMux I__630 (
            .O(N__5032),
            .I(N__5026));
    Span4Mux_h I__629 (
            .O(N__5029),
            .I(N__5023));
    LocalMux I__628 (
            .O(N__5026),
            .I(N__5020));
    Odrv4 I__627 (
            .O(N__5023),
            .I(\U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ));
    Odrv12 I__626 (
            .O(N__5020),
            .I(\U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ));
    InMux I__625 (
            .O(N__5015),
            .I(\U712_CHIP_RAM.un2_DBR_COUNT_cry_5 ));
    InMux I__624 (
            .O(N__5012),
            .I(\U712_CHIP_RAM.un2_DBR_COUNT_cry_6 ));
    CascadeMux I__623 (
            .O(N__5009),
            .I(N__5004));
    InMux I__622 (
            .O(N__5008),
            .I(N__5001));
    InMux I__621 (
            .O(N__5007),
            .I(N__4996));
    InMux I__620 (
            .O(N__5004),
            .I(N__4996));
    LocalMux I__619 (
            .O(N__5001),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ));
    LocalMux I__618 (
            .O(N__4996),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ));
    InMux I__617 (
            .O(N__4991),
            .I(N__4985));
    InMux I__616 (
            .O(N__4990),
            .I(N__4985));
    LocalMux I__615 (
            .O(N__4985),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ));
    InMux I__614 (
            .O(N__4982),
            .I(N__4979));
    LocalMux I__613 (
            .O(N__4979),
            .I(\U712_REG_SM.N_159 ));
    InMux I__612 (
            .O(N__4976),
            .I(N__4972));
    InMux I__611 (
            .O(N__4975),
            .I(N__4969));
    LocalMux I__610 (
            .O(N__4972),
            .I(N__4966));
    LocalMux I__609 (
            .O(N__4969),
            .I(N__4962));
    Span4Mux_v I__608 (
            .O(N__4966),
            .I(N__4959));
    InMux I__607 (
            .O(N__4965),
            .I(N__4956));
    Span4Mux_h I__606 (
            .O(N__4962),
            .I(N__4953));
    Odrv4 I__605 (
            .O(N__4959),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    LocalMux I__604 (
            .O(N__4956),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    Odrv4 I__603 (
            .O(N__4953),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    InMux I__602 (
            .O(N__4946),
            .I(N__4939));
    InMux I__601 (
            .O(N__4945),
            .I(N__4939));
    InMux I__600 (
            .O(N__4944),
            .I(N__4936));
    LocalMux I__599 (
            .O(N__4939),
            .I(\U712_REG_SM.N_109 ));
    LocalMux I__598 (
            .O(N__4936),
            .I(\U712_REG_SM.N_109 ));
    CascadeMux I__597 (
            .O(N__4931),
            .I(N__4928));
    InMux I__596 (
            .O(N__4928),
            .I(N__4925));
    LocalMux I__595 (
            .O(N__4925),
            .I(\U712_REG_SM.N_164 ));
    InMux I__594 (
            .O(N__4922),
            .I(N__4919));
    LocalMux I__593 (
            .O(N__4919),
            .I(\U712_REG_SM.N_80 ));
    InMux I__592 (
            .O(N__4916),
            .I(N__4908));
    CascadeMux I__591 (
            .O(N__4915),
            .I(N__4904));
    CascadeMux I__590 (
            .O(N__4914),
            .I(N__4899));
    CascadeMux I__589 (
            .O(N__4913),
            .I(N__4895));
    InMux I__588 (
            .O(N__4912),
            .I(N__4890));
    InMux I__587 (
            .O(N__4911),
            .I(N__4890));
    LocalMux I__586 (
            .O(N__4908),
            .I(N__4887));
    CascadeMux I__585 (
            .O(N__4907),
            .I(N__4882));
    InMux I__584 (
            .O(N__4904),
            .I(N__4879));
    InMux I__583 (
            .O(N__4903),
            .I(N__4872));
    InMux I__582 (
            .O(N__4902),
            .I(N__4872));
    InMux I__581 (
            .O(N__4899),
            .I(N__4872));
    InMux I__580 (
            .O(N__4898),
            .I(N__4869));
    InMux I__579 (
            .O(N__4895),
            .I(N__4866));
    LocalMux I__578 (
            .O(N__4890),
            .I(N__4863));
    Span4Mux_h I__577 (
            .O(N__4887),
            .I(N__4860));
    InMux I__576 (
            .O(N__4886),
            .I(N__4855));
    InMux I__575 (
            .O(N__4885),
            .I(N__4855));
    InMux I__574 (
            .O(N__4882),
            .I(N__4852));
    LocalMux I__573 (
            .O(N__4879),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__572 (
            .O(N__4872),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__571 (
            .O(N__4869),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__570 (
            .O(N__4866),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__569 (
            .O(N__4863),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__568 (
            .O(N__4860),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__567 (
            .O(N__4855),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__566 (
            .O(N__4852),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    CascadeMux I__565 (
            .O(N__4835),
            .I(N__4832));
    InMux I__564 (
            .O(N__4832),
            .I(N__4829));
    LocalMux I__563 (
            .O(N__4829),
            .I(\U712_REG_SM.N_96 ));
    CascadeMux I__562 (
            .O(N__4826),
            .I(N__4821));
    InMux I__561 (
            .O(N__4825),
            .I(N__4815));
    InMux I__560 (
            .O(N__4824),
            .I(N__4812));
    InMux I__559 (
            .O(N__4821),
            .I(N__4809));
    InMux I__558 (
            .O(N__4820),
            .I(N__4802));
    InMux I__557 (
            .O(N__4819),
            .I(N__4802));
    InMux I__556 (
            .O(N__4818),
            .I(N__4802));
    LocalMux I__555 (
            .O(N__4815),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__554 (
            .O(N__4812),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__553 (
            .O(N__4809),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__552 (
            .O(N__4802),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    CascadeMux I__551 (
            .O(N__4793),
            .I(\U712_REG_SM.N_96_cascade_ ));
    CascadeMux I__550 (
            .O(N__4790),
            .I(N__4786));
    InMux I__549 (
            .O(N__4789),
            .I(N__4780));
    InMux I__548 (
            .O(N__4786),
            .I(N__4777));
    InMux I__547 (
            .O(N__4785),
            .I(N__4772));
    InMux I__546 (
            .O(N__4784),
            .I(N__4772));
    InMux I__545 (
            .O(N__4783),
            .I(N__4769));
    LocalMux I__544 (
            .O(N__4780),
            .I(N__4766));
    LocalMux I__543 (
            .O(N__4777),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__542 (
            .O(N__4772),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__541 (
            .O(N__4769),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    Odrv4 I__540 (
            .O(N__4766),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    IoInMux I__539 (
            .O(N__4757),
            .I(N__4754));
    LocalMux I__538 (
            .O(N__4754),
            .I(N__4751));
    IoSpan4Mux I__537 (
            .O(N__4751),
            .I(N__4748));
    Sp12to4 I__536 (
            .O(N__4748),
            .I(N__4745));
    Span12Mux_v I__535 (
            .O(N__4745),
            .I(N__4741));
    CascadeMux I__534 (
            .O(N__4744),
            .I(N__4738));
    Span12Mux_h I__533 (
            .O(N__4741),
            .I(N__4735));
    InMux I__532 (
            .O(N__4738),
            .I(N__4732));
    Odrv12 I__531 (
            .O(N__4735),
            .I(UDSn_c));
    LocalMux I__530 (
            .O(N__4732),
            .I(UDSn_c));
    InMux I__529 (
            .O(N__4727),
            .I(N__4724));
    LocalMux I__528 (
            .O(N__4724),
            .I(U712_BYTE_ENABLE_UDS_0));
    InMux I__527 (
            .O(N__4721),
            .I(N__4718));
    LocalMux I__526 (
            .O(N__4718),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__525 (
            .O(N__4715),
            .I(N__4712));
    LocalMux I__524 (
            .O(N__4712),
            .I(\U712_REG_SM.N_166 ));
    IoInMux I__523 (
            .O(N__4709),
            .I(N__4706));
    LocalMux I__522 (
            .O(N__4706),
            .I(N__4703));
    Span4Mux_s3_v I__521 (
            .O(N__4703),
            .I(N__4700));
    Span4Mux_h I__520 (
            .O(N__4700),
            .I(N__4697));
    Span4Mux_h I__519 (
            .O(N__4697),
            .I(N__4694));
    Sp12to4 I__518 (
            .O(N__4694),
            .I(N__4691));
    Span12Mux_s10_v I__517 (
            .O(N__4691),
            .I(N__4687));
    InMux I__516 (
            .O(N__4690),
            .I(N__4684));
    Odrv12 I__515 (
            .O(N__4687),
            .I(LDSn_c));
    LocalMux I__514 (
            .O(N__4684),
            .I(LDSn_c));
    IoInMux I__513 (
            .O(N__4679),
            .I(N__4676));
    LocalMux I__512 (
            .O(N__4676),
            .I(N__4673));
    Span4Mux_s2_v I__511 (
            .O(N__4673),
            .I(N__4670));
    Span4Mux_v I__510 (
            .O(N__4670),
            .I(N__4667));
    Span4Mux_v I__509 (
            .O(N__4667),
            .I(N__4664));
    Span4Mux_v I__508 (
            .O(N__4664),
            .I(N__4660));
    InMux I__507 (
            .O(N__4663),
            .I(N__4657));
    Odrv4 I__506 (
            .O(N__4660),
            .I(DBDIR_c));
    LocalMux I__505 (
            .O(N__4657),
            .I(DBDIR_c));
    InMux I__504 (
            .O(N__4652),
            .I(N__4649));
    LocalMux I__503 (
            .O(N__4649),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_2 ));
    InMux I__502 (
            .O(N__4646),
            .I(\U712_CHIP_RAM.un2_DBR_COUNT_cry_1 ));
    InMux I__501 (
            .O(N__4643),
            .I(N__4640));
    LocalMux I__500 (
            .O(N__4640),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_3 ));
    InMux I__499 (
            .O(N__4637),
            .I(\U712_CHIP_RAM.un2_DBR_COUNT_cry_2 ));
    InMux I__498 (
            .O(N__4634),
            .I(N__4631));
    LocalMux I__497 (
            .O(N__4631),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_4 ));
    InMux I__496 (
            .O(N__4628),
            .I(\U712_CHIP_RAM.un2_DBR_COUNT_cry_3 ));
    InMux I__495 (
            .O(N__4625),
            .I(\U712_CHIP_RAM.un2_DBR_COUNT_cry_4 ));
    CascadeMux I__494 (
            .O(N__4622),
            .I(\U712_REG_SM.N_109_cascade_ ));
    CascadeMux I__493 (
            .O(N__4619),
            .I(\U712_REG_SM.STATE_COUNTc_0_0_cascade_ ));
    InMux I__492 (
            .O(N__4616),
            .I(N__4604));
    InMux I__491 (
            .O(N__4615),
            .I(N__4604));
    InMux I__490 (
            .O(N__4614),
            .I(N__4604));
    InMux I__489 (
            .O(N__4613),
            .I(N__4604));
    LocalMux I__488 (
            .O(N__4604),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    CascadeMux I__487 (
            .O(N__4601),
            .I(\U712_REG_SM.REG_CYCLE_0_sqmuxa_cascade_ ));
    InMux I__486 (
            .O(N__4598),
            .I(N__4594));
    InMux I__485 (
            .O(N__4597),
            .I(N__4591));
    LocalMux I__484 (
            .O(N__4594),
            .I(\U712_REG_SM.N_185 ));
    LocalMux I__483 (
            .O(N__4591),
            .I(\U712_REG_SM.N_185 ));
    InMux I__482 (
            .O(N__4586),
            .I(N__4582));
    InMux I__481 (
            .O(N__4585),
            .I(N__4576));
    LocalMux I__480 (
            .O(N__4582),
            .I(N__4573));
    InMux I__479 (
            .O(N__4581),
            .I(N__4570));
    InMux I__478 (
            .O(N__4580),
            .I(N__4565));
    InMux I__477 (
            .O(N__4579),
            .I(N__4565));
    LocalMux I__476 (
            .O(N__4576),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    Odrv4 I__475 (
            .O(N__4573),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__474 (
            .O(N__4570),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__473 (
            .O(N__4565),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    CascadeMux I__472 (
            .O(N__4556),
            .I(N__4553));
    InMux I__471 (
            .O(N__4553),
            .I(N__4550));
    LocalMux I__470 (
            .O(N__4550),
            .I(\U712_REG_SM.N_109_0 ));
    InMux I__469 (
            .O(N__4547),
            .I(N__4543));
    InMux I__468 (
            .O(N__4546),
            .I(N__4540));
    LocalMux I__467 (
            .O(N__4543),
            .I(\U712_REG_SM.N_105_0 ));
    LocalMux I__466 (
            .O(N__4540),
            .I(\U712_REG_SM.N_105_0 ));
    InMux I__465 (
            .O(N__4535),
            .I(N__4531));
    InMux I__464 (
            .O(N__4534),
            .I(N__4525));
    LocalMux I__463 (
            .O(N__4531),
            .I(N__4522));
    InMux I__462 (
            .O(N__4530),
            .I(N__4519));
    InMux I__461 (
            .O(N__4529),
            .I(N__4516));
    InMux I__460 (
            .O(N__4528),
            .I(N__4513));
    LocalMux I__459 (
            .O(N__4525),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    Odrv4 I__458 (
            .O(N__4522),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__457 (
            .O(N__4519),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__456 (
            .O(N__4516),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__455 (
            .O(N__4513),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    InMux I__454 (
            .O(N__4502),
            .I(N__4499));
    LocalMux I__453 (
            .O(N__4499),
            .I(N__4495));
    IoInMux I__452 (
            .O(N__4498),
            .I(N__4492));
    Span4Mux_h I__451 (
            .O(N__4495),
            .I(N__4489));
    LocalMux I__450 (
            .O(N__4492),
            .I(N__4486));
    Span4Mux_v I__449 (
            .O(N__4489),
            .I(N__4483));
    IoSpan4Mux I__448 (
            .O(N__4486),
            .I(N__4480));
    Span4Mux_v I__447 (
            .O(N__4483),
            .I(N__4477));
    IoSpan4Mux I__446 (
            .O(N__4480),
            .I(N__4474));
    IoSpan4Mux I__445 (
            .O(N__4477),
            .I(N__4469));
    IoSpan4Mux I__444 (
            .O(N__4474),
            .I(N__4469));
    Odrv4 I__443 (
            .O(N__4469),
            .I(C1_c));
    InMux I__442 (
            .O(N__4466),
            .I(N__4462));
    InMux I__441 (
            .O(N__4465),
            .I(N__4459));
    LocalMux I__440 (
            .O(N__4462),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    LocalMux I__439 (
            .O(N__4459),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    InMux I__438 (
            .O(N__4454),
            .I(N__4450));
    InMux I__437 (
            .O(N__4453),
            .I(N__4447));
    LocalMux I__436 (
            .O(N__4450),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    LocalMux I__435 (
            .O(N__4447),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    CascadeMux I__434 (
            .O(N__4442),
            .I(\U712_REG_SM.N_157_cascade_ ));
    InMux I__433 (
            .O(N__4439),
            .I(N__4436));
    LocalMux I__432 (
            .O(N__4436),
            .I(N__4432));
    InMux I__431 (
            .O(N__4435),
            .I(N__4429));
    Span4Mux_h I__430 (
            .O(N__4432),
            .I(N__4424));
    LocalMux I__429 (
            .O(N__4429),
            .I(N__4424));
    Span4Mux_v I__428 (
            .O(N__4424),
            .I(N__4421));
    Span4Mux_h I__427 (
            .O(N__4421),
            .I(N__4418));
    Sp12to4 I__426 (
            .O(N__4418),
            .I(N__4415));
    Odrv12 I__425 (
            .O(N__4415),
            .I(DBRn_c));
    IoInMux I__424 (
            .O(N__4412),
            .I(N__4409));
    LocalMux I__423 (
            .O(N__4409),
            .I(N__4406));
    IoSpan4Mux I__422 (
            .O(N__4406),
            .I(N__4403));
    Span4Mux_s3_v I__421 (
            .O(N__4403),
            .I(N__4400));
    Sp12to4 I__420 (
            .O(N__4400),
            .I(N__4397));
    Span12Mux_s11_v I__419 (
            .O(N__4397),
            .I(N__4393));
    InMux I__418 (
            .O(N__4396),
            .I(N__4390));
    Odrv12 I__417 (
            .O(N__4393),
            .I(REGENn_c));
    LocalMux I__416 (
            .O(N__4390),
            .I(REGENn_c));
    InMux I__415 (
            .O(N__4385),
            .I(N__4381));
    InMux I__414 (
            .O(N__4384),
            .I(N__4378));
    LocalMux I__413 (
            .O(N__4381),
            .I(\U712_REG_SM.START_RSTZ0 ));
    LocalMux I__412 (
            .O(N__4378),
            .I(\U712_REG_SM.START_RSTZ0 ));
    CascadeMux I__411 (
            .O(N__4373),
            .I(\U712_REG_SM.un6_REG_CYCLE_START_cascade_ ));
    InMux I__410 (
            .O(N__4370),
            .I(N__4367));
    LocalMux I__409 (
            .O(N__4367),
            .I(N__4364));
    Span12Mux_h I__408 (
            .O(N__4364),
            .I(N__4361));
    Span12Mux_v I__407 (
            .O(N__4361),
            .I(N__4358));
    Odrv12 I__406 (
            .O(N__4358),
            .I(REGSPACEn_c));
    IoInMux I__405 (
            .O(N__4355),
            .I(N__4352));
    LocalMux I__404 (
            .O(N__4352),
            .I(N__4349));
    IoSpan4Mux I__403 (
            .O(N__4349),
            .I(N__4346));
    IoSpan4Mux I__402 (
            .O(N__4346),
            .I(N__4343));
    Span4Mux_s3_h I__401 (
            .O(N__4343),
            .I(N__4339));
    InMux I__400 (
            .O(N__4342),
            .I(N__4336));
    Span4Mux_h I__399 (
            .O(N__4339),
            .I(N__4333));
    LocalMux I__398 (
            .O(N__4336),
            .I(N__4330));
    Sp12to4 I__397 (
            .O(N__4333),
            .I(N__4327));
    Span4Mux_v I__396 (
            .O(N__4330),
            .I(N__4324));
    Span12Mux_h I__395 (
            .O(N__4327),
            .I(N__4319));
    Sp12to4 I__394 (
            .O(N__4324),
            .I(N__4319));
    Span12Mux_h I__393 (
            .O(N__4319),
            .I(N__4316));
    Odrv12 I__392 (
            .O(N__4316),
            .I(C3_c));
    InMux I__391 (
            .O(N__4313),
            .I(N__4310));
    LocalMux I__390 (
            .O(N__4310),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__389 (
            .O(N__4307),
            .I(N__4304));
    LocalMux I__388 (
            .O(N__4304),
            .I(\U712_REG_SM.STATE_COUNT_1_sqmuxa_1 ));
    InMux I__387 (
            .O(N__4301),
            .I(N__4298));
    LocalMux I__386 (
            .O(N__4298),
            .I(\U712_REG_SM.N_188 ));
    IoInMux I__385 (
            .O(N__4295),
            .I(N__4292));
    LocalMux I__384 (
            .O(N__4292),
            .I(N__4289));
    Span4Mux_s1_h I__383 (
            .O(N__4289),
            .I(N__4286));
    Span4Mux_h I__382 (
            .O(N__4286),
            .I(N__4283));
    Odrv4 I__381 (
            .O(N__4283),
            .I(DBRn_c_i_0));
    IoInMux I__380 (
            .O(N__4280),
            .I(N__4277));
    LocalMux I__379 (
            .O(N__4277),
            .I(N__4274));
    Span4Mux_s3_v I__378 (
            .O(N__4274),
            .I(N__4271));
    Span4Mux_h I__377 (
            .O(N__4271),
            .I(N__4268));
    Odrv4 I__376 (
            .O(N__4268),
            .I(CLK80_PLL_i_i));
    InMux I__375 (
            .O(N__4265),
            .I(N__4262));
    LocalMux I__374 (
            .O(N__4262),
            .I(DBR_SYNCZ0Z_0));
    IoInMux I__373 (
            .O(N__4259),
            .I(N__4256));
    LocalMux I__372 (
            .O(N__4256),
            .I(N__4253));
    IoSpan4Mux I__371 (
            .O(N__4253),
            .I(N__4250));
    Span4Mux_s2_v I__370 (
            .O(N__4250),
            .I(N__4247));
    Sp12to4 I__369 (
            .O(N__4247),
            .I(N__4244));
    Span12Mux_v I__368 (
            .O(N__4244),
            .I(N__4241));
    Odrv12 I__367 (
            .O(N__4241),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__5628));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__5630));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__5624));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__5625));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__5623));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__5627));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__5622));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__5626));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_10_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_13_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__4498),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7688),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4295),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__4355),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_13_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_13_7  (
            .in0(N__9541),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10982),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_3_1_1.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_3_1_1.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_3_1_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_3_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10343),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_0_LC_5_13_1.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_5_13_1.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_5_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_5_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4439),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10337),
            .ce(),
            .sr(N__10953));
    defparam DBR_SYNC_1_LC_5_13_5.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_5_13_5.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_5_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_5_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4265),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10337),
            .ce(),
            .sr(N__10953));
    defparam DBRn_ibuf_RNIBAB_LC_5_14_4.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_5_14_4.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_5_14_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_5_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4435),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_LC_5_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_5_15_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_5_15_4 .LUT_INIT=16'b1111101110101010;
    LogicCell40 \U712_REG_SM.REGENn_LC_5_15_4  (
            .in0(N__4307),
            .in1(N__4301),
            .in2(N__4915),
            .in3(N__4396),
            .lcout(REGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10339),
            .ce(),
            .sr(N__10945));
    defparam \U712_REG_SM.START_RST_LC_6_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_6_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_6_12_4 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.START_RST_LC_6_12_4  (
            .in0(N__4385),
            .in1(N__4454),
            .in2(_gnd_net_),
            .in3(N__4535),
            .lcout(\U712_REG_SM.START_RSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10330),
            .ce(),
            .sr(N__10949));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(N__4384),
            .in2(_gnd_net_),
            .in3(N__4585),
            .lcout(),
            .ltout(\U712_REG_SM.un6_REG_CYCLE_START_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_6_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_6_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_6_13_1 .LUT_INIT=16'b1100000011000100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_6_13_1  (
            .in0(N__5405),
            .in1(N__7879),
            .in2(N__4373),
            .in3(N__4370),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10332),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_0_LC_6_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_6_14_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_6_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4342),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10336),
            .ce(),
            .sr(N__10938));
    defparam \U712_REG_SM.C3_SYNC_1_LC_6_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_6_14_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_6_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4313),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10336),
            .ce(),
            .sr(N__10938));
    defparam \U712_REG_SM.REGENn_RNO_1_LC_6_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_RNO_1_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REGENn_RNO_1_LC_6_15_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_REG_SM.REGENn_RNO_1_LC_6_15_4  (
            .in0(N__4586),
            .in1(N__5513),
            .in2(N__4913),
            .in3(N__4976),
            .lcout(\U712_REG_SM.STATE_COUNT_1_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_RNO_0_LC_6_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_RNO_0_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REGENn_RNO_0_LC_6_15_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_REG_SM.REGENn_RNO_0_LC_6_15_6  (
            .in0(_gnd_net_),
            .in1(N__4530),
            .in2(_gnd_net_),
            .in3(N__5512),
            .lcout(\U712_REG_SM.N_188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_RNO_0_LC_6_16_1 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_6_16_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_6_16_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_REG_SM.LDSn_RNO_0_LC_6_16_1  (
            .in0(N__6774),
            .in1(N__6848),
            .in2(N__7002),
            .in3(N__10805),
            .lcout(\U712_REG_SM.N_166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.WRITE_CYCLE_LC_7_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_7_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_7_11_0 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_REG_SM.WRITE_CYCLE_LC_7_11_0  (
            .in0(N__10813),
            .in1(N__4466),
            .in2(_gnd_net_),
            .in3(N__4453),
            .lcout(\U712_REG_SM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10326),
            .ce(),
            .sr(N__10950));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_7_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_7_12_1 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_7_12_1  (
            .in0(N__5526),
            .in1(N__4912),
            .in2(_gnd_net_),
            .in3(N__4818),
            .lcout(\U712_REG_SM.N_164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_7_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_7_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_7_12_3  (
            .in0(N__4465),
            .in1(N__4820),
            .in2(_gnd_net_),
            .in3(N__4597),
            .lcout(\U712_REG_SM.N_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_7_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_7_12_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_7_12_5  (
            .in0(N__4579),
            .in1(N__4911),
            .in2(N__5534),
            .in3(N__4965),
            .lcout(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_7_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_7_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_7_12_6  (
            .in0(N__4819),
            .in1(N__4944),
            .in2(N__4790),
            .in3(N__4580),
            .lcout(\U712_REG_SM.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_7_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_7_13_0 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_7_13_0  (
            .in0(N__4614),
            .in1(N__4886),
            .in2(N__4826),
            .in3(N__6196),
            .lcout(),
            .ltout(\U712_REG_SM.N_157_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_7_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_7_13_1 .LUT_INIT=16'b0000100000001010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_7_13_1  (
            .in0(N__7878),
            .in1(N__5530),
            .in2(N__4442),
            .in3(N__4903),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10331),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_7_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_7_13_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_7_13_2  (
            .in0(N__4783),
            .in1(N__4885),
            .in2(_gnd_net_),
            .in3(N__5521),
            .lcout(\U712_REG_SM.N_185 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_7_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_7_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__4528),
            .in2(_gnd_net_),
            .in3(N__4613),
            .lcout(\U712_REG_SM.N_109 ),
            .ltout(\U712_REG_SM.N_109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_7_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_7_13_4 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_7_13_4  (
            .in0(N__4902),
            .in1(N__5523),
            .in2(N__4622),
            .in3(N__6198),
            .lcout(),
            .ltout(\U712_REG_SM.STATE_COUNTc_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_7_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_7_13_5 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_7_13_5  (
            .in0(N__7877),
            .in1(N__4547),
            .in2(N__4619),
            .in3(N__4616),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10331),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_7_13_6  (
            .in0(N__4615),
            .in1(N__5522),
            .in2(N__4914),
            .in3(N__6197),
            .lcout(),
            .ltout(\U712_REG_SM.REG_CYCLE_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_7_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_7_13_7 .LUT_INIT=16'b0100010011101100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_7_13_7  (
            .in0(N__7876),
            .in1(N__11634),
            .in2(N__4601),
            .in3(N__4598),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10331),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_7_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_7_14_0 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_7_14_0  (
            .in0(N__7880),
            .in1(N__4546),
            .in2(N__4556),
            .in3(N__4534),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10333),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_14_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_14_6  (
            .in0(N__5524),
            .in1(N__4975),
            .in2(_gnd_net_),
            .in3(N__4581),
            .lcout(\U712_REG_SM.N_109_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_7_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_7_14_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__4898),
            .in2(_gnd_net_),
            .in3(N__5525),
            .lcout(\U712_REG_SM.N_105_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_7_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_7_15_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_7_15_7  (
            .in0(N__4789),
            .in1(N__4529),
            .in2(N__4907),
            .in3(N__5488),
            .lcout(\U712_REG_SM.N_163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_0_LC_7_16_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_7_16_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_7_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4502),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10338),
            .ce(),
            .sr(N__10922));
    defparam \U712_REG_SM.C1_SYNC_1_LC_7_16_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_7_16_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_7_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4721),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10338),
            .ce(),
            .sr(N__10922));
    defparam \U712_REG_SM.LDSn_LC_7_16_7 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_7_16_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_7_16_7 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \U712_REG_SM.LDSn_LC_7_16_7  (
            .in0(N__4690),
            .in1(N__5120),
            .in2(N__5533),
            .in3(N__4715),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10338),
            .ce(),
            .sr(N__10922));
    defparam \U712_CHIP_RAM.DBDIR_LC_8_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_8_9_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_8_9_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_8_9_7  (
            .in0(N__6239),
            .in1(N__4663),
            .in2(_gnd_net_),
            .in3(N__5042),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10312),
            .ce(),
            .sr(N__10954));
    defparam \U712_CHIP_RAM.DBR_COUNT_0_LC_8_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_COUNT_0_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_0_LC_8_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_0_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5008),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10317),
            .ce(),
            .sr(N__5032));
    defparam \U712_CHIP_RAM.un2_DBR_COUNT_cry_1_c_LC_8_11_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.un2_DBR_COUNT_cry_1_c_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.un2_DBR_COUNT_cry_1_c_LC_8_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U712_CHIP_RAM.un2_DBR_COUNT_cry_1_c_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__4990),
            .in2(N__5009),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\U712_CHIP_RAM.un2_DBR_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBR_COUNT_2_LC_8_11_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_2_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_2_LC_8_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_2_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__4652),
            .in2(_gnd_net_),
            .in3(N__4646),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un2_DBR_COUNT_cry_1 ),
            .carryout(\U712_CHIP_RAM.un2_DBR_COUNT_cry_2 ),
            .clk(N__10323),
            .ce(),
            .sr(N__5036));
    defparam \U712_CHIP_RAM.DBR_COUNT_3_LC_8_11_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_3_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_3_LC_8_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_3_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__4643),
            .in2(_gnd_net_),
            .in3(N__4637),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un2_DBR_COUNT_cry_2 ),
            .carryout(\U712_CHIP_RAM.un2_DBR_COUNT_cry_3 ),
            .clk(N__10323),
            .ce(),
            .sr(N__5036));
    defparam \U712_CHIP_RAM.DBR_COUNT_4_LC_8_11_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_4_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_4_LC_8_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_4_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__4634),
            .in2(_gnd_net_),
            .in3(N__4628),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un2_DBR_COUNT_cry_3 ),
            .carryout(\U712_CHIP_RAM.un2_DBR_COUNT_cry_4 ),
            .clk(N__10323),
            .ce(),
            .sr(N__5036));
    defparam \U712_CHIP_RAM.DBR_COUNT_5_LC_8_11_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_5_LC_8_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_5_LC_8_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_5_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__5195),
            .in2(_gnd_net_),
            .in3(N__4625),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un2_DBR_COUNT_cry_4 ),
            .carryout(\U712_CHIP_RAM.un2_DBR_COUNT_cry_5 ),
            .clk(N__10323),
            .ce(),
            .sr(N__5036));
    defparam \U712_CHIP_RAM.DBR_COUNT_6_LC_8_11_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_6_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_6_LC_8_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_6_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__5183),
            .in2(_gnd_net_),
            .in3(N__5015),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un2_DBR_COUNT_cry_5 ),
            .carryout(\U712_CHIP_RAM.un2_DBR_COUNT_cry_6 ),
            .clk(N__10323),
            .ce(),
            .sr(N__5036));
    defparam \U712_CHIP_RAM.DBR_COUNT_7_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_COUNT_7_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_7_LC_8_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_7_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(N__5171),
            .in2(_gnd_net_),
            .in3(N__5012),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10323),
            .ce(),
            .sr(N__5036));
    defparam \U712_CHIP_RAM.DBR_COUNT_1_LC_8_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_COUNT_1_LC_8_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_1_LC_8_11_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_1_LC_8_11_7  (
            .in0(N__4991),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5007),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10323),
            .ce(),
            .sr(N__5036));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_12_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_12_1 .LUT_INIT=16'b1111111100000001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_8_12_1  (
            .in0(N__4946),
            .in1(N__4825),
            .in2(N__4835),
            .in3(N__4982),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10327),
            .ce(),
            .sr(N__10939));
    defparam \U712_REG_SM.REG_TACK_LC_8_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_8_12_6 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_8_12_6  (
            .in0(N__6273),
            .in1(N__4945),
            .in2(N__4931),
            .in3(N__4922),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10327),
            .ce(),
            .sr(N__10939));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_8_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_8_13_5 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_8_13_5  (
            .in0(N__4784),
            .in1(N__4916),
            .in2(_gnd_net_),
            .in3(N__5531),
            .lcout(\U712_REG_SM.N_96 ),
            .ltout(\U712_REG_SM.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_8_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_8_13_6 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_8_13_6  (
            .in0(N__7853),
            .in1(N__4824),
            .in2(N__4793),
            .in3(N__4785),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10329),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDSn_LC_8_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_8_15_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_8_15_3 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \U712_REG_SM.UDSn_LC_8_15_3  (
            .in0(N__4727),
            .in1(N__5119),
            .in2(N__4744),
            .in3(N__5517),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10334),
            .ce(),
            .sr(N__10923));
    defparam \U712_BYTE_ENABLE.UDS_LC_8_16_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UDS_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UDS_LC_8_16_0 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \U712_BYTE_ENABLE.UDS_LC_8_16_0  (
            .in0(N__6862),
            .in1(N__6971),
            .in2(N__6818),
            .in3(N__10806),
            .lcout(U712_BYTE_ENABLE_UDS_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_RNO_LC_8_16_6 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_8_16_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_REG_SM.ASn_ess_RNO_LC_8_16_6  (
            .in0(N__10980),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5118),
            .lcout(\U712_REG_SM.N_163_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pll_RNI8MQ3_LC_9_8_6.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_9_8_6.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_9_8_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 pll_RNI8MQ3_LC_9_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5901),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_9_2 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_9_2  (
            .in0(N__6036),
            .in1(N__6283),
            .in2(_gnd_net_),
            .in3(N__7090),
            .lcout(\U712_CYCLE_TERM.N_47_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_9_5 .LUT_INIT=16'b0000000000110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_9_5  (
            .in0(N__7091),
            .in1(N__6037),
            .in2(N__6287),
            .in3(N__6072),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_51_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_9_6 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_9_9_6  (
            .in0(N__6038),
            .in1(N__7850),
            .in2(N__5045),
            .in3(N__5888),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10308),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI1KG35_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI1KG35_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI1KG35_LC_9_9_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI1KG35_LC_9_9_7  (
            .in0(N__8011),
            .in1(N__7269),
            .in2(_gnd_net_),
            .in3(N__7394),
            .lcout(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_10_1 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_10_1  (
            .in0(N__5729),
            .in1(N__5546),
            .in2(_gnd_net_),
            .in3(N__7849),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10313),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_9_10_7 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_9_10_7  (
            .in0(N__6205),
            .in1(N__7848),
            .in2(_gnd_net_),
            .in3(N__6151),
            .lcout(\U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_11_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_11_1  (
            .in0(N__7792),
            .in1(N__7977),
            .in2(_gnd_net_),
            .in3(N__5804),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10318),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIGHLF1_0_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIGHLF1_0_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIGHLF1_0_LC_9_11_4 .LUT_INIT=16'b1010111011111111;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNIGHLF1_0_LC_9_11_4  (
            .in0(N__5727),
            .in1(N__5670),
            .in2(N__6157),
            .in3(N__7197),
            .lcout(\U712_CHIP_RAM.N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__7791),
            .in2(_gnd_net_),
            .in3(N__5671),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10318),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNO_0_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNO_0_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNO_0_LC_9_11_7 .LUT_INIT=16'b0000111100001000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNO_0_LC_9_11_7  (
            .in0(N__5194),
            .in1(N__5182),
            .in2(N__7307),
            .in3(N__5170),
            .lcout(\U712_CHIP_RAM.N_152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIF9JU1_2_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIF9JU1_2_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIF9JU1_2_LC_9_12_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIF9JU1_2_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__5740),
            .in2(_gnd_net_),
            .in3(N__8219),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_1_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_13_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_13_0  (
            .in0(N__5540),
            .in1(N__5993),
            .in2(N__8035),
            .in3(N__5126),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_9_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_9_13_1 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_9_13_1  (
            .in0(N__7851),
            .in1(N__5140),
            .in2(N__5159),
            .in3(N__5783),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10328),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_2_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_2_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_2_LC_9_13_2 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_2_LC_9_13_2  (
            .in0(N__8319),
            .in1(N__8112),
            .in2(_gnd_net_),
            .in3(N__8213),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_13_3 .LUT_INIT=16'b1111011111111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_13_3  (
            .in0(N__7852),
            .in1(N__8224),
            .in2(N__5129),
            .in3(N__7547),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_29_i_a2_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_3_LC_9_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_3_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_3_LC_9_13_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_3_LC_9_13_5  (
            .in0(N__6391),
            .in1(N__6373),
            .in2(N__6356),
            .in3(N__6331),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_2_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_2_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_2_LC_9_13_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_2_LC_9_13_6  (
            .in0(N__8320),
            .in1(N__8113),
            .in2(_gnd_net_),
            .in3(N__8214),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_9_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_9_13_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_9_13_7  (
            .in0(N__8212),
            .in1(N__7546),
            .in2(N__8121),
            .in3(N__8318),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER16_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_LC_9_16_0 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_LC_9_16_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_ess_LC_9_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.ASn_ess_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5532),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10335),
            .ce(N__5417),
            .sr(N__10913));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_20_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_20_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__5401),
            .in2(_gnd_net_),
            .in3(N__5375),
            .lcout(\U712_CHIP_RAM.un3_CPU_CYCLE_START ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_10_2_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_10_2_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_10_2_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_10_2_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_LC_10_6_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_LC_10_6_6  (
            .in0(N__9337),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11653),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_10_8_0 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_LC_10_8_0  (
            .in0(N__6085),
            .in1(N__5273),
            .in2(_gnd_net_),
            .in3(N__5330),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10304),
            .ce(),
            .sr(N__10951));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_8_7 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_8_7 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_10_8_7  (
            .in0(N__5213),
            .in1(N__6119),
            .in2(N__5903),
            .in3(N__6065),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10304),
            .ce(),
            .sr(N__10951));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_9_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_9_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__5558),
            .in2(_gnd_net_),
            .in3(N__5198),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__5629),
            .ce(),
            .sr(N__6023));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_9_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_9_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__5585),
            .in2(_gnd_net_),
            .in3(N__5651),
            .lcout(\U712_CHIP_RAM.REFRESH5lto1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__5629),
            .ce(),
            .sr(N__6023));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_9_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_9_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__5597),
            .in2(_gnd_net_),
            .in3(N__5648),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__5629),
            .ce(),
            .sr(N__6023));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_9_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_9_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__5704),
            .in2(_gnd_net_),
            .in3(N__5645),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__5629),
            .ce(),
            .sr(N__6023));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_9_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_9_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__5572),
            .in2(_gnd_net_),
            .in3(N__5642),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__5629),
            .ce(),
            .sr(N__6023));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_9_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_9_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__5753),
            .in2(_gnd_net_),
            .in3(N__5639),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__5629),
            .ce(),
            .sr(N__6023));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_9_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_9_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__5765),
            .in2(_gnd_net_),
            .in3(N__5636),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__5629),
            .ce(),
            .sr(N__6023));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_9_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_9_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__5777),
            .in2(_gnd_net_),
            .in3(N__5633),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5629),
            .ce(),
            .sr(N__6023));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_10_2 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_10_2  (
            .in0(N__5596),
            .in1(N__5584),
            .in2(N__5573),
            .in3(N__5557),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_10_10_4 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_10_10_4  (
            .in0(N__5728),
            .in1(N__8686),
            .in2(N__5675),
            .in3(N__6152),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_START_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_10_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_10_6  (
            .in0(N__5776),
            .in1(N__5764),
            .in2(_gnd_net_),
            .in3(N__5752),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_7 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_7  (
            .in0(N__7969),
            .in1(N__5741),
            .in2(_gnd_net_),
            .in3(N__7380),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_i_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNI2NL01_0_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNI2NL01_0_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNI2NL01_0_LC_10_11_0 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNI2NL01_0_LC_10_11_0  (
            .in0(N__6153),
            .in1(N__5726),
            .in2(_gnd_net_),
            .in3(N__5669),
            .lcout(\U712_CHIP_RAM.N_119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_11_1 .LUT_INIT=16'b0011000010110000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_10_11_1  (
            .in0(N__5705),
            .in1(N__5690),
            .in2(N__7820),
            .in3(N__5684),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10314),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGI6A1_2_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGI6A1_2_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGI6A1_2_LC_10_11_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIGI6A1_2_LC_10_11_2  (
            .in0(N__7785),
            .in1(N__7942),
            .in2(_gnd_net_),
            .in3(N__8198),
            .lcout(\U712_CHIP_RAM.N_187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_10_11_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_3_LC_10_11_3  (
            .in0(N__7636),
            .in1(N__8328),
            .in2(_gnd_net_),
            .in3(N__8448),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER18 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_10_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_10_11_4 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__7943),
            .in2(N__5678),
            .in3(N__7790),
            .lcout(\U712_CHIP_RAM.N_154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_11_5 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_10_11_5  (
            .in0(N__10580),
            .in1(N__7784),
            .in2(_gnd_net_),
            .in3(N__10667),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10314),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_10_11_6 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_10_11_6  (
            .in0(N__7145),
            .in1(N__8199),
            .in2(_gnd_net_),
            .in3(N__7618),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER33_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_11_7 .LUT_INIT=16'b0111111100110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_11_7  (
            .in0(N__7944),
            .in1(N__7786),
            .in2(N__5840),
            .in3(N__5789),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4HBB7_LC_10_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4HBB7_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4HBB7_LC_10_12_1 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI4HBB7_LC_10_12_1  (
            .in0(N__7968),
            .in1(N__7375),
            .in2(_gnd_net_),
            .in3(N__7617),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH3D4G_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH3D4G_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH3D4G_LC_10_12_2 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH3D4G_LC_10_12_2  (
            .in0(N__7973),
            .in1(N__5803),
            .in2(N__5837),
            .in3(N__6428),
            .lcout(\U712_CHIP_RAM.N_64 ),
            .ltout(\U712_CHIP_RAM.N_64_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_12_3 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_12_3  (
            .in0(N__6582),
            .in1(N__5978),
            .in2(N__5834),
            .in3(N__7172),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10319),
            .ce(N__5921),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIT7PC1_1_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIT7PC1_1_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIT7PC1_1_LC_10_12_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIT7PC1_1_LC_10_12_4  (
            .in0(N__8303),
            .in1(N__8092),
            .in2(_gnd_net_),
            .in3(N__8197),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER37_0_a3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_12_5 .LUT_INIT=16'b0001001011011110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_12_5  (
            .in0(N__5827),
            .in1(N__5951),
            .in2(N__7559),
            .in3(N__5810),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10319),
            .ce(N__5921),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_LC_10_12_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_LC_10_12_6  (
            .in0(N__8087),
            .in1(N__7537),
            .in2(_gnd_net_),
            .in3(N__8196),
            .lcout(\U712_CHIP_RAM.N_177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_12_7 .LUT_INIT=16'b0011000011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_12_7  (
            .in0(N__5802),
            .in1(N__7579),
            .in2(N__8010),
            .in3(N__7374),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_cnst_ss0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_13_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_13_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_13_0  (
            .in0(_gnd_net_),
            .in1(N__7558),
            .in2(_gnd_net_),
            .in3(N__8687),
            .lcout(\U712_CHIP_RAM.LATCH_CLK_6 ),
            .ltout(),
            .carryin(bfn_10_13_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_13_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_13_1  (
            .in0(N__5952),
            .in1(N__8108),
            .in2(_gnd_net_),
            .in3(N__5981),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__10324),
            .ce(N__5920),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_13_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__8225),
            .in2(_gnd_net_),
            .in3(N__5969),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_13_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_13_3  (
            .in0(N__5953),
            .in1(N__8326),
            .in2(_gnd_net_),
            .in3(N__5966),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__10324),
            .ce(N__5920),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_13_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_13_4  (
            .in0(N__5948),
            .in1(N__6354),
            .in2(_gnd_net_),
            .in3(N__5963),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__10324),
            .ce(N__5920),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_13_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_13_5  (
            .in0(N__5954),
            .in1(N__6374),
            .in2(_gnd_net_),
            .in3(N__5960),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__10324),
            .ce(N__5920),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_13_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_13_6  (
            .in0(N__5949),
            .in1(N__6392),
            .in2(_gnd_net_),
            .in3(N__5957),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__10324),
            .ce(N__5920),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_13_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_13_7  (
            .in0(N__6332),
            .in1(N__5950),
            .in2(_gnd_net_),
            .in3(N__5924),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10324),
            .ce(N__5920),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIHHJP6_0_LC_10_14_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIHHJP6_0_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIHHJP6_0_LC_10_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIHHJP6_0_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6557),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UUBE_LC_10_17_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_LC_10_17_3 .LUT_INIT=16'b0101010010101000;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_LC_10_17_3  (
            .in0(N__7011),
            .in1(N__6932),
            .in2(N__6894),
            .in3(N__6817),
            .lcout(UUBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_8_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_11_8_1  (
            .in0(N__7845),
            .in1(N__5902),
            .in2(_gnd_net_),
            .in3(N__6073),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10298),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_8_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__7847),
            .in2(_gnd_net_),
            .in3(N__6118),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10298),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_8_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_11_8_5  (
            .in0(N__7846),
            .in1(_gnd_net_),
            .in2(N__6104),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10298),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_8_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_8_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__6117),
            .in2(_gnd_net_),
            .in3(N__6100),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_11_9_2 .LUT_INIT=16'b1111101010001010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_11_9_2  (
            .in0(N__9299),
            .in1(N__7148),
            .in2(N__8045),
            .in3(N__6452),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10305),
            .ce(),
            .sr(N__10940));
    defparam \U712_CHIP_RAM.DBENn_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_11_9_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_11_9_3 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_11_9_3  (
            .in0(N__6248),
            .in1(N__8703),
            .in2(N__7397),
            .in3(N__9983),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10305),
            .ce(),
            .sr(N__10940));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_9_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_9_4 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_9_4 .LUT_INIT=16'b0000111000001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_11_9_4  (
            .in0(N__6092),
            .in1(N__6086),
            .in2(N__6074),
            .in3(N__6254),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10305),
            .ce(),
            .sr(N__10940));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_10_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_10_0  (
            .in0(N__9768),
            .in1(N__9864),
            .in2(N__9698),
            .in3(N__9485),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_LC_11_10_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_LC_11_10_1 .LUT_INIT=16'b0101000111110011;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_LC_11_10_1  (
            .in0(N__6524),
            .in1(N__8654),
            .in2(N__10598),
            .in3(N__9249),
            .lcout(CLMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNITQTQ3_LC_11_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNITQTQ3_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNITQTQ3_LC_11_10_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNITQTQ3_LC_11_10_2  (
            .in0(N__10720),
            .in1(N__7560),
            .in2(N__6311),
            .in3(N__8475),
            .lcout(\U712_CHIP_RAM.LATCH_CLK_0_sqmuxa ),
            .ltout(\U712_CHIP_RAM.LATCH_CLK_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI17CI7_0_LC_11_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI17CI7_0_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI17CI7_0_LC_11_10_3 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI17CI7_0_LC_11_10_3  (
            .in0(N__8476),
            .in1(N__7565),
            .in2(N__6290),
            .in3(N__6310),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER38_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_10_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_10_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_10_4  (
            .in0(N__6282),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7080),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2RSLC_LC_11_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2RSLC_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2RSLC_LC_11_10_6 .LUT_INIT=16'b1000000011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2RSLC_LC_11_10_6  (
            .in0(N__7379),
            .in1(N__7247),
            .in2(N__8044),
            .in3(N__7146),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_10_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6242),
            .in3(N__10981),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_7_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIQJ661_LC_11_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIQJ661_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIQJ661_LC_11_11_0 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIQJ661_LC_11_11_0  (
            .in0(N__7656),
            .in1(N__7196),
            .in2(_gnd_net_),
            .in3(N__7299),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERlde_0_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_11_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_11_11_1 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_11_11_1  (
            .in0(N__10801),
            .in1(N__7248),
            .in2(_gnd_net_),
            .in3(N__6235),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_LC_11_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_LC_11_11_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_DISABLE_LC_11_11_2  (
            .in0(N__6209),
            .in1(N__6170),
            .in2(N__6161),
            .in3(N__7782),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_DISABLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10309),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_11_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_11_11_3 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_11_11_3  (
            .in0(N__10722),
            .in1(_gnd_net_),
            .in2(N__8125),
            .in3(N__9250),
            .lcout(\U712_CHIP_RAM.CLK_EN_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_11_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_11_11_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_11_11_5  (
            .in0(N__10721),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7554),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE4LR1_1_LC_11_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE4LR1_1_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE4LR1_1_LC_11_11_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIE4LR1_1_LC_11_11_6  (
            .in0(N__8220),
            .in1(N__8009),
            .in2(N__6434),
            .in3(N__8117),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIEL6M4_3_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIEL6M4_3_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIEL6M4_3_LC_11_11_7 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIEL6M4_3_LC_11_11_7  (
            .in0(N__7783),
            .in1(N__8337),
            .in2(N__6431),
            .in3(N__8465),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_i_0_68_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_11_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_11_12_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_11_12_0  (
            .in0(N__8471),
            .in1(N__8034),
            .in2(N__8238),
            .in3(N__6398),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_11_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_11_12_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_11_12_1 .LUT_INIT=16'b0000110011111100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__6409),
            .in2(N__6422),
            .in3(N__6599),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10315),
            .ce(),
            .sr(N__10924));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_11_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_11_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_11_12_2  (
            .in0(N__7545),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8302),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7MG83_1_LC_11_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7MG83_1_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7MG83_1_LC_11_12_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI7MG83_1_LC_11_12_3  (
            .in0(N__8301),
            .in1(N__8227),
            .in2(N__8474),
            .in3(N__8090),
            .lcout(\U712_CHIP_RAM.N_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_12_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_12_4  (
            .in0(N__6390),
            .in1(N__6372),
            .in2(N__6355),
            .in3(N__6330),
            .lcout(\U712_CHIP_RAM.N_331_3 ),
            .ltout(\U712_CHIP_RAM.N_331_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_11_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_11_12_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_11_12_5  (
            .in0(N__8297),
            .in1(N__8088),
            .in2(N__6314),
            .in3(N__7542),
            .lcout(\U712_CHIP_RAM.N_172 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU95J5_0_LC_11_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU95J5_0_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIU95J5_0_LC_11_12_6 .LUT_INIT=16'b0011101100111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIU95J5_0_LC_11_12_6  (
            .in0(N__7544),
            .in1(N__8457),
            .in2(N__6515),
            .in3(N__6306),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_11_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_11_12_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_11_12_7  (
            .in0(N__8200),
            .in1(N__7543),
            .in2(N__8327),
            .in3(N__8089),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_11_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_11_13_0 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_0_LC_11_13_0  (
            .in0(N__6461),
            .in1(N__7268),
            .in2(N__7395),
            .in3(N__9518),
            .lcout(),
            .ltout(\U712_CHIP_RAM.BANK0_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_LC_11_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_LC_11_13_1 .LUT_INIT=16'b0000111101001110;
    LogicCell40 \U712_CHIP_RAM.BANK0_LC_11_13_1  (
            .in0(N__8552),
            .in1(N__6490),
            .in2(N__6506),
            .in3(N__8515),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10320),
            .ce(),
            .sr(N__10917));
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_11_13_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_1_LC_11_13_2  (
            .in0(N__11297),
            .in1(N__6479),
            .in2(_gnd_net_),
            .in3(N__6448),
            .lcout(\U712_CHIP_RAM.A_m_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_3_LC_11_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_3_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_3_LC_11_13_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_1_3_LC_11_13_3  (
            .in0(N__8459),
            .in1(N__8330),
            .in2(N__8234),
            .in3(N__7118),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER15 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNI0NAU5_LC_11_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNI0NAU5_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNI0NAU5_LC_11_13_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNI0NAU5_LC_11_13_4  (
            .in0(N__7283),
            .in1(N__7267),
            .in2(N__6455),
            .in3(N__7208),
            .lcout(\U712_CHIP_RAM.A_m_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_11_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_11_13_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__8091),
            .in2(_gnd_net_),
            .in3(N__7541),
            .lcout(\U712_CHIP_RAM.N_94 ),
            .ltout(\U712_CHIP_RAM.N_94_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_3_LC_11_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_3_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_3_LC_11_13_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_3_LC_11_13_6  (
            .in0(N__8329),
            .in1(N__8215),
            .in2(N__6437),
            .in3(N__8458),
            .lcout(\U712_CHIP_RAM.N_173 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRU1VF_3_LC_11_14_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRU1VF_3_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRU1VF_3_LC_11_14_0 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRU1VF_3_LC_11_14_0  (
            .in0(N__6584),
            .in1(N__6556),
            .in2(N__6536),
            .in3(N__6542),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIG5PHK_LC_11_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIG5PHK_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIG5PHK_LC_11_14_1 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIG5PHK_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6587),
            .in3(N__8356),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIHHJP6_LC_11_14_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIHHJP6_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIHHJP6_LC_11_14_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNIHHJP6_LC_11_14_2  (
            .in0(N__6583),
            .in1(N__6566),
            .in2(N__7271),
            .in3(N__7619),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGELS1_2_LC_11_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGELS1_2_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGELS1_2_LC_11_14_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIGELS1_2_LC_11_14_3  (
            .in0(N__7854),
            .in1(N__7119),
            .in2(_gnd_net_),
            .in3(N__8226),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_3_LC_11_14_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_3_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_3_LC_11_14_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_3_LC_11_14_4  (
            .in0(N__8322),
            .in1(N__8015),
            .in2(N__6545),
            .in3(N__8473),
            .lcout(\U712_CHIP_RAM.N_155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_11_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_11_14_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_11_14_5  (
            .in0(N__8472),
            .in1(N__7120),
            .in2(_gnd_net_),
            .in3(N__8321),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_14_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_14_6 .LUT_INIT=16'b0000011000000111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_14_6  (
            .in0(N__9757),
            .in1(N__9624),
            .in2(N__9486),
            .in3(N__9839),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_CMA28_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_14_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_14_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_11_14_7  (
            .in0(N__10979),
            .in1(_gnd_net_),
            .in2(N__6527),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LMBE_i_LC_11_16_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LMBE_i_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LMBE_i_LC_11_16_1 .LUT_INIT=16'b1010111001011101;
    LogicCell40 \U712_BYTE_ENABLE.LMBE_i_LC_11_16_1  (
            .in0(N__7009),
            .in1(N__6934),
            .in2(N__6875),
            .in3(N__6822),
            .lcout(\U712_BYTE_ENABLE.N_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_i_LC_11_16_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_i_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_i_LC_11_16_2 .LUT_INIT=16'b1111100010101111;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_i_LC_11_16_2  (
            .in0(N__6933),
            .in1(N__6863),
            .in2(N__6824),
            .in3(N__7008),
            .lcout(\U712_BYTE_ENABLE.N_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_LC_11_16_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_LC_11_16_3 .LUT_INIT=16'b0100010010001010;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_LC_11_16_3  (
            .in0(N__7010),
            .in1(N__6935),
            .in2(N__6876),
            .in3(N__6823),
            .lcout(UMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_56_i_LC_11_18_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_56_i_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_56_i_LC_11_18_0 .LUT_INIT=16'b0001000100101010;
    LogicCell40 \U712_BYTE_ENABLE.N_56_i_LC_11_18_0  (
            .in0(N__7012),
            .in1(N__6930),
            .in2(N__6895),
            .in3(N__6815),
            .lcout(N_56_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_58_i_LC_11_18_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_58_i_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_58_i_LC_11_18_2 .LUT_INIT=16'b0101000110100010;
    LogicCell40 \U712_BYTE_ENABLE.N_58_i_LC_11_18_2  (
            .in0(N__7013),
            .in1(N__6931),
            .in2(N__6896),
            .in3(N__6816),
            .lcout(N_58_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DMA_LATCH_EN_LC_11_20_4 .C_ON=1'b0;
    defparam \U712_BUFFERS.DMA_LATCH_EN_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DMA_LATCH_EN_LC_11_20_4 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U712_BUFFERS.DMA_LATCH_EN_LC_11_20_4  (
            .in0(N__10661),
            .in1(N__10584),
            .in2(_gnd_net_),
            .in3(N__10738),
            .lcout(DMA_LATCH_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_9_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_9_0  (
            .in0(N__8042),
            .in1(N__7270),
            .in2(_gnd_net_),
            .in3(N__7396),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10297),
            .ce(N__6710),
            .sr(N__10930));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_10_2  (
            .in0(N__6701),
            .in1(N__6683),
            .in2(_gnd_net_),
            .in3(N__9660),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_10_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_10_3  (
            .in0(N__6668),
            .in1(_gnd_net_),
            .in2(N__9690),
            .in3(N__6647),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_10_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_10_4  (
            .in0(N__6632),
            .in1(N__6617),
            .in2(_gnd_net_),
            .in3(N__9659),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_12_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_12_11_0 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_12_11_0  (
            .in0(N__9313),
            .in1(N__6598),
            .in2(N__7472),
            .in3(N__10724),
            .lcout(\U712_CHIP_RAM.CPU_TACK_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNICP6N_LC_12_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNICP6N_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNICP6N_LC_12_11_2 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_DISABLE_RNICP6N_LC_12_11_2  (
            .in0(N__7300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7657),
            .lcout(\U712_CHIP_RAM.N_95 ),
            .ltout(\U712_CHIP_RAM.N_95_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNI1VCF5_LC_12_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNI1VCF5_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNI1VCF5_LC_12_11_3 .LUT_INIT=16'b1010101100000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNI1VCF5_LC_12_11_3  (
            .in0(N__7257),
            .in1(N__7204),
            .in2(N__7175),
            .in3(N__7616),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_3_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_3_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR7N96_2_LC_12_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR7N96_2_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIR7N96_2_LC_12_11_4 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIR7N96_2_LC_12_11_4  (
            .in0(N__8030),
            .in1(_gnd_net_),
            .in2(N__7160),
            .in3(N__8239),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_12_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_12_11_5 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_12_11_5  (
            .in0(N__7762),
            .in1(N__10725),
            .in2(N__7157),
            .in3(N__7154),
            .lcout(WRITE_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10306),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_12_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_12_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_12_11_6  (
            .in0(N__7147),
            .in1(N__7322),
            .in2(N__8043),
            .in3(N__7124),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER42_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_12_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_12_11_7 .LUT_INIT=16'b0000100010101000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_12_11_7  (
            .in0(N__7761),
            .in1(N__7084),
            .in2(N__7100),
            .in3(N__7097),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10306),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_12_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_12_0  (
            .in0(N__7064),
            .in1(N__7052),
            .in2(_gnd_net_),
            .in3(N__9629),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGMF8A_3_LC_12_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGMF8A_3_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGMF8A_3_LC_12_12_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIGMF8A_3_LC_12_12_1  (
            .in0(N__7614),
            .in1(N__7037),
            .in2(_gnd_net_),
            .in3(N__7480),
            .lcout(\U712_CHIP_RAM.N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_12_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_12_12_2 .LUT_INIT=16'b1010101000100000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_12_12_2  (
            .in0(N__7803),
            .in1(N__9303),
            .in2(N__7661),
            .in3(N__7676),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10307),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_12_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_12_12_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_3_LC_12_12_3  (
            .in0(N__8027),
            .in1(N__8342),
            .in2(N__7640),
            .in3(N__8467),
            .lcout(\U712_CHIP_RAM.N_151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_12_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_12_12_4 .LUT_INIT=16'b1100000001010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_12_12_4  (
            .in0(N__7409),
            .in1(N__7615),
            .in2(N__7583),
            .in3(N__8026),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER17_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_12_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_12_12_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__7564),
            .in2(_gnd_net_),
            .in3(N__7481),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER34 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_12_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_12_12_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_12_12_6  (
            .in0(N__10723),
            .in1(_gnd_net_),
            .in2(N__7460),
            .in3(N__8025),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_7_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_12_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_12_7  (
            .in0(N__9628),
            .in1(N__7457),
            .in2(_gnd_net_),
            .in3(N__7438),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI2MJA9_1_LC_12_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI2MJA9_1_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI2MJA9_1_LC_12_13_2 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI2MJA9_1_LC_12_13_2  (
            .in0(N__7418),
            .in1(N__7408),
            .in2(_gnd_net_),
            .in3(N__8466),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER17_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH9ULN_LC_12_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH9ULN_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH9ULN_LC_12_13_3 .LUT_INIT=16'b0001000010111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH9ULN_LC_12_13_3  (
            .in0(N__8028),
            .in1(N__7387),
            .in2(N__7325),
            .in3(N__7321),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER19_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER19_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI7JQ5O_LC_12_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI7JQ5O_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI7JQ5O_LC_12_13_4 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI7JQ5O_LC_12_13_4  (
            .in0(N__7806),
            .in1(_gnd_net_),
            .in2(N__7310),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_38_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_12_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_12_13_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_12_13_5  (
            .in0(N__8558),
            .in1(N__8551),
            .in2(N__8537),
            .in3(N__8534),
            .lcout(\U712_CHIP_RAM.N_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_13_6 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_12_13_6  (
            .in0(N__7804),
            .in1(N__8528),
            .in2(N__8516),
            .in3(N__8501),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10311),
            .ce(N__8492),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_12_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_12_13_7 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_12_13_7  (
            .in0(N__8500),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7805),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10311),
            .ce(N__8492),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_12_14_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_12_14_0 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_12_14_0  (
            .in0(N__7886),
            .in1(N__8477),
            .in2(_gnd_net_),
            .in3(N__8393),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_61_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_12_14_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_12_14_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_12_14_1  (
            .in0(N__8363),
            .in1(N__8378),
            .in2(N__8381),
            .in3(N__9758),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10316),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_12_14_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_12_14_4 .LUT_INIT=16'b1111000010110001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_12_14_4  (
            .in0(N__8377),
            .in1(N__8369),
            .in2(N__9863),
            .in3(N__8362),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10316),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_12_14_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_12_14_7 .LUT_INIT=16'b0001110011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_2_LC_12_14_7  (
            .in0(N__8338),
            .in1(N__8240),
            .in2(N__8126),
            .in3(N__8029),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_29_i_a2_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_4.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_4.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_17_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7812),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un3_CUMBEn_1_LC_13_10_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un3_CUMBEn_1_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un3_CUMBEn_1_LC_13_10_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_BYTE_ENABLE.un3_CUMBEn_1_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__8719),
            .in2(_gnd_net_),
            .in3(N__8679),
            .lcout(\U712_BYTE_ENABLE.un3_CUMBEnZ0Z_1 ),
            .ltout(\U712_BYTE_ENABLE.un3_CUMBEnZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_LC_13_10_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_LC_13_10_1 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_LC_13_10_1  (
            .in0(N__9308),
            .in1(N__8830),
            .in2(N__8801),
            .in3(N__10666),
            .lcout(CUMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_LC_13_10_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_LC_13_10_3 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_LC_13_10_3  (
            .in0(N__9309),
            .in1(N__8780),
            .in2(N__8753),
            .in3(N__10588),
            .lcout(CUUBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un3_CLLBEn_0_LC_13_10_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un3_CLLBEn_0_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un3_CLLBEn_0_LC_13_10_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_BYTE_ENABLE.un3_CLLBEn_0_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__8718),
            .in2(_gnd_net_),
            .in3(N__8678),
            .lcout(\U712_BYTE_ENABLE.un3_CLLBEnZ0Z_0 ),
            .ltout(\U712_BYTE_ENABLE.un3_CLLBEnZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_LC_13_10_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_LC_13_10_7 .LUT_INIT=16'b0111011100000111;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_LC_13_10_7  (
            .in0(N__9307),
            .in1(N__8645),
            .in2(N__8630),
            .in3(N__10665),
            .lcout(CLLBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_13_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_13_11_7  (
            .in0(N__8585),
            .in1(N__8963),
            .in2(_gnd_net_),
            .in3(N__9014),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10310),
            .ce(N__10177),
            .sr(N__10926));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_12_0 .LUT_INIT=16'b1100111110101111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_12_0  (
            .in0(N__11549),
            .in1(N__8992),
            .in2(N__9429),
            .in3(N__9324),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_13_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_13_12_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_13_12_1  (
            .in0(N__8579),
            .in1(_gnd_net_),
            .in2(N__9339),
            .in3(N__9896),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_12_2 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_13_12_2  (
            .in0(N__10399),
            .in1(_gnd_net_),
            .in2(N__9017),
            .in3(N__9643),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_12_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_12_3  (
            .in0(N__9642),
            .in1(N__9008),
            .in2(N__9342),
            .in3(N__11603),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_12_5 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_12_5  (
            .in0(N__8991),
            .in1(N__9420),
            .in2(N__9341),
            .in3(N__11548),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_12_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__9767),
            .in2(_gnd_net_),
            .in3(N__9856),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_12_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_12_7  (
            .in0(N__9641),
            .in1(N__8957),
            .in2(N__9340),
            .in3(N__9995),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_13_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_13_13_0  (
            .in0(N__8951),
            .in1(N__8933),
            .in2(_gnd_net_),
            .in3(N__9627),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_13_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_13_13_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_13_13_3  (
            .in0(N__9626),
            .in1(N__8915),
            .in2(_gnd_net_),
            .in3(N__8890),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_13_6 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_13_6  (
            .in0(N__9756),
            .in1(N__9625),
            .in2(_gnd_net_),
            .in3(N__9843),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_6_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_14_6_2  (
            .in0(N__9775),
            .in1(N__9706),
            .in2(N__9499),
            .in3(N__9868),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10294),
            .ce(N__10198),
            .sr(N__10956));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_14_6_3 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_14_6_3  (
            .in0(N__9436),
            .in1(N__9122),
            .in2(N__9344),
            .in3(N__9080),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10294),
            .ce(N__10198),
            .sr(N__10956));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_9_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_9_5  (
            .in0(N__11451),
            .in1(N__11234),
            .in2(_gnd_net_),
            .in3(N__11132),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11066),
            .ce(N__11025),
            .sr(N__10946));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_10_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_14_10_5  (
            .in0(N__11131),
            .in1(N__11233),
            .in2(_gnd_net_),
            .in3(N__11456),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__11023),
            .sr(N__10941));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_11_5  (
            .in0(N__11229),
            .in1(N__11366),
            .in2(_gnd_net_),
            .in3(N__10133),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11067),
            .ce(N__11021),
            .sr(N__10931));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_12_1 .LUT_INIT=16'b0000111100100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_12_1  (
            .in0(N__9044),
            .in1(N__9332),
            .in2(N__9705),
            .in3(N__10398),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_14_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_14_12_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_14_12_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(N__9035),
            .in2(N__9071),
            .in3(N__9068),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10321),
            .ce(N__10178),
            .sr(N__10927));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_14_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_14_12_4 .LUT_INIT=16'b0000111011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_14_12_4  (
            .in0(N__9331),
            .in1(N__9043),
            .in2(N__10411),
            .in3(N__9691),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_14_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_14_13_3 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_14_13_3  (
            .in0(N__9314),
            .in1(N__9029),
            .in2(N__9905),
            .in3(N__9670),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_14_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_14_13_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_14_13_4  (
            .in0(N__9669),
            .in1(N__9023),
            .in2(N__9343),
            .in3(N__9884),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_A20_LC_14_14_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_14_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_14_14_4 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_14_14_4  (
            .in0(N__11124),
            .in1(N__11288),
            .in2(N__9542),
            .in3(N__9514),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__10918));
    defparam \U712_CHIP_RAM.CRCSn_LC_15_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_15_5_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_15_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_15_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9500),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10295),
            .ce(),
            .sr(N__10962));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_15_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_15_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_15_6_5 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_15_6_5  (
            .in0(N__9437),
            .in1(N__9401),
            .in2(N__9338),
            .in3(N__11081),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10299),
            .ce(N__10199),
            .sr(N__10958));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_15_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_15_9_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(N__9333),
            .in2(_gnd_net_),
            .in3(N__9699),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_15_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_15_10_0 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_15_10_0  (
            .in0(N__9362),
            .in1(N__9306),
            .in2(N__9968),
            .in3(N__9686),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_10_1 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_15_10_1  (
            .in0(N__9304),
            .in1(N__9353),
            .in2(N__9703),
            .in3(N__9158),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_10_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_15_10_5  (
            .in0(N__9305),
            .in1(N__9173),
            .in2(N__9704),
            .in3(N__9164),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_11_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_11_2  (
            .in0(N__11365),
            .in1(N__11275),
            .in2(_gnd_net_),
            .in3(N__10132),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__11022),
            .sr(N__10942));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_15_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_15_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_15_12_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_15_12_0  (
            .in0(N__10464),
            .in1(N__11468),
            .in2(N__10435),
            .in3(N__9152),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10325),
            .ce(N__10190),
            .sr(N__10932));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_15_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_15_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_15_12_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_15_12_4  (
            .in0(N__10465),
            .in1(N__9878),
            .in2(N__10436),
            .in3(N__9956),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10325),
            .ce(N__10190),
            .sr(N__10932));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_15_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_15_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_15_12_7 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_15_12_7  (
            .in0(N__10425),
            .in1(N__10466),
            .in2(N__10004),
            .in3(N__9932),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10325),
            .ce(N__10190),
            .sr(N__10932));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_13_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_13_1  (
            .in0(N__11290),
            .in1(N__10081),
            .in2(_gnd_net_),
            .in3(N__10046),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__11026),
            .sr(N__10928));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_13_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_13_2  (
            .in0(N__10045),
            .in1(N__11593),
            .in2(_gnd_net_),
            .in3(N__11289),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__11026),
            .sr(N__10928));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_13_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_13_3  (
            .in0(N__11291),
            .in1(N__10131),
            .in2(_gnd_net_),
            .in3(N__10082),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__11026),
            .sr(N__10928));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_14_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_14_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_14_0  (
            .in0(N__10044),
            .in1(N__11287),
            .in2(_gnd_net_),
            .in3(N__11594),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11069),
            .ce(N__11028),
            .sr(N__10925));
    defparam \U712_CHIP_RAM.WEn_LC_16_2_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_16_2_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_16_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_16_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9869),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10293),
            .ce(),
            .sr(N__10966));
    defparam \U712_CHIP_RAM.RASn_LC_16_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_16_4_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_16_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_16_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9779),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10296),
            .ce(),
            .sr(N__10964));
    defparam \U712_CHIP_RAM.CASn_LC_16_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_16_5_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_16_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_16_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9707),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10300),
            .ce(),
            .sr(N__10963));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_16_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_16_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_16_10_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_16_10_0  (
            .in0(N__10455),
            .in1(N__11318),
            .in2(N__10438),
            .in3(N__10514),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10322),
            .ce(N__10197),
            .sr(N__10952));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_16_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_16_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_16_10_4 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_16_10_4  (
            .in0(N__10454),
            .in1(N__10493),
            .in2(N__10437),
            .in3(N__10088),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10322),
            .ce(N__10197),
            .sr(N__10952));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_16_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_16_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_16_10_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_16_10_6  (
            .in0(N__10456),
            .in1(N__11411),
            .in2(N__10439),
            .in3(N__10370),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10322),
            .ce(N__10197),
            .sr(N__10952));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_11_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_16_11_7  (
            .in0(N__10080),
            .in1(N__11274),
            .in2(_gnd_net_),
            .in3(N__10130),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11063),
            .ce(N__11024),
            .sr(N__10947));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_16_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_16_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_16_12_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_16_12_1  (
            .in0(N__11285),
            .in1(N__10079),
            .in2(_gnd_net_),
            .in3(N__10043),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11064),
            .ce(N__11027),
            .sr(N__10943));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_16_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_16_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_16_13_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_16_13_2  (
            .in0(N__11589),
            .in1(N__11283),
            .in2(_gnd_net_),
            .in3(N__11534),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__11029),
            .sr(N__10933));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_16_14_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_16_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_16_14_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_16_14_3  (
            .in0(N__11281),
            .in1(N__11523),
            .in2(_gnd_net_),
            .in3(N__11492),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__11032),
            .sr(N__10929));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_10_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_10_1  (
            .in0(N__11455),
            .in1(N__11286),
            .in2(_gnd_net_),
            .in3(N__11395),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__11030),
            .sr(N__10955));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_12_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_12_3  (
            .in0(N__11284),
            .in1(N__11402),
            .in2(_gnd_net_),
            .in3(N__11358),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__11031),
            .sr(N__10948));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_17_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_17_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_17_13_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_17_13_4  (
            .in0(N__11579),
            .in1(N__11282),
            .in2(_gnd_net_),
            .in3(N__11530),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11065),
            .ce(N__11033),
            .sr(N__10944));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_17_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_17_14_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_17_14_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_17_14_5  (
            .in0(N__11280),
            .in1(N__11522),
            .in2(_gnd_net_),
            .in3(N__11491),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11068),
            .ce(N__11035),
            .sr(N__10934));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_18_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_18_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_18_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_18_10_6  (
            .in0(N__11293),
            .in1(N__11447),
            .in2(_gnd_net_),
            .in3(N__11394),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11062),
            .ce(N__11034),
            .sr(N__10957));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_18_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_18_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_18_10_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_18_10_7  (
            .in0(N__11393),
            .in1(N__11292),
            .in2(_gnd_net_),
            .in3(N__11352),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11062),
            .ce(N__11034),
            .sr(N__10957));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_9_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_9_3  (
            .in0(N__11309),
            .in1(N__11279),
            .in2(_gnd_net_),
            .in3(N__11123),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11061),
            .ce(N__11036),
            .sr(N__10965));
    defparam \U712_BUFFERS.DRDDIR_LC_24_20_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_LC_24_20_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_LC_24_20_1 .LUT_INIT=16'b0100011100001111;
    LogicCell40 \U712_BUFFERS.DRDDIR_LC_24_20_1  (
            .in0(N__10814),
            .in1(N__10558),
            .in2(N__10745),
            .in3(N__10636),
            .lcout(DRDDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_DRDENn_LC_24_20_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_LC_24_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_LC_24_20_2 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_LC_24_20_2  (
            .in0(N__10637),
            .in1(_gnd_net_),
            .in2(N__10573),
            .in3(N__11654),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

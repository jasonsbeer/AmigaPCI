-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Feb 8 2025 11:10:31

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    A : in std_logic_vector(20 downto 0);
    RAMENn : out std_logic;
    TSn : in std_logic;
    DMA_LATCH : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__11113\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \N_1012_i\ : std_logic;
signal \bfn_7_5_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_a3_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_223_i_0_en_cascade_\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \U712_CYCLE_TERM.N_223_i_0_en_0\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \N_242\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \U712_CHIP_RAM.N_381_cascade_\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_16\ : std_logic;
signal \N_187_i\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_0_a3_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_273\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_328_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_332_cascade_\ : std_logic;
signal \U712_CHIP_RAM.A_m_2_20\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.A_m_2_20_cascade_\ : std_logic;
signal \U712_CHIP_RAM.BANK0_esr_RNOZ0Z_1_cascade_\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_10_0_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_e_1\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_243\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_REG_SM.N_225\ : std_logic;
signal \U712_REG_SM.N_225_cascade_\ : std_logic;
signal \U712_REG_SM.N_292\ : std_logic;
signal \U712_REG_SM.REG_TACK_RNOZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_i_0_3_cascade_\ : std_logic;
signal \U712_REG_SM.N_289\ : std_logic;
signal \U712_REG_SM.N_289_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U712_CHIP_RAM.N_261_cascade_\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.N_260\ : std_logic;
signal \U712_CHIP_RAM.N_342_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_381\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_1_cascade_\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.N_270_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_0_0_i_1\ : std_logic;
signal \U712_CHIP_RAM.N_211_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_87\ : std_logic;
signal \U712_CHIP_RAM.N_266\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a3_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_264\ : std_logic;
signal \U712_CHIP_RAM.N_264_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_36_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_209\ : std_logic;
signal \U712_CHIP_RAM.N_209_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_263\ : std_logic;
signal \U712_CHIP_RAM.N_246\ : std_logic;
signal \U712_CHIP_RAM.N_332\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_203\ : std_logic;
signal \U712_CHIP_RAM.N_203_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_3_0\ : std_logic;
signal \U712_CHIP_RAM.N_341\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_SYNCZ0Z_1\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_2\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_1_2_cascade_\ : std_logic;
signal \U712_REG_SM.N_245\ : std_logic;
signal \U712_REG_SM.N_215\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_215_cascade_\ : std_logic;
signal \U712_REG_SM.N_228_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_i_0_1_cascade_\ : std_logic;
signal \C1_c\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_347_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_284\ : std_logic;
signal \U712_CHIP_RAM.N_211\ : std_logic;
signal \U712_CHIP_RAM.N_64_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_64_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_340\ : std_logic;
signal \U712_CHIP_RAM.N_340_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_267\ : std_logic;
signal \U712_CHIP_RAM.N_281_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.N_207_i\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_1_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \bfn_10_8_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_36\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_285\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_a3_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.N_342\ : std_logic;
signal \U712_CHIP_RAM.N_328\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_2_i_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_2_i_2\ : std_logic;
signal \U712_REG_SM.N_210\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_248_cascade_\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0\ : std_logic;
signal \U712_REG_SM.DS_EN_RNOZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_300\ : std_logic;
signal \U712_REG_SM.N_228\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \A_c_10\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\ : std_logic;
signal \U712_REG_SM.ASn_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.N_226\ : std_logic;
signal \ASn_c\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \U712_CHIP_RAM.un5_DMA_CYCLE_START_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10_cascade_\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_BYTE_ENABLE.N_315_cascade_\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_iZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \U712_BYTE_ENABLE.N_311\ : std_logic;
signal \U712_BYTE_ENABLE.N_313\ : std_logic;
signal \N_170\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_iZ0Z_0\ : std_logic;
signal \N_174_i\ : std_logic;
signal \N_172_i\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLMBEn_iZ0Z_0\ : std_logic;
signal \N_176_i\ : std_logic;
signal \A_c_1\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \U712_BYTE_ENABLE.N_309_cascade_\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUUBEn_iZ0Z_0\ : std_logic;
signal \DS_ENm\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \N_168\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \DMA_LATCH_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    \RESETn_wire\ <= RESETn;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    DMA_LATCH <= \DMA_LATCH_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__3792\,
            RESETB => \N__7044\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11113\,
            DIN => \N__11112\,
            DOUT => \N__11111\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11113\,
            PADOUT => \N__11112\,
            PADIN => \N__11111\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9396\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11104\,
            DIN => \N__11103\,
            DOUT => \N__11102\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11104\,
            PADOUT => \N__11103\,
            PADIN => \N__11102\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11095\,
            DIN => \N__11094\,
            DOUT => \N__11093\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11095\,
            PADOUT => \N__11094\,
            PADIN => \N__11093\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8298\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11086\,
            DIN => \N__11085\,
            DOUT => \N__11084\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11086\,
            PADOUT => \N__11085\,
            PADIN => \N__11084\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4008\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11077\,
            DIN => \N__11076\,
            DOUT => \N__11075\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11077\,
            PADOUT => \N__11076\,
            PADIN => \N__11075\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11068\,
            DIN => \N__11067\,
            DOUT => \N__11066\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11068\,
            PADOUT => \N__11067\,
            PADIN => \N__11066\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11059\,
            DIN => \N__11058\,
            DOUT => \N__11057\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11059\,
            PADOUT => \N__11058\,
            PADIN => \N__11057\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11050\,
            DIN => \N__11049\,
            DOUT => \N__11048\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11050\,
            PADOUT => \N__11049\,
            PADIN => \N__11048\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11041\,
            DIN => \N__11040\,
            DOUT => \N__11039\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11041\,
            PADOUT => \N__11040\,
            PADIN => \N__11039\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11032\,
            DIN => \N__11031\,
            DOUT => \N__11030\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11032\,
            PADOUT => \N__11031\,
            PADIN => \N__11030\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11023\,
            DIN => \N__11022\,
            DOUT => \N__11021\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11023\,
            PADOUT => \N__11022\,
            PADIN => \N__11021\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11014\,
            DIN => \N__11013\,
            DOUT => \N__11012\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11014\,
            PADOUT => \N__11013\,
            PADIN => \N__11012\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7167\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11005\,
            DIN => \N__11004\,
            DOUT => \N__11003\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11005\,
            PADOUT => \N__11004\,
            PADIN => \N__11003\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10996\,
            DIN => \N__10995\,
            DOUT => \N__10994\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10996\,
            PADOUT => \N__10995\,
            PADIN => \N__10994\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4418\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10987\,
            DIN => \N__10986\,
            DOUT => \N__10985\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10987\,
            PADOUT => \N__10986\,
            PADIN => \N__10985\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10978\,
            DIN => \N__10977\,
            DOUT => \N__10976\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10978\,
            PADOUT => \N__10977\,
            PADIN => \N__10976\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10969\,
            DIN => \N__10968\,
            DOUT => \N__10967\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10969\,
            PADOUT => \N__10968\,
            PADIN => \N__10967\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3930\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10960\,
            DIN => \N__10959\,
            DOUT => \N__10958\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10960\,
            PADOUT => \N__10959\,
            PADIN => \N__10958\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10951\,
            DIN => \N__10950\,
            DOUT => \N__10949\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10951\,
            PADOUT => \N__10950\,
            PADIN => \N__10949\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10942\,
            DIN => \N__10941\,
            DOUT => \N__10940\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10942\,
            PADOUT => \N__10941\,
            PADIN => \N__10940\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7017\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10933\,
            DIN => \N__10932\,
            DOUT => \N__10931\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10933\,
            PADOUT => \N__10932\,
            PADIN => \N__10931\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10924\,
            DIN => \N__10923\,
            DOUT => \N__10922\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10924\,
            PADOUT => \N__10923\,
            PADIN => \N__10922\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8787\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10915\,
            DIN => \N__10914\,
            DOUT => \N__10913\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10915\,
            PADOUT => \N__10914\,
            PADIN => \N__10913\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10906\,
            DIN => \N__10905\,
            DOUT => \N__10904\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10906\,
            PADOUT => \N__10905\,
            PADIN => \N__10904\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10897\,
            DIN => \N__10896\,
            DOUT => \N__10895\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10897\,
            PADOUT => \N__10896\,
            PADIN => \N__10895\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10888\,
            DIN => \N__10887\,
            DOUT => \N__10886\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10888\,
            PADOUT => \N__10887\,
            PADIN => \N__10886\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10879\,
            DIN => \N__10878\,
            DOUT => \N__10877\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10879\,
            PADOUT => \N__10878\,
            PADIN => \N__10877\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10870\,
            DIN => \N__10869\,
            DOUT => \N__10868\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10870\,
            PADOUT => \N__10869\,
            PADIN => \N__10868\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10861\,
            DIN => \N__10860\,
            DOUT => \N__10859\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10861\,
            PADOUT => \N__10860\,
            PADIN => \N__10859\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10852\,
            DIN => \N__10851\,
            DOUT => \N__10850\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10852\,
            PADOUT => \N__10851\,
            PADIN => \N__10850\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10843\,
            DIN => \N__10842\,
            DOUT => \N__10841\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10843\,
            PADOUT => \N__10842\,
            PADIN => \N__10841\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10834\,
            DIN => \N__10833\,
            DOUT => \N__10832\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10834\,
            PADOUT => \N__10833\,
            PADIN => \N__10832\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10825\,
            DIN => \N__10824\,
            DOUT => \N__10823\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10825\,
            PADOUT => \N__10824\,
            PADIN => \N__10823\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10816\,
            DIN => \N__10815\,
            DOUT => \N__10814\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10816\,
            PADOUT => \N__10815\,
            PADIN => \N__10814\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10807\,
            DIN => \N__10806\,
            DOUT => \N__10805\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10807\,
            PADOUT => \N__10806\,
            PADIN => \N__10805\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10798\,
            DIN => \N__10797\,
            DOUT => \N__10796\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10798\,
            PADOUT => \N__10797\,
            PADIN => \N__10796\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9933\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10789\,
            DIN => \N__10788\,
            DOUT => \N__10787\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10789\,
            PADOUT => \N__10788\,
            PADIN => \N__10787\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7870\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10780\,
            DIN => \N__10779\,
            DOUT => \N__10778\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10780\,
            PADOUT => \N__10779\,
            PADIN => \N__10778\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10771\,
            DIN => \N__10770\,
            DOUT => \N__10769\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10771\,
            PADOUT => \N__10770\,
            PADIN => \N__10769\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7500\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10762\,
            DIN => \N__10761\,
            DOUT => \N__10760\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10762\,
            PADOUT => \N__10761\,
            PADIN => \N__10760\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10753\,
            DIN => \N__10752\,
            DOUT => \N__10751\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10753\,
            PADOUT => \N__10752\,
            PADIN => \N__10751\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4320\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10744\,
            DIN => \N__10743\,
            DOUT => \N__10742\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10744\,
            PADOUT => \N__10743\,
            PADIN => \N__10742\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7872\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10735\,
            DIN => \N__10734\,
            DOUT => \N__10733\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10735\,
            PADOUT => \N__10734\,
            PADIN => \N__10733\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3849\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10726\,
            DIN => \N__10725\,
            DOUT => \N__10724\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10726\,
            PADOUT => \N__10725\,
            PADIN => \N__10724\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10717\,
            DIN => \N__10716\,
            DOUT => \N__10715\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10717\,
            PADOUT => \N__10716\,
            PADIN => \N__10715\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7074\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10708\,
            DIN => \N__10707\,
            DOUT => \N__10706\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10708\,
            PADOUT => \N__10707\,
            PADIN => \N__10706\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6954\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10699\,
            DIN => \N__10698\,
            DOUT => \N__10697\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10699\,
            PADOUT => \N__10698\,
            PADIN => \N__10697\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10690\,
            DIN => \N__10689\,
            DOUT => \N__10688\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10690\,
            PADOUT => \N__10689\,
            PADIN => \N__10688\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10681\,
            DIN => \N__10680\,
            DOUT => \N__10679\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10681\,
            PADOUT => \N__10680\,
            PADIN => \N__10679\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__10672\,
            DIN => \N__10671\,
            DOUT => \N__10670\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10672\,
            PADOUT => \N__10671\,
            PADIN => \N__10670\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10663\,
            DIN => \N__10662\,
            DOUT => \N__10661\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10663\,
            PADOUT => \N__10662\,
            PADIN => \N__10661\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7029\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10654\,
            DIN => \N__10653\,
            DOUT => \N__10652\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10654\,
            PADOUT => \N__10653\,
            PADIN => \N__10652\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10645\,
            DIN => \N__10644\,
            DOUT => \N__10643\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10645\,
            PADOUT => \N__10644\,
            PADIN => \N__10643\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7871\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10636\,
            DIN => \N__10635\,
            DOUT => \N__10634\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10636\,
            PADOUT => \N__10635\,
            PADIN => \N__10634\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7224\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10627\,
            DIN => \N__10626\,
            DOUT => \N__10625\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10627\,
            PADOUT => \N__10626\,
            PADIN => \N__10625\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8487\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10618\,
            DIN => \N__10617\,
            DOUT => \N__10616\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10618\,
            PADOUT => \N__10617\,
            PADIN => \N__10616\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4122\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10609\,
            DIN => \N__10608\,
            DOUT => \N__10607\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10609\,
            PADOUT => \N__10608\,
            PADIN => \N__10607\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7428\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10600\,
            DIN => \N__10599\,
            DOUT => \N__10598\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10600\,
            PADOUT => \N__10599\,
            PADIN => \N__10598\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6468\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10591\,
            DIN => \N__10590\,
            DOUT => \N__10589\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10591\,
            PADOUT => \N__10590\,
            PADIN => \N__10589\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10582\,
            DIN => \N__10581\,
            DOUT => \N__10580\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10582\,
            PADOUT => \N__10581\,
            PADIN => \N__10580\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10573\,
            DIN => \N__10572\,
            DOUT => \N__10571\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10573\,
            PADOUT => \N__10572\,
            PADIN => \N__10571\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9795\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10564\,
            DIN => \N__10563\,
            DOUT => \N__10562\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10564\,
            PADOUT => \N__10563\,
            PADIN => \N__10562\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8229\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10555\,
            DIN => \N__10554\,
            DOUT => \N__10553\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10555\,
            PADOUT => \N__10554\,
            PADIN => \N__10553\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3891\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10546\,
            DIN => \N__10545\,
            DOUT => \N__10544\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10546\,
            PADOUT => \N__10545\,
            PADIN => \N__10544\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9909\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10537\,
            DIN => \N__10536\,
            DOUT => \N__10535\,
            PACKAGEPIN => \DMA_LATCH_wire\
        );

    \DMA_LATCH_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10537\,
            PADOUT => \N__10536\,
            PADIN => \N__10535\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10528\,
            DIN => \N__10527\,
            DOUT => \N__10526\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10528\,
            PADOUT => \N__10527\,
            PADIN => \N__10526\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10519\,
            DIN => \N__10518\,
            DOUT => \N__10517\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10519\,
            PADOUT => \N__10518\,
            PADIN => \N__10517\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10510\,
            DIN => \N__10509\,
            DOUT => \N__10508\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10510\,
            PADOUT => \N__10509\,
            PADIN => \N__10508\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10501\,
            DIN => \N__10500\,
            DOUT => \N__10499\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10501\,
            PADOUT => \N__10500\,
            PADIN => \N__10499\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10492\,
            DIN => \N__10491\,
            DOUT => \N__10490\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10492\,
            PADOUT => \N__10491\,
            PADIN => \N__10490\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6387\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10483\,
            DIN => \N__10482\,
            DOUT => \N__10481\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10483\,
            PADOUT => \N__10482\,
            PADIN => \N__10481\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10474\,
            DIN => \N__10473\,
            DOUT => \N__10472\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10474\,
            PADOUT => \N__10473\,
            PADIN => \N__10472\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9897\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10465\,
            DIN => \N__10464\,
            DOUT => \N__10463\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__10465\,
            PADOUT => \N__10464\,
            PADIN => \N__10463\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3831\,
            DIN0 => OPEN,
            DOUT0 => \N__4269\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10456\,
            DIN => \N__10455\,
            DOUT => \N__10454\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10456\,
            PADOUT => \N__10455\,
            PADIN => \N__10454\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6423\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10447\,
            DIN => \N__10446\,
            DOUT => \N__10445\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10447\,
            PADOUT => \N__10446\,
            PADIN => \N__10445\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10438\,
            DIN => \N__10437\,
            DOUT => \N__10436\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10438\,
            PADOUT => \N__10437\,
            PADIN => \N__10436\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10429\,
            DIN => \N__10428\,
            DOUT => \N__10427\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10429\,
            PADOUT => \N__10428\,
            PADIN => \N__10427\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6981\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10420\,
            DIN => \N__10419\,
            DOUT => \N__10418\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10420\,
            PADOUT => \N__10419\,
            PADIN => \N__10418\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10411\,
            DIN => \N__10410\,
            DOUT => \N__10409\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10411\,
            PADOUT => \N__10410\,
            PADIN => \N__10409\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10402\,
            DIN => \N__10401\,
            DOUT => \N__10400\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10402\,
            PADOUT => \N__10401\,
            PADIN => \N__10400\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10393\,
            DIN => \N__10392\,
            DOUT => \N__10391\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10393\,
            PADOUT => \N__10392\,
            PADIN => \N__10391\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10384\,
            DIN => \N__10383\,
            DOUT => \N__10382\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10384\,
            PADOUT => \N__10383\,
            PADIN => \N__10382\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6879\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10375\,
            DIN => \N__10374\,
            DOUT => \N__10373\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10375\,
            PADOUT => \N__10374\,
            PADIN => \N__10373\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10152\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10366\,
            DIN => \N__10365\,
            DOUT => \N__10364\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10366\,
            PADOUT => \N__10365\,
            PADIN => \N__10364\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4548\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10357\,
            DIN => \N__10356\,
            DOUT => \N__10355\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10357\,
            PADOUT => \N__10356\,
            PADIN => \N__10355\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10348\,
            DIN => \N__10347\,
            DOUT => \N__10346\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10348\,
            PADOUT => \N__10347\,
            PADIN => \N__10346\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10339\,
            DIN => \N__10338\,
            DOUT => \N__10337\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10339\,
            PADOUT => \N__10338\,
            PADIN => \N__10337\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6930\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2505\ : InMux
    port map (
            O => \N__10320\,
            I => \N__10316\
        );

    \I__2504\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10313\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10316\,
            I => \N__10308\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10313\,
            I => \N__10308\
        );

    \I__2501\ : Span12Mux_h
    port map (
            O => \N__10308\,
            I => \N__10304\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10307\,
            I => \N__10301\
        );

    \I__2499\ : Odrv12
    port map (
            O => \N__10304\,
            I => \DS_ENm\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__10301\,
            I => \DS_ENm\
        );

    \I__2497\ : InMux
    port map (
            O => \N__10296\,
            I => \N__10293\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10293\,
            I => \N__10288\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10281\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10291\,
            I => \N__10281\
        );

    \I__2493\ : Span4Mux_h
    port map (
            O => \N__10288\,
            I => \N__10278\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10287\,
            I => \N__10275\
        );

    \I__2491\ : InMux
    port map (
            O => \N__10286\,
            I => \N__10271\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10281\,
            I => \N__10268\
        );

    \I__2489\ : Span4Mux_v
    port map (
            O => \N__10278\,
            I => \N__10265\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__10275\,
            I => \N__10262\
        );

    \I__2487\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10259\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__10271\,
            I => \N__10254\
        );

    \I__2485\ : Sp12to4
    port map (
            O => \N__10268\,
            I => \N__10254\
        );

    \I__2484\ : Span4Mux_v
    port map (
            O => \N__10265\,
            I => \N__10249\
        );

    \I__2483\ : Span4Mux_v
    port map (
            O => \N__10262\,
            I => \N__10249\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__10259\,
            I => \N__10246\
        );

    \I__2481\ : Span12Mux_v
    port map (
            O => \N__10254\,
            I => \N__10239\
        );

    \I__2480\ : Sp12to4
    port map (
            O => \N__10249\,
            I => \N__10239\
        );

    \I__2479\ : Span12Mux_s10_v
    port map (
            O => \N__10246\,
            I => \N__10239\
        );

    \I__2478\ : Span12Mux_h
    port map (
            O => \N__10239\,
            I => \N__10236\
        );

    \I__2477\ : Odrv12
    port map (
            O => \N__10236\,
            I => \A_c_0\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__10233\,
            I => \N__10228\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__10232\,
            I => \N__10225\
        );

    \I__2474\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10222\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10228\,
            I => \N__10217\
        );

    \I__2472\ : InMux
    port map (
            O => \N__10225\,
            I => \N__10217\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__10222\,
            I => \N__10211\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__10217\,
            I => \N__10211\
        );

    \I__2469\ : InMux
    port map (
            O => \N__10216\,
            I => \N__10208\
        );

    \I__2468\ : Span4Mux_v
    port map (
            O => \N__10211\,
            I => \N__10204\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__10208\,
            I => \N__10201\
        );

    \I__2466\ : InMux
    port map (
            O => \N__10207\,
            I => \N__10197\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__10204\,
            I => \N__10194\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__10201\,
            I => \N__10191\
        );

    \I__2463\ : InMux
    port map (
            O => \N__10200\,
            I => \N__10188\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__10197\,
            I => \N__10185\
        );

    \I__2461\ : Sp12to4
    port map (
            O => \N__10194\,
            I => \N__10182\
        );

    \I__2460\ : Span4Mux_v
    port map (
            O => \N__10191\,
            I => \N__10179\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__10188\,
            I => \N__10176\
        );

    \I__2458\ : Span12Mux_v
    port map (
            O => \N__10185\,
            I => \N__10173\
        );

    \I__2457\ : Span12Mux_h
    port map (
            O => \N__10182\,
            I => \N__10170\
        );

    \I__2456\ : Sp12to4
    port map (
            O => \N__10179\,
            I => \N__10165\
        );

    \I__2455\ : Span12Mux_v
    port map (
            O => \N__10176\,
            I => \N__10165\
        );

    \I__2454\ : Span12Mux_v
    port map (
            O => \N__10173\,
            I => \N__10162\
        );

    \I__2453\ : Span12Mux_v
    port map (
            O => \N__10170\,
            I => \N__10157\
        );

    \I__2452\ : Span12Mux_h
    port map (
            O => \N__10165\,
            I => \N__10157\
        );

    \I__2451\ : Odrv12
    port map (
            O => \N__10162\,
            I => \SIZ_c_0\
        );

    \I__2450\ : Odrv12
    port map (
            O => \N__10157\,
            I => \SIZ_c_0\
        );

    \I__2449\ : IoInMux
    port map (
            O => \N__10152\,
            I => \N__10149\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__10149\,
            I => \N__10146\
        );

    \I__2447\ : Span12Mux_s6_v
    port map (
            O => \N__10146\,
            I => \N__10143\
        );

    \I__2446\ : Odrv12
    port map (
            O => \N__10143\,
            I => \N_168\
        );

    \I__2445\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10133\
        );

    \I__2444\ : InMux
    port map (
            O => \N__10139\,
            I => \N__10130\
        );

    \I__2443\ : InMux
    port map (
            O => \N__10138\,
            I => \N__10127\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10137\,
            I => \N__10124\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10121\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__10133\,
            I => \N__10112\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__10130\,
            I => \N__10105\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__10127\,
            I => \N__10102\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10124\,
            I => \N__10075\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__10121\,
            I => \N__10072\
        );

    \I__2435\ : SRMux
    port map (
            O => \N__10120\,
            I => \N__9993\
        );

    \I__2434\ : SRMux
    port map (
            O => \N__10119\,
            I => \N__9993\
        );

    \I__2433\ : SRMux
    port map (
            O => \N__10118\,
            I => \N__9993\
        );

    \I__2432\ : SRMux
    port map (
            O => \N__10117\,
            I => \N__9993\
        );

    \I__2431\ : SRMux
    port map (
            O => \N__10116\,
            I => \N__9993\
        );

    \I__2430\ : SRMux
    port map (
            O => \N__10115\,
            I => \N__9993\
        );

    \I__2429\ : Glb2LocalMux
    port map (
            O => \N__10112\,
            I => \N__9993\
        );

    \I__2428\ : SRMux
    port map (
            O => \N__10111\,
            I => \N__9993\
        );

    \I__2427\ : SRMux
    port map (
            O => \N__10110\,
            I => \N__9993\
        );

    \I__2426\ : SRMux
    port map (
            O => \N__10109\,
            I => \N__9993\
        );

    \I__2425\ : SRMux
    port map (
            O => \N__10108\,
            I => \N__9993\
        );

    \I__2424\ : Glb2LocalMux
    port map (
            O => \N__10105\,
            I => \N__9993\
        );

    \I__2423\ : Glb2LocalMux
    port map (
            O => \N__10102\,
            I => \N__9993\
        );

    \I__2422\ : SRMux
    port map (
            O => \N__10101\,
            I => \N__9993\
        );

    \I__2421\ : SRMux
    port map (
            O => \N__10100\,
            I => \N__9993\
        );

    \I__2420\ : SRMux
    port map (
            O => \N__10099\,
            I => \N__9993\
        );

    \I__2419\ : SRMux
    port map (
            O => \N__10098\,
            I => \N__9993\
        );

    \I__2418\ : SRMux
    port map (
            O => \N__10097\,
            I => \N__9993\
        );

    \I__2417\ : SRMux
    port map (
            O => \N__10096\,
            I => \N__9993\
        );

    \I__2416\ : SRMux
    port map (
            O => \N__10095\,
            I => \N__9993\
        );

    \I__2415\ : SRMux
    port map (
            O => \N__10094\,
            I => \N__9993\
        );

    \I__2414\ : SRMux
    port map (
            O => \N__10093\,
            I => \N__9993\
        );

    \I__2413\ : SRMux
    port map (
            O => \N__10092\,
            I => \N__9993\
        );

    \I__2412\ : SRMux
    port map (
            O => \N__10091\,
            I => \N__9993\
        );

    \I__2411\ : SRMux
    port map (
            O => \N__10090\,
            I => \N__9993\
        );

    \I__2410\ : SRMux
    port map (
            O => \N__10089\,
            I => \N__9993\
        );

    \I__2409\ : SRMux
    port map (
            O => \N__10088\,
            I => \N__9993\
        );

    \I__2408\ : SRMux
    port map (
            O => \N__10087\,
            I => \N__9993\
        );

    \I__2407\ : SRMux
    port map (
            O => \N__10086\,
            I => \N__9993\
        );

    \I__2406\ : SRMux
    port map (
            O => \N__10085\,
            I => \N__9993\
        );

    \I__2405\ : SRMux
    port map (
            O => \N__10084\,
            I => \N__9993\
        );

    \I__2404\ : SRMux
    port map (
            O => \N__10083\,
            I => \N__9993\
        );

    \I__2403\ : SRMux
    port map (
            O => \N__10082\,
            I => \N__9993\
        );

    \I__2402\ : SRMux
    port map (
            O => \N__10081\,
            I => \N__9993\
        );

    \I__2401\ : SRMux
    port map (
            O => \N__10080\,
            I => \N__9993\
        );

    \I__2400\ : SRMux
    port map (
            O => \N__10079\,
            I => \N__9993\
        );

    \I__2399\ : SRMux
    port map (
            O => \N__10078\,
            I => \N__9993\
        );

    \I__2398\ : Glb2LocalMux
    port map (
            O => \N__10075\,
            I => \N__9993\
        );

    \I__2397\ : Glb2LocalMux
    port map (
            O => \N__10072\,
            I => \N__9993\
        );

    \I__2396\ : GlobalMux
    port map (
            O => \N__9993\,
            I => \N__9990\
        );

    \I__2395\ : gio2CtrlBuf
    port map (
            O => \N__9990\,
            I => \RESETn_c_i_g\
        );

    \I__2394\ : InMux
    port map (
            O => \N__9987\,
            I => \N__9983\
        );

    \I__2393\ : CascadeMux
    port map (
            O => \N__9986\,
            I => \N__9979\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__9983\,
            I => \N__9976\
        );

    \I__2391\ : InMux
    port map (
            O => \N__9982\,
            I => \N__9973\
        );

    \I__2390\ : InMux
    port map (
            O => \N__9979\,
            I => \N__9970\
        );

    \I__2389\ : Span4Mux_h
    port map (
            O => \N__9976\,
            I => \N__9965\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__9973\,
            I => \N__9965\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__9970\,
            I => \N__9962\
        );

    \I__2386\ : Span4Mux_v
    port map (
            O => \N__9965\,
            I => \N__9959\
        );

    \I__2385\ : Span12Mux_v
    port map (
            O => \N__9962\,
            I => \N__9954\
        );

    \I__2384\ : Sp12to4
    port map (
            O => \N__9959\,
            I => \N__9954\
        );

    \I__2383\ : Span12Mux_h
    port map (
            O => \N__9954\,
            I => \N__9951\
        );

    \I__2382\ : Span12Mux_v
    port map (
            O => \N__9951\,
            I => \N__9948\
        );

    \I__2381\ : Odrv12
    port map (
            O => \N__9948\,
            I => \CASLn_c\
        );

    \I__2380\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9942\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__9942\,
            I => \U712_BYTE_ENABLE.N_311\
        );

    \I__2378\ : InMux
    port map (
            O => \N__9939\,
            I => \N__9936\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__9936\,
            I => \U712_BYTE_ENABLE.N_313\
        );

    \I__2376\ : IoInMux
    port map (
            O => \N__9933\,
            I => \N__9930\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__9930\,
            I => \N__9927\
        );

    \I__2374\ : Span4Mux_s2_v
    port map (
            O => \N__9927\,
            I => \N__9924\
        );

    \I__2373\ : Span4Mux_h
    port map (
            O => \N__9924\,
            I => \N__9921\
        );

    \I__2372\ : Span4Mux_v
    port map (
            O => \N__9921\,
            I => \N__9918\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__9918\,
            I => \N_170\
        );

    \I__2370\ : InMux
    port map (
            O => \N__9915\,
            I => \N__9912\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__9912\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_iZ0Z_0\
        );

    \I__2368\ : IoInMux
    port map (
            O => \N__9909\,
            I => \N__9906\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__9906\,
            I => \N__9903\
        );

    \I__2366\ : Span12Mux_s11_h
    port map (
            O => \N__9903\,
            I => \N__9900\
        );

    \I__2365\ : Odrv12
    port map (
            O => \N__9900\,
            I => \N_174_i\
        );

    \I__2364\ : IoInMux
    port map (
            O => \N__9897\,
            I => \N__9894\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__9894\,
            I => \N__9891\
        );

    \I__2362\ : IoSpan4Mux
    port map (
            O => \N__9891\,
            I => \N__9888\
        );

    \I__2361\ : Span4Mux_s3_h
    port map (
            O => \N__9888\,
            I => \N__9885\
        );

    \I__2360\ : Span4Mux_h
    port map (
            O => \N__9885\,
            I => \N__9882\
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__9882\,
            I => \N_172_i\
        );

    \I__2358\ : InMux
    port map (
            O => \N__9879\,
            I => \N__9872\
        );

    \I__2357\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9867\
        );

    \I__2356\ : InMux
    port map (
            O => \N__9877\,
            I => \N__9867\
        );

    \I__2355\ : CascadeMux
    port map (
            O => \N__9876\,
            I => \N__9864\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__9875\,
            I => \N__9861\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__9872\,
            I => \N__9855\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__9867\,
            I => \N__9855\
        );

    \I__2351\ : InMux
    port map (
            O => \N__9864\,
            I => \N__9852\
        );

    \I__2350\ : InMux
    port map (
            O => \N__9861\,
            I => \N__9849\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__9860\,
            I => \N__9846\
        );

    \I__2348\ : Span4Mux_v
    port map (
            O => \N__9855\,
            I => \N__9839\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__9852\,
            I => \N__9839\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__9849\,
            I => \N__9839\
        );

    \I__2345\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9836\
        );

    \I__2344\ : Span4Mux_h
    port map (
            O => \N__9839\,
            I => \N__9833\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__9836\,
            I => \N__9830\
        );

    \I__2342\ : Span4Mux_v
    port map (
            O => \N__9833\,
            I => \N__9827\
        );

    \I__2341\ : Span4Mux_h
    port map (
            O => \N__9830\,
            I => \N__9824\
        );

    \I__2340\ : Sp12to4
    port map (
            O => \N__9827\,
            I => \N__9821\
        );

    \I__2339\ : Span4Mux_v
    port map (
            O => \N__9824\,
            I => \N__9818\
        );

    \I__2338\ : Span12Mux_h
    port map (
            O => \N__9821\,
            I => \N__9815\
        );

    \I__2337\ : Sp12to4
    port map (
            O => \N__9818\,
            I => \N__9812\
        );

    \I__2336\ : Span12Mux_v
    port map (
            O => \N__9815\,
            I => \N__9809\
        );

    \I__2335\ : Span12Mux_v
    port map (
            O => \N__9812\,
            I => \N__9806\
        );

    \I__2334\ : Odrv12
    port map (
            O => \N__9809\,
            I => \SIZ_c_1\
        );

    \I__2333\ : Odrv12
    port map (
            O => \N__9806\,
            I => \SIZ_c_1\
        );

    \I__2332\ : InMux
    port map (
            O => \N__9801\,
            I => \N__9798\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__9798\,
            I => \U712_BYTE_ENABLE.un1_CLMBEn_iZ0Z_0\
        );

    \I__2330\ : IoInMux
    port map (
            O => \N__9795\,
            I => \N__9792\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__9792\,
            I => \N__9789\
        );

    \I__2328\ : IoSpan4Mux
    port map (
            O => \N__9789\,
            I => \N__9786\
        );

    \I__2327\ : Span4Mux_s1_h
    port map (
            O => \N__9786\,
            I => \N__9783\
        );

    \I__2326\ : Sp12to4
    port map (
            O => \N__9783\,
            I => \N__9780\
        );

    \I__2325\ : Span12Mux_v
    port map (
            O => \N__9780\,
            I => \N__9777\
        );

    \I__2324\ : Odrv12
    port map (
            O => \N__9777\,
            I => \N_176_i\
        );

    \I__2323\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9771\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__9771\,
            I => \N__9767\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__9770\,
            I => \N__9763\
        );

    \I__2320\ : Span4Mux_v
    port map (
            O => \N__9767\,
            I => \N__9759\
        );

    \I__2319\ : InMux
    port map (
            O => \N__9766\,
            I => \N__9756\
        );

    \I__2318\ : InMux
    port map (
            O => \N__9763\,
            I => \N__9751\
        );

    \I__2317\ : InMux
    port map (
            O => \N__9762\,
            I => \N__9751\
        );

    \I__2316\ : Span4Mux_v
    port map (
            O => \N__9759\,
            I => \N__9748\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__9756\,
            I => \N__9743\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__9751\,
            I => \N__9743\
        );

    \I__2313\ : Span4Mux_v
    port map (
            O => \N__9748\,
            I => \N__9740\
        );

    \I__2312\ : Sp12to4
    port map (
            O => \N__9743\,
            I => \N__9737\
        );

    \I__2311\ : Sp12to4
    port map (
            O => \N__9740\,
            I => \N__9732\
        );

    \I__2310\ : Span12Mux_v
    port map (
            O => \N__9737\,
            I => \N__9732\
        );

    \I__2309\ : Span12Mux_h
    port map (
            O => \N__9732\,
            I => \N__9729\
        );

    \I__2308\ : Odrv12
    port map (
            O => \N__9729\,
            I => \A_c_1\
        );

    \I__2307\ : CascadeMux
    port map (
            O => \N__9726\,
            I => \N__9719\
        );

    \I__2306\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9713\
        );

    \I__2305\ : InMux
    port map (
            O => \N__9724\,
            I => \N__9713\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__9723\,
            I => \N__9710\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__9722\,
            I => \N__9706\
        );

    \I__2302\ : InMux
    port map (
            O => \N__9719\,
            I => \N__9702\
        );

    \I__2301\ : InMux
    port map (
            O => \N__9718\,
            I => \N__9699\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__9713\,
            I => \N__9692\
        );

    \I__2299\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9689\
        );

    \I__2298\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9685\
        );

    \I__2297\ : InMux
    port map (
            O => \N__9706\,
            I => \N__9680\
        );

    \I__2296\ : InMux
    port map (
            O => \N__9705\,
            I => \N__9677\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__9702\,
            I => \N__9674\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__9699\,
            I => \N__9671\
        );

    \I__2293\ : InMux
    port map (
            O => \N__9698\,
            I => \N__9664\
        );

    \I__2292\ : InMux
    port map (
            O => \N__9697\,
            I => \N__9664\
        );

    \I__2291\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9664\
        );

    \I__2290\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9661\
        );

    \I__2289\ : Span4Mux_v
    port map (
            O => \N__9692\,
            I => \N__9655\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__9689\,
            I => \N__9655\
        );

    \I__2287\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9652\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__9685\,
            I => \N__9649\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__9684\,
            I => \N__9643\
        );

    \I__2284\ : InMux
    port map (
            O => \N__9683\,
            I => \N__9636\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__9680\,
            I => \N__9631\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__9677\,
            I => \N__9631\
        );

    \I__2281\ : Span4Mux_h
    port map (
            O => \N__9674\,
            I => \N__9622\
        );

    \I__2280\ : Span4Mux_v
    port map (
            O => \N__9671\,
            I => \N__9622\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__9664\,
            I => \N__9622\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__9661\,
            I => \N__9622\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__9660\,
            I => \N__9616\
        );

    \I__2276\ : Span4Mux_h
    port map (
            O => \N__9655\,
            I => \N__9610\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__9652\,
            I => \N__9610\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__9649\,
            I => \N__9607\
        );

    \I__2273\ : InMux
    port map (
            O => \N__9648\,
            I => \N__9602\
        );

    \I__2272\ : InMux
    port map (
            O => \N__9647\,
            I => \N__9602\
        );

    \I__2271\ : InMux
    port map (
            O => \N__9646\,
            I => \N__9599\
        );

    \I__2270\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9594\
        );

    \I__2269\ : InMux
    port map (
            O => \N__9642\,
            I => \N__9594\
        );

    \I__2268\ : InMux
    port map (
            O => \N__9641\,
            I => \N__9589\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9640\,
            I => \N__9589\
        );

    \I__2266\ : InMux
    port map (
            O => \N__9639\,
            I => \N__9586\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__9636\,
            I => \N__9583\
        );

    \I__2264\ : Span4Mux_v
    port map (
            O => \N__9631\,
            I => \N__9578\
        );

    \I__2263\ : Span4Mux_h
    port map (
            O => \N__9622\,
            I => \N__9578\
        );

    \I__2262\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9573\
        );

    \I__2261\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9573\
        );

    \I__2260\ : InMux
    port map (
            O => \N__9619\,
            I => \N__9570\
        );

    \I__2259\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9567\
        );

    \I__2258\ : InMux
    port map (
            O => \N__9615\,
            I => \N__9564\
        );

    \I__2257\ : Span4Mux_h
    port map (
            O => \N__9610\,
            I => \N__9561\
        );

    \I__2256\ : Sp12to4
    port map (
            O => \N__9607\,
            I => \N__9550\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__9602\,
            I => \N__9550\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__9599\,
            I => \N__9550\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__9594\,
            I => \N__9550\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__9589\,
            I => \N__9550\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__9586\,
            I => \N__9543\
        );

    \I__2250\ : Span4Mux_h
    port map (
            O => \N__9583\,
            I => \N__9543\
        );

    \I__2249\ : Span4Mux_h
    port map (
            O => \N__9578\,
            I => \N__9543\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__9573\,
            I => \CPU_CYCLEm\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__9570\,
            I => \CPU_CYCLEm\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__9567\,
            I => \CPU_CYCLEm\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__9564\,
            I => \CPU_CYCLEm\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__9561\,
            I => \CPU_CYCLEm\
        );

    \I__2243\ : Odrv12
    port map (
            O => \N__9550\,
            I => \CPU_CYCLEm\
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__9543\,
            I => \CPU_CYCLEm\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__9525\,
            I => \N__9519\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__9524\,
            I => \N__9515\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9510\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9507\
        );

    \I__2236\ : Span4Mux_v
    port map (
            O => \N__9519\,
            I => \N__9504\
        );

    \I__2235\ : InMux
    port map (
            O => \N__9518\,
            I => \N__9501\
        );

    \I__2234\ : InMux
    port map (
            O => \N__9515\,
            I => \N__9498\
        );

    \I__2233\ : InMux
    port map (
            O => \N__9514\,
            I => \N__9495\
        );

    \I__2232\ : InMux
    port map (
            O => \N__9513\,
            I => \N__9492\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9510\,
            I => \N__9489\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__9507\,
            I => \N__9486\
        );

    \I__2229\ : Sp12to4
    port map (
            O => \N__9504\,
            I => \N__9477\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__9501\,
            I => \N__9477\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__9498\,
            I => \N__9477\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9495\,
            I => \N__9477\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__9492\,
            I => \N__9473\
        );

    \I__2224\ : Span12Mux_s8_v
    port map (
            O => \N__9489\,
            I => \N__9470\
        );

    \I__2223\ : Span12Mux_v
    port map (
            O => \N__9486\,
            I => \N__9465\
        );

    \I__2222\ : Span12Mux_h
    port map (
            O => \N__9477\,
            I => \N__9465\
        );

    \I__2221\ : InMux
    port map (
            O => \N__9476\,
            I => \N__9462\
        );

    \I__2220\ : Span4Mux_h
    port map (
            O => \N__9473\,
            I => \N__9459\
        );

    \I__2219\ : Odrv12
    port map (
            O => \N__9470\,
            I => \DMA_CYCLEm\
        );

    \I__2218\ : Odrv12
    port map (
            O => \N__9465\,
            I => \DMA_CYCLEm\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__9462\,
            I => \DMA_CYCLEm\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__9459\,
            I => \DMA_CYCLEm\
        );

    \I__2215\ : InMux
    port map (
            O => \N__9450\,
            I => \N__9446\
        );

    \I__2214\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9443\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__9446\,
            I => \N__9439\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__9443\,
            I => \N__9436\
        );

    \I__2211\ : InMux
    port map (
            O => \N__9442\,
            I => \N__9433\
        );

    \I__2210\ : Span4Mux_v
    port map (
            O => \N__9439\,
            I => \N__9430\
        );

    \I__2209\ : Span4Mux_v
    port map (
            O => \N__9436\,
            I => \N__9427\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__9433\,
            I => \N__9424\
        );

    \I__2207\ : Sp12to4
    port map (
            O => \N__9430\,
            I => \N__9419\
        );

    \I__2206\ : Sp12to4
    port map (
            O => \N__9427\,
            I => \N__9419\
        );

    \I__2205\ : Span4Mux_v
    port map (
            O => \N__9424\,
            I => \N__9416\
        );

    \I__2204\ : Span12Mux_h
    port map (
            O => \N__9419\,
            I => \N__9413\
        );

    \I__2203\ : Sp12to4
    port map (
            O => \N__9416\,
            I => \N__9410\
        );

    \I__2202\ : Span12Mux_v
    port map (
            O => \N__9413\,
            I => \N__9407\
        );

    \I__2201\ : Span12Mux_v
    port map (
            O => \N__9410\,
            I => \N__9404\
        );

    \I__2200\ : Odrv12
    port map (
            O => \N__9407\,
            I => \CASUn_c\
        );

    \I__2199\ : Odrv12
    port map (
            O => \N__9404\,
            I => \CASUn_c\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__9399\,
            I => \U712_BYTE_ENABLE.N_309_cascade_\
        );

    \I__2197\ : IoInMux
    port map (
            O => \N__9396\,
            I => \N__9393\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__9393\,
            I => \N__9389\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9386\
        );

    \I__2194\ : IoSpan4Mux
    port map (
            O => \N__9389\,
            I => \N__9382\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__9386\,
            I => \N__9379\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9385\,
            I => \N__9376\
        );

    \I__2191\ : Sp12to4
    port map (
            O => \N__9382\,
            I => \N__9371\
        );

    \I__2190\ : Span4Mux_v
    port map (
            O => \N__9379\,
            I => \N__9368\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__9376\,
            I => \N__9365\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9362\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9374\,
            I => \N__9359\
        );

    \I__2186\ : Span12Mux_s7_v
    port map (
            O => \N__9371\,
            I => \N__9355\
        );

    \I__2185\ : Sp12to4
    port map (
            O => \N__9368\,
            I => \N__9346\
        );

    \I__2184\ : Sp12to4
    port map (
            O => \N__9365\,
            I => \N__9346\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__9362\,
            I => \N__9346\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__9359\,
            I => \N__9346\
        );

    \I__2181\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9343\
        );

    \I__2180\ : Odrv12
    port map (
            O => \N__9355\,
            I => \DBENn_c\
        );

    \I__2179\ : Odrv12
    port map (
            O => \N__9346\,
            I => \DBENn_c\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9343\,
            I => \DBENn_c\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9336\,
            I => \N__9333\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9333\,
            I => \U712_BYTE_ENABLE.un1_CUUBEn_iZ0Z_0\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9330\,
            I => \N__9325\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9319\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9319\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9325\,
            I => \N__9316\
        );

    \I__2171\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9313\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9319\,
            I => \N__9310\
        );

    \I__2169\ : Span4Mux_h
    port map (
            O => \N__9316\,
            I => \N__9305\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__9313\,
            I => \N__9305\
        );

    \I__2167\ : Span4Mux_v
    port map (
            O => \N__9310\,
            I => \N__9302\
        );

    \I__2166\ : Span4Mux_v
    port map (
            O => \N__9305\,
            I => \N__9299\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__9302\,
            I => \N__9296\
        );

    \I__2164\ : Span4Mux_v
    port map (
            O => \N__9299\,
            I => \N__9293\
        );

    \I__2163\ : Sp12to4
    port map (
            O => \N__9296\,
            I => \N__9290\
        );

    \I__2162\ : Sp12to4
    port map (
            O => \N__9293\,
            I => \N__9287\
        );

    \I__2161\ : Span12Mux_h
    port map (
            O => \N__9290\,
            I => \N__9284\
        );

    \I__2160\ : Span12Mux_h
    port map (
            O => \N__9287\,
            I => \N__9281\
        );

    \I__2159\ : Odrv12
    port map (
            O => \N__9284\,
            I => \DRA_c_4\
        );

    \I__2158\ : Odrv12
    port map (
            O => \N__9281\,
            I => \DRA_c_4\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9276\,
            I => \N__9273\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__9273\,
            I => \N__9268\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9263\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9271\,
            I => \N__9263\
        );

    \I__2153\ : Span4Mux_h
    port map (
            O => \N__9268\,
            I => \N__9258\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__9263\,
            I => \N__9258\
        );

    \I__2151\ : Span4Mux_v
    port map (
            O => \N__9258\,
            I => \N__9254\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9251\
        );

    \I__2149\ : Span4Mux_v
    port map (
            O => \N__9254\,
            I => \N__9248\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9251\,
            I => \N__9245\
        );

    \I__2147\ : Sp12to4
    port map (
            O => \N__9248\,
            I => \N__9240\
        );

    \I__2146\ : Span12Mux_v
    port map (
            O => \N__9245\,
            I => \N__9240\
        );

    \I__2145\ : Span12Mux_h
    port map (
            O => \N__9240\,
            I => \N__9237\
        );

    \I__2144\ : Odrv12
    port map (
            O => \N__9237\,
            I => \DRA_c_3\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9231\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9231\,
            I => \N__9228\
        );

    \I__2141\ : Span4Mux_h
    port map (
            O => \N__9228\,
            I => \N__9225\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__9225\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9217\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9214\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9211\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9217\,
            I => \N__9207\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__9214\,
            I => \N__9202\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9211\,
            I => \N__9202\
        );

    \I__2133\ : InMux
    port map (
            O => \N__9210\,
            I => \N__9199\
        );

    \I__2132\ : Span4Mux_v
    port map (
            O => \N__9207\,
            I => \N__9196\
        );

    \I__2131\ : Sp12to4
    port map (
            O => \N__9202\,
            I => \N__9191\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__9199\,
            I => \N__9191\
        );

    \I__2129\ : Sp12to4
    port map (
            O => \N__9196\,
            I => \N__9188\
        );

    \I__2128\ : Span12Mux_v
    port map (
            O => \N__9191\,
            I => \N__9185\
        );

    \I__2127\ : Span12Mux_h
    port map (
            O => \N__9188\,
            I => \N__9182\
        );

    \I__2126\ : Span12Mux_h
    port map (
            O => \N__9185\,
            I => \N__9179\
        );

    \I__2125\ : Odrv12
    port map (
            O => \N__9182\,
            I => \DRA_c_8\
        );

    \I__2124\ : Odrv12
    port map (
            O => \N__9179\,
            I => \DRA_c_8\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9174\,
            I => \N__9171\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9171\,
            I => \N__9168\
        );

    \I__2121\ : Span4Mux_h
    port map (
            O => \N__9168\,
            I => \N__9165\
        );

    \I__2120\ : Odrv4
    port map (
            O => \N__9165\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9162\,
            I => \N__9159\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9159\,
            I => \N__9155\
        );

    \I__2117\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9152\
        );

    \I__2116\ : Span4Mux_v
    port map (
            O => \N__9155\,
            I => \N__9149\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9152\,
            I => \N__9146\
        );

    \I__2114\ : Sp12to4
    port map (
            O => \N__9149\,
            I => \N__9143\
        );

    \I__2113\ : Span12Mux_v
    port map (
            O => \N__9146\,
            I => \N__9140\
        );

    \I__2112\ : Span12Mux_h
    port map (
            O => \N__9143\,
            I => \N__9137\
        );

    \I__2111\ : Span12Mux_h
    port map (
            O => \N__9140\,
            I => \N__9134\
        );

    \I__2110\ : Odrv12
    port map (
            O => \N__9137\,
            I => \RAS0n_c\
        );

    \I__2109\ : Odrv12
    port map (
            O => \N__9134\,
            I => \RAS0n_c\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9129\,
            I => \N__9126\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__9126\,
            I => \N__9115\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9125\,
            I => \N__9112\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__9124\,
            I => \N__9108\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__9123\,
            I => \N__9105\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__9122\,
            I => \N__9102\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__9121\,
            I => \N__9096\
        );

    \I__2101\ : CascadeMux
    port map (
            O => \N__9120\,
            I => \N__9093\
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__9119\,
            I => \N__9089\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__9118\,
            I => \N__9085\
        );

    \I__2098\ : Span4Mux_h
    port map (
            O => \N__9115\,
            I => \N__9080\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__9112\,
            I => \N__9077\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9111\,
            I => \N__9063\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9108\,
            I => \N__9063\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9105\,
            I => \N__9063\
        );

    \I__2093\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9063\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9063\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9100\,
            I => \N__9063\
        );

    \I__2090\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9060\
        );

    \I__2089\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9045\
        );

    \I__2088\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9045\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9045\
        );

    \I__2086\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9045\
        );

    \I__2085\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9045\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9085\,
            I => \N__9045\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9045\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__9083\,
            I => \N__9042\
        );

    \I__2081\ : Span4Mux_v
    port map (
            O => \N__9080\,
            I => \N__9035\
        );

    \I__2080\ : Span4Mux_v
    port map (
            O => \N__9077\,
            I => \N__9035\
        );

    \I__2079\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9032\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__9063\,
            I => \N__9029\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__9060\,
            I => \N__9026\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9045\,
            I => \N__9023\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9042\,
            I => \N__9018\
        );

    \I__2074\ : InMux
    port map (
            O => \N__9041\,
            I => \N__9018\
        );

    \I__2073\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9015\
        );

    \I__2072\ : Sp12to4
    port map (
            O => \N__9035\,
            I => \N__9011\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__9032\,
            I => \N__9008\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__9029\,
            I => \N__9003\
        );

    \I__2069\ : Span4Mux_h
    port map (
            O => \N__9026\,
            I => \N__9003\
        );

    \I__2068\ : Span4Mux_v
    port map (
            O => \N__9023\,
            I => \N__9000\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__9018\,
            I => \N__8995\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9015\,
            I => \N__8995\
        );

    \I__2065\ : InMux
    port map (
            O => \N__9014\,
            I => \N__8992\
        );

    \I__2064\ : Span12Mux_h
    port map (
            O => \N__9011\,
            I => \N__8983\
        );

    \I__2063\ : Span12Mux_v
    port map (
            O => \N__9008\,
            I => \N__8983\
        );

    \I__2062\ : Sp12to4
    port map (
            O => \N__9003\,
            I => \N__8983\
        );

    \I__2061\ : Sp12to4
    port map (
            O => \N__9000\,
            I => \N__8983\
        );

    \I__2060\ : Sp12to4
    port map (
            O => \N__8995\,
            I => \N__8978\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__8992\,
            I => \N__8978\
        );

    \I__2058\ : Span12Mux_v
    port map (
            O => \N__8983\,
            I => \N__8975\
        );

    \I__2057\ : Span12Mux_v
    port map (
            O => \N__8978\,
            I => \N__8972\
        );

    \I__2056\ : Span12Mux_h
    port map (
            O => \N__8975\,
            I => \N__8969\
        );

    \I__2055\ : Span12Mux_h
    port map (
            O => \N__8972\,
            I => \N__8966\
        );

    \I__2054\ : Odrv12
    port map (
            O => \N__8969\,
            I => \AGNUS_REV_c\
        );

    \I__2053\ : Odrv12
    port map (
            O => \N__8966\,
            I => \AGNUS_REV_c\
        );

    \I__2052\ : InMux
    port map (
            O => \N__8961\,
            I => \N__8957\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__8960\,
            I => \N__8954\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__8957\,
            I => \N__8951\
        );

    \I__2049\ : InMux
    port map (
            O => \N__8954\,
            I => \N__8948\
        );

    \I__2048\ : Span4Mux_h
    port map (
            O => \N__8951\,
            I => \N__8941\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__8948\,
            I => \N__8941\
        );

    \I__2046\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8938\
        );

    \I__2045\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8935\
        );

    \I__2044\ : Span4Mux_v
    port map (
            O => \N__8941\,
            I => \N__8932\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__8938\,
            I => \N__8927\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__8935\,
            I => \N__8927\
        );

    \I__2041\ : Sp12to4
    port map (
            O => \N__8932\,
            I => \N__8922\
        );

    \I__2040\ : Span12Mux_v
    port map (
            O => \N__8927\,
            I => \N__8922\
        );

    \I__2039\ : Span12Mux_h
    port map (
            O => \N__8922\,
            I => \N__8919\
        );

    \I__2038\ : Span12Mux_v
    port map (
            O => \N__8919\,
            I => \N__8916\
        );

    \I__2037\ : Odrv12
    port map (
            O => \N__8916\,
            I => \DRA_c_9\
        );

    \I__2036\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8910\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__8910\,
            I => \N__8907\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__8907\,
            I => \N__8904\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__8904\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2032\ : InMux
    port map (
            O => \N__8901\,
            I => \N__8898\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__8898\,
            I => \N__8890\
        );

    \I__2030\ : ClkMux
    port map (
            O => \N__8897\,
            I => \N__8877\
        );

    \I__2029\ : ClkMux
    port map (
            O => \N__8896\,
            I => \N__8877\
        );

    \I__2028\ : ClkMux
    port map (
            O => \N__8895\,
            I => \N__8877\
        );

    \I__2027\ : ClkMux
    port map (
            O => \N__8894\,
            I => \N__8877\
        );

    \I__2026\ : ClkMux
    port map (
            O => \N__8893\,
            I => \N__8877\
        );

    \I__2025\ : Glb2LocalMux
    port map (
            O => \N__8890\,
            I => \N__8877\
        );

    \I__2024\ : GlobalMux
    port map (
            O => \N__8877\,
            I => \N__8874\
        );

    \I__2023\ : gio2CtrlBuf
    port map (
            O => \N__8874\,
            I => \C3_c_g\
        );

    \I__2022\ : CEMux
    port map (
            O => \N__8871\,
            I => \N__8867\
        );

    \I__2021\ : CEMux
    port map (
            O => \N__8870\,
            I => \N__8863\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__8867\,
            I => \N__8860\
        );

    \I__2019\ : CEMux
    port map (
            O => \N__8866\,
            I => \N__8857\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__8863\,
            I => \N__8849\
        );

    \I__2017\ : Span4Mux_v
    port map (
            O => \N__8860\,
            I => \N__8849\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__8857\,
            I => \N__8849\
        );

    \I__2015\ : CEMux
    port map (
            O => \N__8856\,
            I => \N__8846\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__8849\,
            I => \N__8841\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__8846\,
            I => \N__8841\
        );

    \I__2012\ : Span4Mux_v
    port map (
            O => \N__8841\,
            I => \N__8838\
        );

    \I__2011\ : Odrv4
    port map (
            O => \N__8838\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__8835\,
            I => \N__8831\
        );

    \I__2009\ : InMux
    port map (
            O => \N__8834\,
            I => \N__8828\
        );

    \I__2008\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8825\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__8828\,
            I => \N__8822\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__8825\,
            I => \N__8818\
        );

    \I__2005\ : Span4Mux_v
    port map (
            O => \N__8822\,
            I => \N__8815\
        );

    \I__2004\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8810\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__8818\,
            I => \N__8807\
        );

    \I__2002\ : Span4Mux_h
    port map (
            O => \N__8815\,
            I => \N__8804\
        );

    \I__2001\ : InMux
    port map (
            O => \N__8814\,
            I => \N__8801\
        );

    \I__2000\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8798\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__8810\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__8807\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__8804\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__8801\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__8798\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1994\ : IoInMux
    port map (
            O => \N__8787\,
            I => \N__8784\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__8784\,
            I => \N__8781\
        );

    \I__1992\ : Span4Mux_s3_v
    port map (
            O => \N__8781\,
            I => \N__8778\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__8778\,
            I => \N__8775\
        );

    \I__1990\ : Span4Mux_h
    port map (
            O => \N__8775\,
            I => \N__8772\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__8772\,
            I => \CRCSn_c\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__8769\,
            I => \U712_BYTE_ENABLE.N_315_cascade_\
        );

    \I__1987\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8763\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8763\,
            I => \N__8760\
        );

    \I__1985\ : Span4Mux_v
    port map (
            O => \N__8760\,
            I => \N__8757\
        );

    \I__1984\ : Span4Mux_h
    port map (
            O => \N__8757\,
            I => \N__8754\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__8754\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_iZ0Z_0\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8751\,
            I => \N__8747\
        );

    \I__1981\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8744\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__8747\,
            I => \N__8739\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__8744\,
            I => \N__8739\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__8739\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1977\ : InMux
    port map (
            O => \N__8736\,
            I => \N__8733\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__8733\,
            I => \N__8707\
        );

    \I__1975\ : ClkMux
    port map (
            O => \N__8732\,
            I => \N__8628\
        );

    \I__1974\ : ClkMux
    port map (
            O => \N__8731\,
            I => \N__8628\
        );

    \I__1973\ : ClkMux
    port map (
            O => \N__8730\,
            I => \N__8628\
        );

    \I__1972\ : ClkMux
    port map (
            O => \N__8729\,
            I => \N__8628\
        );

    \I__1971\ : ClkMux
    port map (
            O => \N__8728\,
            I => \N__8628\
        );

    \I__1970\ : ClkMux
    port map (
            O => \N__8727\,
            I => \N__8628\
        );

    \I__1969\ : ClkMux
    port map (
            O => \N__8726\,
            I => \N__8628\
        );

    \I__1968\ : ClkMux
    port map (
            O => \N__8725\,
            I => \N__8628\
        );

    \I__1967\ : ClkMux
    port map (
            O => \N__8724\,
            I => \N__8628\
        );

    \I__1966\ : ClkMux
    port map (
            O => \N__8723\,
            I => \N__8628\
        );

    \I__1965\ : ClkMux
    port map (
            O => \N__8722\,
            I => \N__8628\
        );

    \I__1964\ : ClkMux
    port map (
            O => \N__8721\,
            I => \N__8628\
        );

    \I__1963\ : ClkMux
    port map (
            O => \N__8720\,
            I => \N__8628\
        );

    \I__1962\ : ClkMux
    port map (
            O => \N__8719\,
            I => \N__8628\
        );

    \I__1961\ : ClkMux
    port map (
            O => \N__8718\,
            I => \N__8628\
        );

    \I__1960\ : ClkMux
    port map (
            O => \N__8717\,
            I => \N__8628\
        );

    \I__1959\ : ClkMux
    port map (
            O => \N__8716\,
            I => \N__8628\
        );

    \I__1958\ : ClkMux
    port map (
            O => \N__8715\,
            I => \N__8628\
        );

    \I__1957\ : ClkMux
    port map (
            O => \N__8714\,
            I => \N__8628\
        );

    \I__1956\ : ClkMux
    port map (
            O => \N__8713\,
            I => \N__8628\
        );

    \I__1955\ : ClkMux
    port map (
            O => \N__8712\,
            I => \N__8628\
        );

    \I__1954\ : ClkMux
    port map (
            O => \N__8711\,
            I => \N__8628\
        );

    \I__1953\ : ClkMux
    port map (
            O => \N__8710\,
            I => \N__8628\
        );

    \I__1952\ : Glb2LocalMux
    port map (
            O => \N__8707\,
            I => \N__8628\
        );

    \I__1951\ : ClkMux
    port map (
            O => \N__8706\,
            I => \N__8628\
        );

    \I__1950\ : ClkMux
    port map (
            O => \N__8705\,
            I => \N__8628\
        );

    \I__1949\ : ClkMux
    port map (
            O => \N__8704\,
            I => \N__8628\
        );

    \I__1948\ : ClkMux
    port map (
            O => \N__8703\,
            I => \N__8628\
        );

    \I__1947\ : ClkMux
    port map (
            O => \N__8702\,
            I => \N__8628\
        );

    \I__1946\ : ClkMux
    port map (
            O => \N__8701\,
            I => \N__8628\
        );

    \I__1945\ : ClkMux
    port map (
            O => \N__8700\,
            I => \N__8628\
        );

    \I__1944\ : ClkMux
    port map (
            O => \N__8699\,
            I => \N__8628\
        );

    \I__1943\ : ClkMux
    port map (
            O => \N__8698\,
            I => \N__8628\
        );

    \I__1942\ : ClkMux
    port map (
            O => \N__8697\,
            I => \N__8628\
        );

    \I__1941\ : GlobalMux
    port map (
            O => \N__8628\,
            I => \CLK80_PLL\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8622\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__8622\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1938\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8616\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__8616\,
            I => \N__8613\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__8613\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1935\ : InMux
    port map (
            O => \N__8610\,
            I => \N__8602\
        );

    \I__1934\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8602\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8608\,
            I => \N__8599\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8607\,
            I => \N__8596\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__8602\,
            I => \N__8589\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__8599\,
            I => \N__8589\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__8596\,
            I => \N__8589\
        );

    \I__1928\ : Span4Mux_v
    port map (
            O => \N__8589\,
            I => \N__8586\
        );

    \I__1927\ : Sp12to4
    port map (
            O => \N__8586\,
            I => \N__8583\
        );

    \I__1926\ : Span12Mux_h
    port map (
            O => \N__8583\,
            I => \N__8580\
        );

    \I__1925\ : Odrv12
    port map (
            O => \N__8580\,
            I => \DRA_c_7\
        );

    \I__1924\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8574\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__8574\,
            I => \N__8571\
        );

    \I__1922\ : Span4Mux_h
    port map (
            O => \N__8571\,
            I => \N__8568\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__8568\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1920\ : CEMux
    port map (
            O => \N__8565\,
            I => \N__8562\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__8562\,
            I => \N__8558\
        );

    \I__1918\ : CEMux
    port map (
            O => \N__8561\,
            I => \N__8554\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__8558\,
            I => \N__8551\
        );

    \I__1916\ : CEMux
    port map (
            O => \N__8557\,
            I => \N__8548\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__8554\,
            I => \N__8545\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__8551\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8548\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\
        );

    \I__1912\ : Odrv12
    port map (
            O => \N__8545\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\
        );

    \I__1911\ : InMux
    port map (
            O => \N__8538\,
            I => \N__8535\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__8535\,
            I => \N__8531\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8528\
        );

    \I__1908\ : Odrv12
    port map (
            O => \N__8531\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8528\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1906\ : InMux
    port map (
            O => \N__8523\,
            I => \N__8520\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8520\,
            I => \N__8516\
        );

    \I__1904\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8513\
        );

    \I__1903\ : Sp12to4
    port map (
            O => \N__8516\,
            I => \N__8509\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__8513\,
            I => \N__8506\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8503\
        );

    \I__1900\ : Span12Mux_v
    port map (
            O => \N__8509\,
            I => \N__8500\
        );

    \I__1899\ : Span4Mux_v
    port map (
            O => \N__8506\,
            I => \N__8497\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__8503\,
            I => \N__8494\
        );

    \I__1897\ : Odrv12
    port map (
            O => \N__8500\,
            I => \REG_CYCLEm\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__8497\,
            I => \REG_CYCLEm\
        );

    \I__1895\ : Odrv12
    port map (
            O => \N__8494\,
            I => \REG_CYCLEm\
        );

    \I__1894\ : IoInMux
    port map (
            O => \N__8487\,
            I => \N__8484\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__8484\,
            I => \N__8481\
        );

    \I__1892\ : IoSpan4Mux
    port map (
            O => \N__8481\,
            I => \N__8478\
        );

    \I__1891\ : IoSpan4Mux
    port map (
            O => \N__8478\,
            I => \N__8475\
        );

    \I__1890\ : Sp12to4
    port map (
            O => \N__8475\,
            I => \N__8472\
        );

    \I__1889\ : Span12Mux_s7_h
    port map (
            O => \N__8472\,
            I => \N__8469\
        );

    \I__1888\ : Odrv12
    port map (
            O => \N__8469\,
            I => \DRDENn_c\
        );

    \I__1887\ : InMux
    port map (
            O => \N__8466\,
            I => \N__8463\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__8463\,
            I => \N__8453\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__8462\,
            I => \N__8450\
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__8461\,
            I => \N__8447\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__8460\,
            I => \N__8444\
        );

    \I__1882\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8440\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__8458\,
            I => \N__8437\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__8457\,
            I => \N__8434\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__8456\,
            I => \N__8431\
        );

    \I__1878\ : Span4Mux_h
    port map (
            O => \N__8453\,
            I => \N__8427\
        );

    \I__1877\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8420\
        );

    \I__1876\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8420\
        );

    \I__1875\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8420\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8443\,
            I => \N__8417\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__8440\,
            I => \N__8414\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8411\
        );

    \I__1871\ : InMux
    port map (
            O => \N__8434\,
            I => \N__8408\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8431\,
            I => \N__8400\
        );

    \I__1869\ : CascadeMux
    port map (
            O => \N__8430\,
            I => \N__8393\
        );

    \I__1868\ : Span4Mux_v
    port map (
            O => \N__8427\,
            I => \N__8386\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8420\,
            I => \N__8386\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__8417\,
            I => \N__8386\
        );

    \I__1865\ : Span4Mux_h
    port map (
            O => \N__8414\,
            I => \N__8379\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8411\,
            I => \N__8379\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__8408\,
            I => \N__8379\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8407\,
            I => \N__8370\
        );

    \I__1861\ : InMux
    port map (
            O => \N__8406\,
            I => \N__8370\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8405\,
            I => \N__8370\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8370\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__8403\,
            I => \N__8365\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__8400\,
            I => \N__8361\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__8399\,
            I => \N__8357\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8398\,
            I => \N__8350\
        );

    \I__1854\ : InMux
    port map (
            O => \N__8397\,
            I => \N__8350\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8396\,
            I => \N__8350\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8347\
        );

    \I__1851\ : Span4Mux_h
    port map (
            O => \N__8386\,
            I => \N__8344\
        );

    \I__1850\ : Span4Mux_v
    port map (
            O => \N__8379\,
            I => \N__8339\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8370\,
            I => \N__8339\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8369\,
            I => \N__8336\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8368\,
            I => \N__8333\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8328\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8328\
        );

    \I__1844\ : Span4Mux_h
    port map (
            O => \N__8361\,
            I => \N__8325\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8320\
        );

    \I__1842\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8320\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8350\,
            I => \N__8317\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8347\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1839\ : Odrv4
    port map (
            O => \N__8344\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1838\ : Odrv4
    port map (
            O => \N__8339\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8336\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__8333\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8328\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__8325\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__8320\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1832\ : Odrv4
    port map (
            O => \N__8317\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1831\ : IoInMux
    port map (
            O => \N__8298\,
            I => \N__8295\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8295\,
            I => \N__8292\
        );

    \I__1829\ : Span4Mux_s0_v
    port map (
            O => \N__8292\,
            I => \N__8289\
        );

    \I__1828\ : Sp12to4
    port map (
            O => \N__8289\,
            I => \N__8286\
        );

    \I__1827\ : Span12Mux_h
    port map (
            O => \N__8286\,
            I => \N__8283\
        );

    \I__1826\ : Odrv12
    port map (
            O => \N__8283\,
            I => \CASn_c\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8276\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8273\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8276\,
            I => \N__8266\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8273\,
            I => \N__8263\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8272\,
            I => \N__8256\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8271\,
            I => \N__8256\
        );

    \I__1819\ : InMux
    port map (
            O => \N__8270\,
            I => \N__8256\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__8269\,
            I => \N__8252\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__8266\,
            I => \N__8249\
        );

    \I__1816\ : Span4Mux_v
    port map (
            O => \N__8263\,
            I => \N__8244\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8256\,
            I => \N__8244\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8255\,
            I => \N__8241\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8252\,
            I => \N__8238\
        );

    \I__1812\ : Odrv4
    port map (
            O => \N__8249\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__8244\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8241\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__8238\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1808\ : IoInMux
    port map (
            O => \N__8229\,
            I => \N__8226\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__8226\,
            I => \N__8223\
        );

    \I__1806\ : Span4Mux_s2_h
    port map (
            O => \N__8223\,
            I => \N__8220\
        );

    \I__1805\ : Sp12to4
    port map (
            O => \N__8220\,
            I => \N__8217\
        );

    \I__1804\ : Span12Mux_s7_v
    port map (
            O => \N__8217\,
            I => \N__8214\
        );

    \I__1803\ : Span12Mux_h
    port map (
            O => \N__8214\,
            I => \N__8211\
        );

    \I__1802\ : Odrv12
    port map (
            O => \N__8211\,
            I => \WEn_c\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8208\,
            I => \N__8202\
        );

    \I__1800\ : InMux
    port map (
            O => \N__8207\,
            I => \N__8199\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8196\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8193\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__8202\,
            I => \N__8184\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8199\,
            I => \N__8184\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__8196\,
            I => \N__8184\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__8193\,
            I => \N__8184\
        );

    \I__1793\ : Sp12to4
    port map (
            O => \N__8184\,
            I => \N__8181\
        );

    \I__1792\ : Span12Mux_v
    port map (
            O => \N__8181\,
            I => \N__8178\
        );

    \I__1791\ : Span12Mux_h
    port map (
            O => \N__8178\,
            I => \N__8175\
        );

    \I__1790\ : Odrv12
    port map (
            O => \N__8175\,
            I => \DRA_c_5\
        );

    \I__1789\ : InMux
    port map (
            O => \N__8172\,
            I => \N__8169\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8169\,
            I => \N__8163\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8168\,
            I => \N__8160\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8157\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8166\,
            I => \N__8154\
        );

    \I__1784\ : Span4Mux_h
    port map (
            O => \N__8163\,
            I => \N__8147\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8160\,
            I => \N__8147\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8157\,
            I => \N__8147\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__8154\,
            I => \N__8142\
        );

    \I__1780\ : Sp12to4
    port map (
            O => \N__8147\,
            I => \N__8142\
        );

    \I__1779\ : Span12Mux_v
    port map (
            O => \N__8142\,
            I => \N__8139\
        );

    \I__1778\ : Span12Mux_h
    port map (
            O => \N__8139\,
            I => \N__8136\
        );

    \I__1777\ : Odrv12
    port map (
            O => \N__8136\,
            I => \DRA_c_6\
        );

    \I__1776\ : InMux
    port map (
            O => \N__8133\,
            I => \N__8127\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8127\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__8127\,
            I => \N__8124\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__8124\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1772\ : InMux
    port map (
            O => \N__8121\,
            I => \N__8118\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__8118\,
            I => \N__8115\
        );

    \I__1770\ : Span4Mux_h
    port map (
            O => \N__8115\,
            I => \N__8112\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__8112\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__1768\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8106\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__8106\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8100\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8100\,
            I => \N__8097\
        );

    \I__1764\ : Odrv4
    port map (
            O => \N__8097\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1763\ : CascadeMux
    port map (
            O => \N__8094\,
            I => \N__8091\
        );

    \I__1762\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8088\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8088\,
            I => \N__8085\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__8085\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__1759\ : InMux
    port map (
            O => \N__8082\,
            I => \N__8078\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8081\,
            I => \N__8075\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8078\,
            I => \N__8072\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8075\,
            I => \N__8069\
        );

    \I__1755\ : Span4Mux_v
    port map (
            O => \N__8072\,
            I => \N__8066\
        );

    \I__1754\ : Span4Mux_h
    port map (
            O => \N__8069\,
            I => \N__8063\
        );

    \I__1753\ : Sp12to4
    port map (
            O => \N__8066\,
            I => \N__8060\
        );

    \I__1752\ : Sp12to4
    port map (
            O => \N__8063\,
            I => \N__8057\
        );

    \I__1751\ : Span12Mux_h
    port map (
            O => \N__8060\,
            I => \N__8054\
        );

    \I__1750\ : Span12Mux_v
    port map (
            O => \N__8057\,
            I => \N__8051\
        );

    \I__1749\ : Span12Mux_v
    port map (
            O => \N__8054\,
            I => \N__8048\
        );

    \I__1748\ : Span12Mux_h
    port map (
            O => \N__8051\,
            I => \N__8045\
        );

    \I__1747\ : Odrv12
    port map (
            O => \N__8048\,
            I => \DRA_c_0\
        );

    \I__1746\ : Odrv12
    port map (
            O => \N__8045\,
            I => \DRA_c_0\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8040\,
            I => \N__8037\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__8037\,
            I => \N__8034\
        );

    \I__1743\ : Span4Mux_h
    port map (
            O => \N__8034\,
            I => \N__8031\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__8031\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8028\,
            I => \N__8022\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8027\,
            I => \N__8022\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8022\,
            I => \N__8017\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8021\,
            I => \N__8012\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8020\,
            I => \N__8012\
        );

    \I__1736\ : Span4Mux_h
    port map (
            O => \N__8017\,
            I => \N__8007\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8012\,
            I => \N__8007\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__8007\,
            I => \N__8004\
        );

    \I__1733\ : Sp12to4
    port map (
            O => \N__8004\,
            I => \N__8001\
        );

    \I__1732\ : Span12Mux_v
    port map (
            O => \N__8001\,
            I => \N__7998\
        );

    \I__1731\ : Span12Mux_h
    port map (
            O => \N__7998\,
            I => \N__7995\
        );

    \I__1730\ : Odrv12
    port map (
            O => \N__7995\,
            I => \DRA_c_1\
        );

    \I__1729\ : InMux
    port map (
            O => \N__7992\,
            I => \N__7989\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__7986\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1726\ : InMux
    port map (
            O => \N__7983\,
            I => \N__7975\
        );

    \I__1725\ : InMux
    port map (
            O => \N__7982\,
            I => \N__7975\
        );

    \I__1724\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7970\
        );

    \I__1723\ : InMux
    port map (
            O => \N__7980\,
            I => \N__7970\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__7975\,
            I => \N__7965\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__7970\,
            I => \N__7965\
        );

    \I__1720\ : Sp12to4
    port map (
            O => \N__7965\,
            I => \N__7962\
        );

    \I__1719\ : Span12Mux_v
    port map (
            O => \N__7962\,
            I => \N__7959\
        );

    \I__1718\ : Span12Mux_h
    port map (
            O => \N__7959\,
            I => \N__7956\
        );

    \I__1717\ : Odrv12
    port map (
            O => \N__7956\,
            I => \DRA_c_2\
        );

    \I__1716\ : InMux
    port map (
            O => \N__7953\,
            I => \N__7950\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__7950\,
            I => \N__7947\
        );

    \I__1714\ : Span4Mux_h
    port map (
            O => \N__7947\,
            I => \N__7944\
        );

    \I__1713\ : Odrv4
    port map (
            O => \N__7944\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1712\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7938\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__7938\,
            I => \N__7935\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__7935\,
            I => \N__7932\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__7932\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1708\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7926\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__7926\,
            I => \N__7923\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__7923\,
            I => \N__7920\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__7920\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__7917\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10_cascade_\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__7914\,
            I => \N__7909\
        );

    \I__1702\ : InMux
    port map (
            O => \N__7913\,
            I => \N__7905\
        );

    \I__1701\ : InMux
    port map (
            O => \N__7912\,
            I => \N__7898\
        );

    \I__1700\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7898\
        );

    \I__1699\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7898\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__7905\,
            I => \N__7895\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__7898\,
            I => \N__7892\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__7895\,
            I => \N__7889\
        );

    \I__1695\ : Span4Mux_v
    port map (
            O => \N__7892\,
            I => \N__7886\
        );

    \I__1694\ : Span4Mux_v
    port map (
            O => \N__7889\,
            I => \N__7881\
        );

    \I__1693\ : Span4Mux_h
    port map (
            O => \N__7886\,
            I => \N__7881\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__7881\,
            I => \N__7878\
        );

    \I__1691\ : Span4Mux_v
    port map (
            O => \N__7878\,
            I => \N__7875\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__7875\,
            I => \CLK40_PLL_i\
        );

    \I__1689\ : IoInMux
    port map (
            O => \N__7872\,
            I => \N__7867\
        );

    \I__1688\ : IoInMux
    port map (
            O => \N__7871\,
            I => \N__7864\
        );

    \I__1687\ : IoInMux
    port map (
            O => \N__7870\,
            I => \N__7861\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__7867\,
            I => \N__7858\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__7864\,
            I => \N__7855\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__7861\,
            I => \N__7852\
        );

    \I__1683\ : Span4Mux_s3_v
    port map (
            O => \N__7858\,
            I => \N__7849\
        );

    \I__1682\ : Span4Mux_s3_h
    port map (
            O => \N__7855\,
            I => \N__7846\
        );

    \I__1681\ : Span12Mux_s3_v
    port map (
            O => \N__7852\,
            I => \N__7843\
        );

    \I__1680\ : Sp12to4
    port map (
            O => \N__7849\,
            I => \N__7840\
        );

    \I__1679\ : Span4Mux_h
    port map (
            O => \N__7846\,
            I => \N__7837\
        );

    \I__1678\ : Span12Mux_v
    port map (
            O => \N__7843\,
            I => \N__7834\
        );

    \I__1677\ : Span12Mux_h
    port map (
            O => \N__7840\,
            I => \N__7831\
        );

    \I__1676\ : Span4Mux_h
    port map (
            O => \N__7837\,
            I => \N__7828\
        );

    \I__1675\ : Span12Mux_h
    port map (
            O => \N__7834\,
            I => \N__7825\
        );

    \I__1674\ : Span12Mux_v
    port map (
            O => \N__7831\,
            I => \N__7822\
        );

    \I__1673\ : Span4Mux_h
    port map (
            O => \N__7828\,
            I => \N__7819\
        );

    \I__1672\ : Odrv12
    port map (
            O => \N__7825\,
            I => \CLK40_PLL_i_i\
        );

    \I__1671\ : Odrv12
    port map (
            O => \N__7822\,
            I => \CLK40_PLL_i_i\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__7819\,
            I => \CLK40_PLL_i_i\
        );

    \I__1669\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7808\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7805\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__7808\,
            I => \N__7801\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__7805\,
            I => \N__7798\
        );

    \I__1665\ : InMux
    port map (
            O => \N__7804\,
            I => \N__7795\
        );

    \I__1664\ : Span4Mux_h
    port map (
            O => \N__7801\,
            I => \N__7790\
        );

    \I__1663\ : Span4Mux_v
    port map (
            O => \N__7798\,
            I => \N__7790\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7795\,
            I => \N__7786\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__7790\,
            I => \N__7783\
        );

    \I__1660\ : InMux
    port map (
            O => \N__7789\,
            I => \N__7780\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__7786\,
            I => \N__7777\
        );

    \I__1658\ : Span4Mux_v
    port map (
            O => \N__7783\,
            I => \N__7772\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__7780\,
            I => \N__7772\
        );

    \I__1656\ : Sp12to4
    port map (
            O => \N__7777\,
            I => \N__7769\
        );

    \I__1655\ : Span4Mux_h
    port map (
            O => \N__7772\,
            I => \N__7766\
        );

    \I__1654\ : Span12Mux_h
    port map (
            O => \N__7769\,
            I => \N__7763\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__7766\,
            I => \N__7760\
        );

    \I__1652\ : Span12Mux_v
    port map (
            O => \N__7763\,
            I => \N__7757\
        );

    \I__1651\ : Span4Mux_h
    port map (
            O => \N__7760\,
            I => \N__7754\
        );

    \I__1650\ : Odrv12
    port map (
            O => \N__7757\,
            I => \DBRn_c\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__7754\,
            I => \DBRn_c\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7749\,
            I => \N__7743\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7748\,
            I => \N__7740\
        );

    \I__1646\ : InMux
    port map (
            O => \N__7747\,
            I => \N__7735\
        );

    \I__1645\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7735\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7743\,
            I => \N__7727\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7740\,
            I => \N__7724\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__7735\,
            I => \N__7721\
        );

    \I__1641\ : ClkMux
    port map (
            O => \N__7734\,
            I => \N__7704\
        );

    \I__1640\ : ClkMux
    port map (
            O => \N__7733\,
            I => \N__7704\
        );

    \I__1639\ : ClkMux
    port map (
            O => \N__7732\,
            I => \N__7704\
        );

    \I__1638\ : ClkMux
    port map (
            O => \N__7731\,
            I => \N__7704\
        );

    \I__1637\ : ClkMux
    port map (
            O => \N__7730\,
            I => \N__7704\
        );

    \I__1636\ : Glb2LocalMux
    port map (
            O => \N__7727\,
            I => \N__7704\
        );

    \I__1635\ : Glb2LocalMux
    port map (
            O => \N__7724\,
            I => \N__7704\
        );

    \I__1634\ : Glb2LocalMux
    port map (
            O => \N__7721\,
            I => \N__7704\
        );

    \I__1633\ : GlobalMux
    port map (
            O => \N__7704\,
            I => \N__7701\
        );

    \I__1632\ : gio2CtrlBuf
    port map (
            O => \N__7701\,
            I => \C1_c_g\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7698\,
            I => \N__7689\
        );

    \I__1630\ : InMux
    port map (
            O => \N__7697\,
            I => \N__7686\
        );

    \I__1629\ : InMux
    port map (
            O => \N__7696\,
            I => \N__7682\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7695\,
            I => \N__7677\
        );

    \I__1627\ : InMux
    port map (
            O => \N__7694\,
            I => \N__7677\
        );

    \I__1626\ : InMux
    port map (
            O => \N__7693\,
            I => \N__7672\
        );

    \I__1625\ : InMux
    port map (
            O => \N__7692\,
            I => \N__7672\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7689\,
            I => \N__7667\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__7686\,
            I => \N__7667\
        );

    \I__1622\ : InMux
    port map (
            O => \N__7685\,
            I => \N__7664\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__7682\,
            I => \N__7658\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__7677\,
            I => \N__7654\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7672\,
            I => \N__7647\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__7667\,
            I => \N__7647\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__7664\,
            I => \N__7647\
        );

    \I__1616\ : InMux
    port map (
            O => \N__7663\,
            I => \N__7644\
        );

    \I__1615\ : InMux
    port map (
            O => \N__7662\,
            I => \N__7641\
        );

    \I__1614\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7638\
        );

    \I__1613\ : Span4Mux_h
    port map (
            O => \N__7658\,
            I => \N__7635\
        );

    \I__1612\ : InMux
    port map (
            O => \N__7657\,
            I => \N__7632\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__7654\,
            I => \N__7629\
        );

    \I__1610\ : Span4Mux_h
    port map (
            O => \N__7647\,
            I => \N__7624\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__7644\,
            I => \N__7624\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__7641\,
            I => \N__7621\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__7638\,
            I => \N__7618\
        );

    \I__1606\ : Sp12to4
    port map (
            O => \N__7635\,
            I => \N__7607\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__7632\,
            I => \N__7607\
        );

    \I__1604\ : Span4Mux_v
    port map (
            O => \N__7629\,
            I => \N__7602\
        );

    \I__1603\ : Span4Mux_v
    port map (
            O => \N__7624\,
            I => \N__7602\
        );

    \I__1602\ : Span4Mux_v
    port map (
            O => \N__7621\,
            I => \N__7597\
        );

    \I__1601\ : Span4Mux_v
    port map (
            O => \N__7618\,
            I => \N__7597\
        );

    \I__1600\ : InMux
    port map (
            O => \N__7617\,
            I => \N__7588\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7616\,
            I => \N__7588\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7615\,
            I => \N__7588\
        );

    \I__1597\ : InMux
    port map (
            O => \N__7614\,
            I => \N__7588\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7613\,
            I => \N__7583\
        );

    \I__1595\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7583\
        );

    \I__1594\ : Span12Mux_v
    port map (
            O => \N__7607\,
            I => \N__7578\
        );

    \I__1593\ : Sp12to4
    port map (
            O => \N__7602\,
            I => \N__7578\
        );

    \I__1592\ : Sp12to4
    port map (
            O => \N__7597\,
            I => \N__7571\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__7588\,
            I => \N__7571\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__7583\,
            I => \N__7571\
        );

    \I__1589\ : Span12Mux_h
    port map (
            O => \N__7578\,
            I => \N__7568\
        );

    \I__1588\ : Span12Mux_h
    port map (
            O => \N__7571\,
            I => \N__7565\
        );

    \I__1587\ : Odrv12
    port map (
            O => \N__7568\,
            I => \RESETn_c\
        );

    \I__1586\ : Odrv12
    port map (
            O => \N__7565\,
            I => \RESETn_c\
        );

    \I__1585\ : IoInMux
    port map (
            O => \N__7560\,
            I => \N__7557\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7557\,
            I => \N__7554\
        );

    \I__1583\ : Odrv12
    port map (
            O => \N__7554\,
            I => \RESETn_c_i\
        );

    \I__1582\ : InMux
    port map (
            O => \N__7551\,
            I => \N__7547\
        );

    \I__1581\ : InMux
    port map (
            O => \N__7550\,
            I => \N__7544\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__7547\,
            I => \N__7541\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7544\,
            I => \N__7537\
        );

    \I__1578\ : Span4Mux_h
    port map (
            O => \N__7541\,
            I => \N__7534\
        );

    \I__1577\ : InMux
    port map (
            O => \N__7540\,
            I => \N__7527\
        );

    \I__1576\ : Span4Mux_v
    port map (
            O => \N__7537\,
            I => \N__7522\
        );

    \I__1575\ : Span4Mux_v
    port map (
            O => \N__7534\,
            I => \N__7522\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7533\,
            I => \N__7517\
        );

    \I__1573\ : InMux
    port map (
            O => \N__7532\,
            I => \N__7517\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7531\,
            I => \N__7514\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7530\,
            I => \N__7511\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7527\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1569\ : Odrv4
    port map (
            O => \N__7522\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7517\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__7514\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7511\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1565\ : IoInMux
    port map (
            O => \N__7500\,
            I => \N__7497\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__7497\,
            I => \N__7494\
        );

    \I__1563\ : IoSpan4Mux
    port map (
            O => \N__7494\,
            I => \N__7491\
        );

    \I__1562\ : Sp12to4
    port map (
            O => \N__7491\,
            I => \N__7488\
        );

    \I__1561\ : Span12Mux_s7_v
    port map (
            O => \N__7488\,
            I => \N__7485\
        );

    \I__1560\ : Odrv12
    port map (
            O => \N__7485\,
            I => \RASn_c\
        );

    \I__1559\ : InMux
    port map (
            O => \N__7482\,
            I => \N__7478\
        );

    \I__1558\ : InMux
    port map (
            O => \N__7481\,
            I => \N__7475\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7478\,
            I => \N__7472\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7475\,
            I => \N__7469\
        );

    \I__1555\ : Span4Mux_v
    port map (
            O => \N__7472\,
            I => \N__7464\
        );

    \I__1554\ : Span4Mux_v
    port map (
            O => \N__7469\,
            I => \N__7461\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7456\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7467\,
            I => \N__7456\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__7464\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1550\ : Odrv4
    port map (
            O => \N__7461\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7456\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7449\,
            I => \N__7446\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7446\,
            I => \N__7443\
        );

    \I__1546\ : Span4Mux_v
    port map (
            O => \N__7443\,
            I => \N__7440\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__7440\,
            I => \N__7437\
        );

    \I__1544\ : Sp12to4
    port map (
            O => \N__7437\,
            I => \N__7434\
        );

    \I__1543\ : Span12Mux_h
    port map (
            O => \N__7434\,
            I => \N__7431\
        );

    \I__1542\ : Odrv12
    port map (
            O => \N__7431\,
            I => \A_c_19\
        );

    \I__1541\ : IoInMux
    port map (
            O => \N__7428\,
            I => \N__7425\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7425\,
            I => \N__7422\
        );

    \I__1539\ : IoSpan4Mux
    port map (
            O => \N__7422\,
            I => \N__7419\
        );

    \I__1538\ : IoSpan4Mux
    port map (
            O => \N__7419\,
            I => \N__7416\
        );

    \I__1537\ : Span4Mux_s2_h
    port map (
            O => \N__7416\,
            I => \N__7413\
        );

    \I__1536\ : Sp12to4
    port map (
            O => \N__7413\,
            I => \N__7410\
        );

    \I__1535\ : Odrv12
    port map (
            O => \N__7410\,
            I => \CMA_c_9\
        );

    \I__1534\ : CEMux
    port map (
            O => \N__7407\,
            I => \N__7404\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7404\,
            I => \N__7400\
        );

    \I__1532\ : CEMux
    port map (
            O => \N__7403\,
            I => \N__7397\
        );

    \I__1531\ : Span4Mux_v
    port map (
            O => \N__7400\,
            I => \N__7391\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7397\,
            I => \N__7391\
        );

    \I__1529\ : CEMux
    port map (
            O => \N__7396\,
            I => \N__7388\
        );

    \I__1528\ : Span4Mux_v
    port map (
            O => \N__7391\,
            I => \N__7382\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7388\,
            I => \N__7379\
        );

    \I__1526\ : CEMux
    port map (
            O => \N__7387\,
            I => \N__7376\
        );

    \I__1525\ : CEMux
    port map (
            O => \N__7386\,
            I => \N__7373\
        );

    \I__1524\ : CEMux
    port map (
            O => \N__7385\,
            I => \N__7370\
        );

    \I__1523\ : Odrv4
    port map (
            O => \N__7382\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1522\ : Odrv12
    port map (
            O => \N__7379\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7376\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7373\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7370\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__7359\,
            I => \N__7353\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__7358\,
            I => \N__7350\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__7357\,
            I => \N__7343\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__7356\,
            I => \N__7340\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7353\,
            I => \N__7337\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7350\,
            I => \N__7333\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7349\,
            I => \N__7330\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7348\,
            I => \N__7327\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7347\,
            I => \N__7322\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7346\,
            I => \N__7322\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7343\,
            I => \N__7317\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7340\,
            I => \N__7317\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7337\,
            I => \N__7314\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7311\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7333\,
            I => \N__7306\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7330\,
            I => \N__7306\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7327\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7322\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7317\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__7314\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7311\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1497\ : Odrv12
    port map (
            O => \N__7306\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7290\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7290\,
            I => \N__7287\
        );

    \I__1494\ : Odrv4
    port map (
            O => \N__7287\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1493\ : InMux
    port map (
            O => \N__7284\,
            I => \N__7281\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7281\,
            I => \N__7278\
        );

    \I__1491\ : Odrv4
    port map (
            O => \N__7278\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7275\,
            I => \N__7272\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7272\,
            I => \N__7269\
        );

    \I__1488\ : Span4Mux_v
    port map (
            O => \N__7269\,
            I => \N__7266\
        );

    \I__1487\ : Span4Mux_h
    port map (
            O => \N__7266\,
            I => \N__7262\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7265\,
            I => \N__7259\
        );

    \I__1485\ : Odrv4
    port map (
            O => \N__7262\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7259\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7254\,
            I => \N__7251\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7251\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7248\,
            I => \N__7245\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7245\,
            I => \N__7242\
        );

    \I__1479\ : Odrv12
    port map (
            O => \N__7242\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7239\,
            I => \N__7236\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__7236\,
            I => \N__7233\
        );

    \I__1476\ : Span4Mux_h
    port map (
            O => \N__7233\,
            I => \N__7230\
        );

    \I__1475\ : Odrv4
    port map (
            O => \N__7230\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__1474\ : CascadeMux
    port map (
            O => \N__7227\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_\
        );

    \I__1473\ : IoInMux
    port map (
            O => \N__7224\,
            I => \N__7221\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7221\,
            I => \N__7218\
        );

    \I__1471\ : Span12Mux_s4_h
    port map (
            O => \N__7218\,
            I => \N__7215\
        );

    \I__1470\ : Span12Mux_h
    port map (
            O => \N__7215\,
            I => \N__7212\
        );

    \I__1469\ : Odrv12
    port map (
            O => \N__7212\,
            I => \CMA_c_4\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__7209\,
            I => \N__7206\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7206\,
            I => \N__7196\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7205\,
            I => \N__7196\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7204\,
            I => \N__7196\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7203\,
            I => \N__7193\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7196\,
            I => \N__7188\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7193\,
            I => \N__7185\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7180\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7191\,
            I => \N__7180\
        );

    \I__1459\ : Odrv4
    port map (
            O => \N__7188\,
            I => \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5Z0Z_1\
        );

    \I__1458\ : Odrv4
    port map (
            O => \N__7185\,
            I => \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5Z0Z_1\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7180\,
            I => \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5Z0Z_1\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7170\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7170\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1454\ : IoInMux
    port map (
            O => \N__7167\,
            I => \N__7164\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7164\,
            I => \N__7161\
        );

    \I__1452\ : Span4Mux_s2_h
    port map (
            O => \N__7161\,
            I => \N__7158\
        );

    \I__1451\ : Sp12to4
    port map (
            O => \N__7158\,
            I => \N__7155\
        );

    \I__1450\ : Span12Mux_v
    port map (
            O => \N__7155\,
            I => \N__7152\
        );

    \I__1449\ : Span12Mux_h
    port map (
            O => \N__7152\,
            I => \N__7149\
        );

    \I__1448\ : Odrv12
    port map (
            O => \N__7149\,
            I => \CMA_c_7\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7146\,
            I => \N__7143\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7143\,
            I => \N__7140\
        );

    \I__1445\ : Odrv4
    port map (
            O => \N__7140\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7137\,
            I => \N__7134\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7134\,
            I => \N__7130\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7133\,
            I => \N__7127\
        );

    \I__1441\ : Span4Mux_h
    port map (
            O => \N__7130\,
            I => \N__7124\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__7127\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__1439\ : Odrv4
    port map (
            O => \N__7124\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7119\,
            I => \N__7116\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7116\,
            I => \N__7113\
        );

    \I__1436\ : Span4Mux_v
    port map (
            O => \N__7113\,
            I => \N__7110\
        );

    \I__1435\ : Span4Mux_h
    port map (
            O => \N__7110\,
            I => \N__7107\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__7107\,
            I => \U712_CHIP_RAM.un5_DMA_CYCLE_START_0\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7104\,
            I => \N__7101\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7101\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7098\,
            I => \N__7094\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7097\,
            I => \N__7091\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7094\,
            I => \U712_REG_SM.ASn_0_sqmuxa_1\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__7091\,
            I => \U712_REG_SM.ASn_0_sqmuxa_1\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7086\,
            I => \N__7082\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7085\,
            I => \N__7079\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7082\,
            I => \U712_REG_SM.N_226\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7079\,
            I => \U712_REG_SM.N_226\
        );

    \I__1423\ : IoInMux
    port map (
            O => \N__7074\,
            I => \N__7071\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7071\,
            I => \N__7068\
        );

    \I__1421\ : IoSpan4Mux
    port map (
            O => \N__7068\,
            I => \N__7065\
        );

    \I__1420\ : Span4Mux_s1_v
    port map (
            O => \N__7065\,
            I => \N__7062\
        );

    \I__1419\ : Span4Mux_v
    port map (
            O => \N__7062\,
            I => \N__7059\
        );

    \I__1418\ : Sp12to4
    port map (
            O => \N__7059\,
            I => \N__7056\
        );

    \I__1417\ : Span12Mux_h
    port map (
            O => \N__7056\,
            I => \N__7052\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7055\,
            I => \N__7049\
        );

    \I__1415\ : Odrv12
    port map (
            O => \N__7052\,
            I => \ASn_c\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__7049\,
            I => \ASn_c\
        );

    \I__1413\ : IoInMux
    port map (
            O => \N__7044\,
            I => \N__7041\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7041\,
            I => \N__7038\
        );

    \I__1411\ : Span4Mux_s2_v
    port map (
            O => \N__7038\,
            I => \N__7035\
        );

    \I__1410\ : Span4Mux_v
    port map (
            O => \N__7035\,
            I => \N__7032\
        );

    \I__1409\ : Odrv4
    port map (
            O => \N__7032\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1408\ : IoInMux
    port map (
            O => \N__7029\,
            I => \N__7026\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7026\,
            I => \N__7023\
        );

    \I__1406\ : Span12Mux_s8_v
    port map (
            O => \N__7023\,
            I => \N__7020\
        );

    \I__1405\ : Odrv12
    port map (
            O => \N__7020\,
            I => \CMA_c_10\
        );

    \I__1404\ : IoInMux
    port map (
            O => \N__7017\,
            I => \N__7014\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7014\,
            I => \N__7011\
        );

    \I__1402\ : IoSpan4Mux
    port map (
            O => \N__7011\,
            I => \N__7008\
        );

    \I__1401\ : Span4Mux_s2_v
    port map (
            O => \N__7008\,
            I => \N__7005\
        );

    \I__1400\ : Span4Mux_v
    port map (
            O => \N__7005\,
            I => \N__7002\
        );

    \I__1399\ : Span4Mux_v
    port map (
            O => \N__7002\,
            I => \N__6999\
        );

    \I__1398\ : Odrv4
    port map (
            O => \N__6999\,
            I => \CMA_c_0\
        );

    \I__1397\ : InMux
    port map (
            O => \N__6996\,
            I => \N__6993\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__6993\,
            I => \N__6990\
        );

    \I__1395\ : Span12Mux_v
    port map (
            O => \N__6990\,
            I => \N__6987\
        );

    \I__1394\ : Span12Mux_h
    port map (
            O => \N__6987\,
            I => \N__6984\
        );

    \I__1393\ : Odrv12
    port map (
            O => \N__6984\,
            I => \A_c_17\
        );

    \I__1392\ : IoInMux
    port map (
            O => \N__6981\,
            I => \N__6978\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6978\,
            I => \N__6975\
        );

    \I__1390\ : IoSpan4Mux
    port map (
            O => \N__6975\,
            I => \N__6972\
        );

    \I__1389\ : Span4Mux_s2_h
    port map (
            O => \N__6972\,
            I => \N__6969\
        );

    \I__1388\ : Sp12to4
    port map (
            O => \N__6969\,
            I => \N__6966\
        );

    \I__1387\ : Span12Mux_h
    port map (
            O => \N__6966\,
            I => \N__6963\
        );

    \I__1386\ : Odrv12
    port map (
            O => \N__6963\,
            I => \CMA_c_8\
        );

    \I__1385\ : InMux
    port map (
            O => \N__6960\,
            I => \N__6957\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__6957\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1383\ : IoInMux
    port map (
            O => \N__6954\,
            I => \N__6951\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__6951\,
            I => \N__6948\
        );

    \I__1381\ : IoSpan4Mux
    port map (
            O => \N__6948\,
            I => \N__6945\
        );

    \I__1380\ : Span4Mux_s3_h
    port map (
            O => \N__6945\,
            I => \N__6942\
        );

    \I__1379\ : Span4Mux_h
    port map (
            O => \N__6942\,
            I => \N__6939\
        );

    \I__1378\ : Sp12to4
    port map (
            O => \N__6939\,
            I => \N__6936\
        );

    \I__1377\ : Span12Mux_h
    port map (
            O => \N__6936\,
            I => \N__6933\
        );

    \I__1376\ : Odrv12
    port map (
            O => \N__6933\,
            I => \CMA_c_3\
        );

    \I__1375\ : IoInMux
    port map (
            O => \N__6930\,
            I => \N__6927\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__6927\,
            I => \N__6924\
        );

    \I__1373\ : IoSpan4Mux
    port map (
            O => \N__6924\,
            I => \N__6921\
        );

    \I__1372\ : Span4Mux_s3_h
    port map (
            O => \N__6921\,
            I => \N__6918\
        );

    \I__1371\ : Span4Mux_v
    port map (
            O => \N__6918\,
            I => \N__6915\
        );

    \I__1370\ : Span4Mux_h
    port map (
            O => \N__6915\,
            I => \N__6912\
        );

    \I__1369\ : Sp12to4
    port map (
            O => \N__6912\,
            I => \N__6909\
        );

    \I__1368\ : Odrv12
    port map (
            O => \N__6909\,
            I => \CMA_c_6\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6906\,
            I => \N__6903\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__6903\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6897\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__6897\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6894\,
            I => \N__6891\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__6891\,
            I => \N__6888\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__6888\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1360\ : InMux
    port map (
            O => \N__6885\,
            I => \N__6882\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__6882\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1358\ : IoInMux
    port map (
            O => \N__6879\,
            I => \N__6876\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__6876\,
            I => \N__6873\
        );

    \I__1356\ : IoSpan4Mux
    port map (
            O => \N__6873\,
            I => \N__6870\
        );

    \I__1355\ : Span4Mux_s3_h
    port map (
            O => \N__6870\,
            I => \N__6867\
        );

    \I__1354\ : Sp12to4
    port map (
            O => \N__6867\,
            I => \N__6864\
        );

    \I__1353\ : Span12Mux_h
    port map (
            O => \N__6864\,
            I => \N__6861\
        );

    \I__1352\ : Odrv12
    port map (
            O => \N__6861\,
            I => \CMA_c_5\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6858\,
            I => \N__6855\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6855\,
            I => \N__6852\
        );

    \I__1349\ : Span4Mux_v
    port map (
            O => \N__6852\,
            I => \N__6849\
        );

    \I__1348\ : Sp12to4
    port map (
            O => \N__6849\,
            I => \N__6846\
        );

    \I__1347\ : Span12Mux_h
    port map (
            O => \N__6846\,
            I => \N__6843\
        );

    \I__1346\ : Odrv12
    port map (
            O => \N__6843\,
            I => \A_c_9\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6840\,
            I => \N__6837\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__6837\,
            I => \N__6834\
        );

    \I__1343\ : Span4Mux_v
    port map (
            O => \N__6834\,
            I => \N__6831\
        );

    \I__1342\ : Sp12to4
    port map (
            O => \N__6831\,
            I => \N__6828\
        );

    \I__1341\ : Span12Mux_v
    port map (
            O => \N__6828\,
            I => \N__6825\
        );

    \I__1340\ : Span12Mux_h
    port map (
            O => \N__6825\,
            I => \N__6822\
        );

    \I__1339\ : Odrv12
    port map (
            O => \N__6822\,
            I => \A_c_2\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6819\,
            I => \N__6816\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6816\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6813\,
            I => \N__6810\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__6810\,
            I => \N__6807\
        );

    \I__1334\ : Span4Mux_v
    port map (
            O => \N__6807\,
            I => \N__6804\
        );

    \I__1333\ : Sp12to4
    port map (
            O => \N__6804\,
            I => \N__6801\
        );

    \I__1332\ : Span12Mux_h
    port map (
            O => \N__6801\,
            I => \N__6798\
        );

    \I__1331\ : Odrv12
    port map (
            O => \N__6798\,
            I => \A_c_10\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6795\,
            I => \N__6792\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6792\,
            I => \N__6789\
        );

    \I__1328\ : Span12Mux_h
    port map (
            O => \N__6789\,
            I => \N__6786\
        );

    \I__1327\ : Span12Mux_v
    port map (
            O => \N__6786\,
            I => \N__6783\
        );

    \I__1326\ : Odrv12
    port map (
            O => \N__6783\,
            I => \A_c_3\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__6780\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\
        );

    \I__1324\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6774\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__6774\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__6771\,
            I => \N__6768\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6762\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6767\,
            I => \N__6762\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6762\,
            I => \N__6759\
        );

    \I__1318\ : Span4Mux_v
    port map (
            O => \N__6759\,
            I => \N__6756\
        );

    \I__1317\ : Span4Mux_v
    port map (
            O => \N__6756\,
            I => \N__6753\
        );

    \I__1316\ : Sp12to4
    port map (
            O => \N__6753\,
            I => \N__6750\
        );

    \I__1315\ : Span12Mux_h
    port map (
            O => \N__6750\,
            I => \N__6747\
        );

    \I__1314\ : Odrv12
    port map (
            O => \N__6747\,
            I => \A_c_14\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6741\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6741\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1311\ : InMux
    port map (
            O => \N__6738\,
            I => \N__6733\
        );

    \I__1310\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6728\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6728\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__6733\,
            I => \N__6725\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__6728\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1306\ : Odrv4
    port map (
            O => \N__6725\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6716\
        );

    \I__1304\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6713\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6716\,
            I => \N__6710\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__6713\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1301\ : Odrv12
    port map (
            O => \N__6710\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6705\,
            I => \N__6702\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6702\,
            I => \N__6699\
        );

    \I__1298\ : Odrv12
    port map (
            O => \N__6699\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6696\,
            I => \N__6687\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6695\,
            I => \N__6680\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6694\,
            I => \N__6680\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6693\,
            I => \N__6680\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6692\,
            I => \N__6677\
        );

    \I__1292\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6672\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6690\,
            I => \N__6672\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__6687\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6680\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6677\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__6672\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__6663\,
            I => \N__6659\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__6662\,
            I => \N__6654\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6659\,
            I => \N__6648\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6658\,
            I => \N__6648\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6657\,
            I => \N__6645\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6654\,
            I => \N__6642\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6639\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6648\,
            I => \N__6636\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__6645\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6642\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__6639\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__6636\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__1274\ : CascadeMux
    port map (
            O => \N__6627\,
            I => \N__6619\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__6626\,
            I => \N__6616\
        );

    \I__1272\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6613\
        );

    \I__1271\ : InMux
    port map (
            O => \N__6624\,
            I => \N__6608\
        );

    \I__1270\ : InMux
    port map (
            O => \N__6623\,
            I => \N__6608\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6622\,
            I => \N__6605\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6600\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6616\,
            I => \N__6600\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__6613\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6608\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6605\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__6600\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6591\,
            I => \N__6581\
        );

    \I__1261\ : InMux
    port map (
            O => \N__6590\,
            I => \N__6576\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6589\,
            I => \N__6576\
        );

    \I__1259\ : InMux
    port map (
            O => \N__6588\,
            I => \N__6573\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6587\,
            I => \N__6564\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6564\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6585\,
            I => \N__6564\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6584\,
            I => \N__6564\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6581\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__6576\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6573\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__6564\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__6555\,
            I => \N__6551\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6544\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6541\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6536\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6536\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6548\,
            I => \N__6531\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6531\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__6544\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6541\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6536\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__6531\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6519\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6519\,
            I => \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__6516\,
            I => \N__6513\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6513\,
            I => \N__6510\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6510\,
            I => \N__6507\
        );

    \I__1234\ : Odrv4
    port map (
            O => \N__6507\,
            I => \U712_REG_SM.DS_EN_RNOZ0Z_0\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6504\,
            I => \N__6501\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6501\,
            I => \U712_REG_SM.N_300\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6494\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6497\,
            I => \N__6491\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__6494\,
            I => \U712_REG_SM.N_228\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__6491\,
            I => \U712_REG_SM.N_228\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6486\,
            I => \N__6483\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6483\,
            I => \N__6480\
        );

    \I__1225\ : Span4Mux_h
    port map (
            O => \N__6480\,
            I => \N__6476\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6473\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__6476\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__6473\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__1221\ : IoInMux
    port map (
            O => \N__6468\,
            I => \N__6465\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6465\,
            I => \N__6461\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6457\
        );

    \I__1218\ : Span12Mux_s2_v
    port map (
            O => \N__6461\,
            I => \N__6454\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__6460\,
            I => \N__6451\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__6457\,
            I => \N__6448\
        );

    \I__1215\ : Span12Mux_v
    port map (
            O => \N__6454\,
            I => \N__6445\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6451\,
            I => \N__6442\
        );

    \I__1213\ : Span4Mux_v
    port map (
            O => \N__6448\,
            I => \N__6439\
        );

    \I__1212\ : Odrv12
    port map (
            O => \N__6445\,
            I => \REGENn_c\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6442\,
            I => \REGENn_c\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__6439\,
            I => \REGENn_c\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6432\,
            I => \N__6429\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6429\,
            I => \N__6426\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__6426\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1206\ : IoInMux
    port map (
            O => \N__6423\,
            I => \N__6420\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6420\,
            I => \N__6417\
        );

    \I__1204\ : Span12Mux_s9_v
    port map (
            O => \N__6417\,
            I => \N__6414\
        );

    \I__1203\ : Odrv12
    port map (
            O => \N__6414\,
            I => \CMA_c_2\
        );

    \I__1202\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6408\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6408\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6405\,
            I => \N__6402\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6402\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6399\,
            I => \N__6396\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6396\,
            I => \N__6393\
        );

    \I__1196\ : Span4Mux_h
    port map (
            O => \N__6393\,
            I => \N__6390\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__6390\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1194\ : IoInMux
    port map (
            O => \N__6387\,
            I => \N__6384\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6384\,
            I => \N__6381\
        );

    \I__1192\ : Span4Mux_s3_v
    port map (
            O => \N__6381\,
            I => \N__6378\
        );

    \I__1191\ : Span4Mux_v
    port map (
            O => \N__6378\,
            I => \N__6375\
        );

    \I__1190\ : Odrv4
    port map (
            O => \N__6375\,
            I => \CMA_c_1\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6359\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6359\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6370\,
            I => \N__6359\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6369\,
            I => \N__6356\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6349\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6349\
        );

    \I__1183\ : InMux
    port map (
            O => \N__6366\,
            I => \N__6349\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6359\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6356\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6349\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6342\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6339\,
            I => \N__6335\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6338\,
            I => \N__6332\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6335\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6332\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1174\ : CEMux
    port map (
            O => \N__6327\,
            I => \N__6324\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__6324\,
            I => \N__6320\
        );

    \I__1172\ : CEMux
    port map (
            O => \N__6323\,
            I => \N__6317\
        );

    \I__1171\ : Span4Mux_v
    port map (
            O => \N__6320\,
            I => \N__6314\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6317\,
            I => \N__6311\
        );

    \I__1169\ : Span4Mux_h
    port map (
            O => \N__6314\,
            I => \N__6306\
        );

    \I__1168\ : Span4Mux_v
    port map (
            O => \N__6311\,
            I => \N__6306\
        );

    \I__1167\ : Span4Mux_h
    port map (
            O => \N__6306\,
            I => \N__6303\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__6303\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__1165\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6297\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6297\,
            I => \N__6294\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__6294\,
            I => \U712_CHIP_RAM.N_285\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6285\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6290\,
            I => \N__6282\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6289\,
            I => \N__6277\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6288\,
            I => \N__6277\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6285\,
            I => \N__6271\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6282\,
            I => \N__6271\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6277\,
            I => \N__6268\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6276\,
            I => \N__6265\
        );

    \I__1154\ : Odrv4
    port map (
            O => \N__6271\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__6268\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6265\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__6258\,
            I => \N__6253\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6257\,
            I => \N__6243\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6256\,
            I => \N__6243\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6253\,
            I => \N__6243\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__6252\,
            I => \N__6238\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6251\,
            I => \N__6233\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6250\,
            I => \N__6233\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__6243\,
            I => \N__6230\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__6242\,
            I => \N__6227\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6221\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6221\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__6233\,
            I => \N__6218\
        );

    \I__1139\ : Span4Mux_v
    port map (
            O => \N__6230\,
            I => \N__6215\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6227\,
            I => \N__6210\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6210\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6221\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1135\ : Odrv4
    port map (
            O => \N__6218\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__6215\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6210\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6198\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6198\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_a3_0_a3_0\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6192\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6192\,
            I => \N__6189\
        );

    \I__1128\ : Span4Mux_v
    port map (
            O => \N__6189\,
            I => \N__6185\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6182\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__6185\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6182\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6177\,
            I => \N__6174\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6171\
        );

    \I__1122\ : Span4Mux_v
    port map (
            O => \N__6171\,
            I => \N__6165\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6162\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6169\,
            I => \N__6157\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6168\,
            I => \N__6157\
        );

    \I__1118\ : Odrv4
    port map (
            O => \N__6165\,
            I => \U712_CHIP_RAM.N_328\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__6162\,
            I => \U712_CHIP_RAM.N_328\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6157\,
            I => \U712_CHIP_RAM.N_328\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__6150\,
            I => \N__6146\
        );

    \I__1114\ : CascadeMux
    port map (
            O => \N__6149\,
            I => \N__6143\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6146\,
            I => \N__6137\
        );

    \I__1112\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6137\
        );

    \I__1111\ : InMux
    port map (
            O => \N__6142\,
            I => \N__6129\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6137\,
            I => \N__6126\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6136\,
            I => \N__6123\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6135\,
            I => \N__6119\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__6134\,
            I => \N__6114\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6111\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6132\,
            I => \N__6103\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6129\,
            I => \N__6096\
        );

    \I__1103\ : Span4Mux_h
    port map (
            O => \N__6126\,
            I => \N__6096\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6123\,
            I => \N__6096\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__6122\,
            I => \N__6092\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6119\,
            I => \N__6087\
        );

    \I__1099\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6084\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6117\,
            I => \N__6078\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6114\,
            I => \N__6078\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__6111\,
            I => \N__6075\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6070\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6109\,
            I => \N__6070\
        );

    \I__1093\ : InMux
    port map (
            O => \N__6108\,
            I => \N__6063\
        );

    \I__1092\ : InMux
    port map (
            O => \N__6107\,
            I => \N__6063\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6106\,
            I => \N__6063\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__6103\,
            I => \N__6060\
        );

    \I__1089\ : Span4Mux_v
    port map (
            O => \N__6096\,
            I => \N__6057\
        );

    \I__1088\ : InMux
    port map (
            O => \N__6095\,
            I => \N__6048\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6048\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6091\,
            I => \N__6048\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6048\
        );

    \I__1084\ : Span4Mux_v
    port map (
            O => \N__6087\,
            I => \N__6043\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__6084\,
            I => \N__6043\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6083\,
            I => \N__6040\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__6078\,
            I => \N__6037\
        );

    \I__1080\ : Span4Mux_h
    port map (
            O => \N__6075\,
            I => \N__6030\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6070\,
            I => \N__6030\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6063\,
            I => \N__6030\
        );

    \I__1077\ : Odrv12
    port map (
            O => \N__6060\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__6057\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6048\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1074\ : Odrv4
    port map (
            O => \N__6043\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__6040\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1072\ : Odrv4
    port map (
            O => \N__6037\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__6030\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1070\ : CascadeMux
    port map (
            O => \N__6015\,
            I => \N__6008\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__6014\,
            I => \N__6004\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__6013\,
            I => \N__6001\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6012\,
            I => \N__5994\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6011\,
            I => \N__5994\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6008\,
            I => \N__5991\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6007\,
            I => \N__5988\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6004\,
            I => \N__5985\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5982\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__6000\,
            I => \N__5975\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__5999\,
            I => \N__5972\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5994\,
            I => \N__5963\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__5991\,
            I => \N__5963\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__5988\,
            I => \N__5963\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__5985\,
            I => \N__5960\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__5982\,
            I => \N__5957\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5954\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5951\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5948\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5978\,
            I => \N__5941\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5975\,
            I => \N__5941\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5941\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5936\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5970\,
            I => \N__5936\
        );

    \I__1046\ : Span4Mux_v
    port map (
            O => \N__5963\,
            I => \N__5933\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__5960\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__5957\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5954\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5951\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5948\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5941\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5936\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1038\ : Odrv4
    port map (
            O => \N__5933\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5916\,
            I => \N__5908\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5915\,
            I => \N__5908\
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__5914\,
            I => \N__5900\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5913\,
            I => \N__5895\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__5908\,
            I => \N__5891\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__5907\,
            I => \N__5887\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5906\,
            I => \N__5883\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5905\,
            I => \N__5878\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5878\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5903\,
            I => \N__5873\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5900\,
            I => \N__5873\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__5899\,
            I => \N__5870\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5898\,
            I => \N__5865\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__5895\,
            I => \N__5862\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5859\
        );

    \I__1022\ : Span4Mux_v
    port map (
            O => \N__5891\,
            I => \N__5856\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5890\,
            I => \N__5849\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5849\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5886\,
            I => \N__5849\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5883\,
            I => \N__5842\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5878\,
            I => \N__5842\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5873\,
            I => \N__5842\
        );

    \I__1015\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5835\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5835\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5868\,
            I => \N__5835\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5865\,
            I => \N__5830\
        );

    \I__1011\ : Span4Mux_h
    port map (
            O => \N__5862\,
            I => \N__5830\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__5859\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__5856\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5849\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1007\ : Odrv4
    port map (
            O => \N__5842\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__5835\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__5830\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5806\
        );

    \I__1003\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5806\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5815\,
            I => \N__5801\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5814\,
            I => \N__5801\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5813\,
            I => \N__5798\
        );

    \I__999\ : InMux
    port map (
            O => \N__5812\,
            I => \N__5795\
        );

    \I__998\ : InMux
    port map (
            O => \N__5811\,
            I => \N__5784\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5806\,
            I => \N__5778\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5801\,
            I => \N__5775\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5798\,
            I => \N__5771\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5795\,
            I => \N__5768\
        );

    \I__993\ : InMux
    port map (
            O => \N__5794\,
            I => \N__5765\
        );

    \I__992\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5758\
        );

    \I__991\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5758\
        );

    \I__990\ : InMux
    port map (
            O => \N__5791\,
            I => \N__5758\
        );

    \I__989\ : InMux
    port map (
            O => \N__5790\,
            I => \N__5753\
        );

    \I__988\ : InMux
    port map (
            O => \N__5789\,
            I => \N__5753\
        );

    \I__987\ : InMux
    port map (
            O => \N__5788\,
            I => \N__5748\
        );

    \I__986\ : InMux
    port map (
            O => \N__5787\,
            I => \N__5748\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__5784\,
            I => \N__5745\
        );

    \I__984\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5738\
        );

    \I__983\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5738\
        );

    \I__982\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5738\
        );

    \I__981\ : Span4Mux_v
    port map (
            O => \N__5778\,
            I => \N__5733\
        );

    \I__980\ : Span4Mux_h
    port map (
            O => \N__5775\,
            I => \N__5733\
        );

    \I__979\ : InMux
    port map (
            O => \N__5774\,
            I => \N__5730\
        );

    \I__978\ : Odrv4
    port map (
            O => \N__5771\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__977\ : Odrv4
    port map (
            O => \N__5768\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5765\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__5758\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__5753\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__5748\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__972\ : Odrv4
    port map (
            O => \N__5745\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__5738\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__970\ : Odrv4
    port map (
            O => \N__5733\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5730\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__5709\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_2_i_1_cascade_\
        );

    \I__967\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5702\
        );

    \I__966\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5691\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__5702\,
            I => \N__5688\
        );

    \I__964\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5685\
        );

    \I__963\ : InMux
    port map (
            O => \N__5700\,
            I => \N__5682\
        );

    \I__962\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5677\
        );

    \I__961\ : InMux
    port map (
            O => \N__5698\,
            I => \N__5677\
        );

    \I__960\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5672\
        );

    \I__959\ : InMux
    port map (
            O => \N__5696\,
            I => \N__5672\
        );

    \I__958\ : InMux
    port map (
            O => \N__5695\,
            I => \N__5663\
        );

    \I__957\ : InMux
    port map (
            O => \N__5694\,
            I => \N__5660\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5691\,
            I => \N__5655\
        );

    \I__955\ : Span4Mux_h
    port map (
            O => \N__5688\,
            I => \N__5655\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5685\,
            I => \N__5652\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5682\,
            I => \N__5645\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__5677\,
            I => \N__5645\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__5672\,
            I => \N__5645\
        );

    \I__950\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5638\
        );

    \I__949\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5638\
        );

    \I__948\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5638\
        );

    \I__947\ : InMux
    port map (
            O => \N__5668\,
            I => \N__5633\
        );

    \I__946\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5633\
        );

    \I__945\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5630\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5663\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__5660\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__942\ : Odrv4
    port map (
            O => \N__5655\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__941\ : Odrv4
    port map (
            O => \N__5652\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__940\ : Odrv4
    port map (
            O => \N__5645\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5638\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5633\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__5630\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__5613\,
            I => \N__5610\
        );

    \I__935\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5607\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5607\,
            I => \N__5604\
        );

    \I__933\ : Span4Mux_h
    port map (
            O => \N__5604\,
            I => \N__5601\
        );

    \I__932\ : Odrv4
    port map (
            O => \N__5601\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_2_i_2\
        );

    \I__931\ : InMux
    port map (
            O => \N__5598\,
            I => \N__5593\
        );

    \I__930\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5588\
        );

    \I__929\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5588\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5593\,
            I => \U712_REG_SM.N_210\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__5588\,
            I => \U712_REG_SM.N_210\
        );

    \I__926\ : InMux
    port map (
            O => \N__5583\,
            I => \N__5577\
        );

    \I__925\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5570\
        );

    \I__924\ : InMux
    port map (
            O => \N__5581\,
            I => \N__5570\
        );

    \I__923\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5570\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__5577\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__5570\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__5565\,
            I => \U712_REG_SM.N_248_cascade_\
        );

    \I__919\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5555\
        );

    \I__918\ : InMux
    port map (
            O => \N__5561\,
            I => \N__5552\
        );

    \I__917\ : InMux
    port map (
            O => \N__5560\,
            I => \N__5549\
        );

    \I__916\ : InMux
    port map (
            O => \N__5559\,
            I => \N__5544\
        );

    \I__915\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5544\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5555\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5552\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__5549\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5544\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__910\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5532\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5532\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_1_0\
        );

    \I__908\ : InMux
    port map (
            O => \N__5529\,
            I => \N__5526\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5526\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__906\ : InMux
    port map (
            O => \N__5523\,
            I => \bfn_10_8_0_\
        );

    \I__905\ : InMux
    port map (
            O => \N__5520\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__904\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5514\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5514\,
            I => \N__5511\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__5511\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__901\ : InMux
    port map (
            O => \N__5508\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__900\ : InMux
    port map (
            O => \N__5505\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__5502\,
            I => \N__5498\
        );

    \I__898\ : InMux
    port map (
            O => \N__5501\,
            I => \N__5495\
        );

    \I__897\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5492\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5495\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__5492\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__894\ : InMux
    port map (
            O => \N__5487\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__893\ : InMux
    port map (
            O => \N__5484\,
            I => \N__5480\
        );

    \I__892\ : InMux
    port map (
            O => \N__5483\,
            I => \N__5477\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__5480\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5477\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__889\ : InMux
    port map (
            O => \N__5472\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__888\ : InMux
    port map (
            O => \N__5469\,
            I => \N__5465\
        );

    \I__887\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5462\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5465\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5462\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__884\ : InMux
    port map (
            O => \N__5457\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__883\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5450\
        );

    \I__882\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5447\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5450\,
            I => \U712_CHIP_RAM.N_211\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5447\,
            I => \U712_CHIP_RAM.N_211\
        );

    \I__879\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5439\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__5439\,
            I => \N__5436\
        );

    \I__877\ : Odrv4
    port map (
            O => \N__5436\,
            I => \U712_CHIP_RAM.N_64_1\
        );

    \I__876\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5426\
        );

    \I__875\ : InMux
    port map (
            O => \N__5432\,
            I => \N__5426\
        );

    \I__874\ : InMux
    port map (
            O => \N__5431\,
            I => \N__5423\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5426\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5423\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__5418\,
            I => \U712_CHIP_RAM.N_64_1_cascade_\
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__5415\,
            I => \N__5411\
        );

    \I__869\ : InMux
    port map (
            O => \N__5414\,
            I => \N__5407\
        );

    \I__868\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5404\
        );

    \I__867\ : InMux
    port map (
            O => \N__5410\,
            I => \N__5401\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5407\,
            I => \N__5396\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5404\,
            I => \N__5396\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5401\,
            I => \U712_CHIP_RAM.N_340\
        );

    \I__863\ : Odrv4
    port map (
            O => \N__5396\,
            I => \U712_CHIP_RAM.N_340\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__5391\,
            I => \U712_CHIP_RAM.N_340_cascade_\
        );

    \I__861\ : InMux
    port map (
            O => \N__5388\,
            I => \N__5383\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__5387\,
            I => \N__5379\
        );

    \I__859\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5372\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5383\,
            I => \N__5369\
        );

    \I__857\ : InMux
    port map (
            O => \N__5382\,
            I => \N__5366\
        );

    \I__856\ : InMux
    port map (
            O => \N__5379\,
            I => \N__5363\
        );

    \I__855\ : InMux
    port map (
            O => \N__5378\,
            I => \N__5358\
        );

    \I__854\ : InMux
    port map (
            O => \N__5377\,
            I => \N__5358\
        );

    \I__853\ : InMux
    port map (
            O => \N__5376\,
            I => \N__5355\
        );

    \I__852\ : InMux
    port map (
            O => \N__5375\,
            I => \N__5352\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5372\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__5369\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__5366\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5363\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5358\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5355\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__5352\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\
        );

    \I__844\ : InMux
    port map (
            O => \N__5337\,
            I => \N__5334\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__5334\,
            I => \U712_CHIP_RAM.N_267\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__5331\,
            I => \U712_CHIP_RAM.N_281_cascade_\
        );

    \I__841\ : InMux
    port map (
            O => \N__5328\,
            I => \N__5325\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5325\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_0_i_0\
        );

    \I__839\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5316\
        );

    \I__838\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5316\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5316\,
            I => \U712_CHIP_RAM.N_207_i\
        );

    \I__836\ : InMux
    port map (
            O => \N__5313\,
            I => \N__5310\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__5310\,
            I => \N__5307\
        );

    \I__834\ : Span4Mux_v
    port map (
            O => \N__5307\,
            I => \N__5304\
        );

    \I__833\ : Sp12to4
    port map (
            O => \N__5304\,
            I => \N__5301\
        );

    \I__832\ : Span12Mux_h
    port map (
            O => \N__5301\,
            I => \N__5298\
        );

    \I__831\ : Odrv12
    port map (
            O => \N__5298\,
            I => \A_c_11\
        );

    \I__830\ : InMux
    port map (
            O => \N__5295\,
            I => \N__5292\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__5292\,
            I => \N__5289\
        );

    \I__828\ : Span12Mux_v
    port map (
            O => \N__5289\,
            I => \N__5286\
        );

    \I__827\ : Span12Mux_h
    port map (
            O => \N__5286\,
            I => \N__5283\
        );

    \I__826\ : Odrv12
    port map (
            O => \N__5283\,
            I => \A_c_4\
        );

    \I__825\ : InMux
    port map (
            O => \N__5280\,
            I => \N__5277\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5277\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__823\ : SRMux
    port map (
            O => \N__5274\,
            I => \N__5271\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5271\,
            I => \N__5268\
        );

    \I__821\ : Span4Mux_h
    port map (
            O => \N__5268\,
            I => \N__5265\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__5265\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__819\ : InMux
    port map (
            O => \N__5262\,
            I => \N__5259\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5259\,
            I => \N__5256\
        );

    \I__817\ : Span4Mux_v
    port map (
            O => \N__5256\,
            I => \N__5253\
        );

    \I__816\ : Sp12to4
    port map (
            O => \N__5253\,
            I => \N__5250\
        );

    \I__815\ : Span12Mux_h
    port map (
            O => \N__5250\,
            I => \N__5247\
        );

    \I__814\ : Span12Mux_v
    port map (
            O => \N__5247\,
            I => \N__5244\
        );

    \I__813\ : Odrv12
    port map (
            O => \N__5244\,
            I => \A_c_5\
        );

    \I__812\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5238\,
            I => \N__5235\
        );

    \I__810\ : Span12Mux_h
    port map (
            O => \N__5235\,
            I => \N__5232\
        );

    \I__809\ : Odrv12
    port map (
            O => \N__5232\,
            I => \A_c_12\
        );

    \I__808\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5226\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__5226\,
            I => \N__5223\
        );

    \I__806\ : Span4Mux_v
    port map (
            O => \N__5223\,
            I => \N__5220\
        );

    \I__805\ : Span4Mux_v
    port map (
            O => \N__5220\,
            I => \N__5217\
        );

    \I__804\ : Sp12to4
    port map (
            O => \N__5217\,
            I => \N__5214\
        );

    \I__803\ : Span12Mux_h
    port map (
            O => \N__5214\,
            I => \N__5211\
        );

    \I__802\ : Odrv12
    port map (
            O => \N__5211\,
            I => \A_c_7\
        );

    \I__801\ : CascadeMux
    port map (
            O => \N__5208\,
            I => \U712_CHIP_RAM.N_347_cascade_\
        );

    \I__800\ : CascadeMux
    port map (
            O => \N__5205\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_1_cascade_\
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__5202\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_cascade_\
        );

    \I__798\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5196\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5196\,
            I => \U712_CHIP_RAM.N_284\
        );

    \I__796\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5186\
        );

    \I__795\ : InMux
    port map (
            O => \N__5192\,
            I => \N__5186\
        );

    \I__794\ : InMux
    port map (
            O => \N__5191\,
            I => \N__5183\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5186\,
            I => \U712_REG_SM.N_215\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5183\,
            I => \U712_REG_SM.N_215\
        );

    \I__791\ : InMux
    port map (
            O => \N__5178\,
            I => \N__5174\
        );

    \I__790\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5171\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5174\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5171\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__787\ : CascadeMux
    port map (
            O => \N__5166\,
            I => \U712_REG_SM.N_215_cascade_\
        );

    \I__786\ : CascadeMux
    port map (
            O => \N__5163\,
            I => \U712_REG_SM.N_228_cascade_\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__5160\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_i_0_1_cascade_\
        );

    \I__784\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5154\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5154\,
            I => \N__5150\
        );

    \I__782\ : IoInMux
    port map (
            O => \N__5153\,
            I => \N__5147\
        );

    \I__781\ : Span4Mux_v
    port map (
            O => \N__5150\,
            I => \N__5144\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5147\,
            I => \N__5141\
        );

    \I__779\ : Sp12to4
    port map (
            O => \N__5144\,
            I => \N__5138\
        );

    \I__778\ : Span4Mux_s3_h
    port map (
            O => \N__5141\,
            I => \N__5135\
        );

    \I__777\ : Span12Mux_h
    port map (
            O => \N__5138\,
            I => \N__5130\
        );

    \I__776\ : Sp12to4
    port map (
            O => \N__5135\,
            I => \N__5130\
        );

    \I__775\ : Span12Mux_v
    port map (
            O => \N__5130\,
            I => \N__5127\
        );

    \I__774\ : Odrv12
    port map (
            O => \N__5127\,
            I => \C1_c\
        );

    \I__773\ : InMux
    port map (
            O => \N__5124\,
            I => \N__5120\
        );

    \I__772\ : IoInMux
    port map (
            O => \N__5123\,
            I => \N__5117\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5120\,
            I => \N__5114\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5117\,
            I => \N__5111\
        );

    \I__769\ : Span4Mux_v
    port map (
            O => \N__5114\,
            I => \N__5108\
        );

    \I__768\ : IoSpan4Mux
    port map (
            O => \N__5111\,
            I => \N__5105\
        );

    \I__767\ : Sp12to4
    port map (
            O => \N__5108\,
            I => \N__5102\
        );

    \I__766\ : IoSpan4Mux
    port map (
            O => \N__5105\,
            I => \N__5099\
        );

    \I__765\ : Span12Mux_h
    port map (
            O => \N__5102\,
            I => \N__5096\
        );

    \I__764\ : IoSpan4Mux
    port map (
            O => \N__5099\,
            I => \N__5093\
        );

    \I__763\ : Odrv12
    port map (
            O => \N__5096\,
            I => \C3_c\
        );

    \I__762\ : Odrv4
    port map (
            O => \N__5093\,
            I => \C3_c\
        );

    \I__761\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5085\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__5085\,
            I => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_1\
        );

    \I__759\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5079\,
            I => \N__5076\
        );

    \I__757\ : Span12Mux_h
    port map (
            O => \N__5076\,
            I => \N__5073\
        );

    \I__756\ : Odrv12
    port map (
            O => \N__5073\,
            I => \RAS1n_c\
        );

    \I__755\ : InMux
    port map (
            O => \N__5070\,
            I => \N__5064\
        );

    \I__754\ : InMux
    port map (
            O => \N__5069\,
            I => \N__5064\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5064\,
            I => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0\
        );

    \I__752\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5058\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__5058\,
            I => \N__5055\
        );

    \I__750\ : Span4Mux_v
    port map (
            O => \N__5055\,
            I => \N__5051\
        );

    \I__749\ : InMux
    port map (
            O => \N__5054\,
            I => \N__5048\
        );

    \I__748\ : Sp12to4
    port map (
            O => \N__5051\,
            I => \N__5045\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__5048\,
            I => \N__5042\
        );

    \I__746\ : Span12Mux_h
    port map (
            O => \N__5045\,
            I => \N__5039\
        );

    \I__745\ : Span12Mux_h
    port map (
            O => \N__5042\,
            I => \N__5036\
        );

    \I__744\ : Span12Mux_v
    port map (
            O => \N__5039\,
            I => \N__5033\
        );

    \I__743\ : Span12Mux_v
    port map (
            O => \N__5036\,
            I => \N__5030\
        );

    \I__742\ : Odrv12
    port map (
            O => \N__5033\,
            I => \TSn_c\
        );

    \I__741\ : Odrv12
    port map (
            O => \N__5030\,
            I => \TSn_c\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__5025\,
            I => \N__5022\
        );

    \I__739\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5019\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__5019\,
            I => \N__5016\
        );

    \I__737\ : Span4Mux_v
    port map (
            O => \N__5016\,
            I => \N__5013\
        );

    \I__736\ : Span4Mux_v
    port map (
            O => \N__5013\,
            I => \N__5010\
        );

    \I__735\ : Sp12to4
    port map (
            O => \N__5010\,
            I => \N__5007\
        );

    \I__734\ : Span12Mux_h
    port map (
            O => \N__5007\,
            I => \N__5004\
        );

    \I__733\ : Odrv12
    port map (
            O => \N__5004\,
            I => \REGSPACEn_c\
        );

    \I__732\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4998\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4998\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_2\
        );

    \I__730\ : CascadeMux
    port map (
            O => \N__4995\,
            I => \N__4991\
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__4994\,
            I => \N__4988\
        );

    \I__728\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4985\
        );

    \I__727\ : InMux
    port map (
            O => \N__4988\,
            I => \N__4982\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4985\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4982\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__724\ : InMux
    port map (
            O => \N__4977\,
            I => \N__4973\
        );

    \I__723\ : InMux
    port map (
            O => \N__4976\,
            I => \N__4970\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4973\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4970\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__4965\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_1_2_cascade_\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__4962\,
            I => \N__4958\
        );

    \I__718\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4955\
        );

    \I__717\ : InMux
    port map (
            O => \N__4958\,
            I => \N__4952\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4955\,
            I => \U712_REG_SM.N_245\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4952\,
            I => \U712_REG_SM.N_245\
        );

    \I__714\ : InMux
    port map (
            O => \N__4947\,
            I => \N__4944\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__4944\,
            I => \U712_CHIP_RAM.N_209\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__4941\,
            I => \U712_CHIP_RAM.N_209_cascade_\
        );

    \I__711\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4935\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4935\,
            I => \U712_CHIP_RAM.N_263\
        );

    \I__709\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4929\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4929\,
            I => \U712_CHIP_RAM.N_246\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__4926\,
            I => \N__4923\
        );

    \I__706\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4920\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4920\,
            I => \N__4911\
        );

    \I__704\ : InMux
    port map (
            O => \N__4919\,
            I => \N__4908\
        );

    \I__703\ : InMux
    port map (
            O => \N__4918\,
            I => \N__4904\
        );

    \I__702\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4901\
        );

    \I__701\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4898\
        );

    \I__700\ : InMux
    port map (
            O => \N__4915\,
            I => \N__4893\
        );

    \I__699\ : InMux
    port map (
            O => \N__4914\,
            I => \N__4893\
        );

    \I__698\ : Span4Mux_h
    port map (
            O => \N__4911\,
            I => \N__4888\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__4908\,
            I => \N__4888\
        );

    \I__696\ : InMux
    port map (
            O => \N__4907\,
            I => \N__4885\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4904\,
            I => \N__4882\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4901\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4898\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__4893\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__4888\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4885\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__4882\,
            I => \U712_CHIP_RAM.N_332\
        );

    \I__688\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4865\
        );

    \I__687\ : InMux
    port map (
            O => \N__4868\,
            I => \N__4862\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4865\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4862\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__684\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4850\
        );

    \I__683\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4850\
        );

    \I__682\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4847\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4850\,
            I => \N__4844\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4847\,
            I => \U712_CHIP_RAM.N_203\
        );

    \I__679\ : Odrv4
    port map (
            O => \N__4844\,
            I => \U712_CHIP_RAM.N_203\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__4839\,
            I => \U712_CHIP_RAM.N_203_cascade_\
        );

    \I__677\ : CascadeMux
    port map (
            O => \N__4836\,
            I => \N__4833\
        );

    \I__676\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4830\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__4830\,
            I => \N__4827\
        );

    \I__674\ : Odrv4
    port map (
            O => \N__4827\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_3_0\
        );

    \I__673\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4818\
        );

    \I__672\ : InMux
    port map (
            O => \N__4823\,
            I => \N__4818\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4818\,
            I => \U712_CHIP_RAM.N_341\
        );

    \I__670\ : CEMux
    port map (
            O => \N__4815\,
            I => \N__4812\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__4812\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__4809\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7_cascade_\
        );

    \I__667\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4803\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__4803\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_0_0_i_1\
        );

    \I__665\ : CascadeMux
    port map (
            O => \N__4800\,
            I => \U712_CHIP_RAM.N_211_cascade_\
        );

    \I__664\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4794\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__4794\,
            I => \U712_CHIP_RAM.N_87\
        );

    \I__662\ : InMux
    port map (
            O => \N__4791\,
            I => \N__4788\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4788\,
            I => \U712_CHIP_RAM.N_266\
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__4785\,
            I => \N__4778\
        );

    \I__659\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4775\
        );

    \I__658\ : InMux
    port map (
            O => \N__4783\,
            I => \N__4772\
        );

    \I__657\ : InMux
    port map (
            O => \N__4782\,
            I => \N__4767\
        );

    \I__656\ : InMux
    port map (
            O => \N__4781\,
            I => \N__4767\
        );

    \I__655\ : InMux
    port map (
            O => \N__4778\,
            I => \N__4763\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4775\,
            I => \N__4756\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4772\,
            I => \N__4756\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__4767\,
            I => \N__4756\
        );

    \I__651\ : InMux
    port map (
            O => \N__4766\,
            I => \N__4753\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4763\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__649\ : Odrv4
    port map (
            O => \N__4756\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4753\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__647\ : CascadeMux
    port map (
            O => \N__4746\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a3_0_0_cascade_\
        );

    \I__646\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4739\
        );

    \I__645\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4736\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4739\,
            I => \N__4733\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4736\,
            I => \U712_CHIP_RAM.N_264\
        );

    \I__642\ : Odrv4
    port map (
            O => \N__4733\,
            I => \U712_CHIP_RAM.N_264\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__4728\,
            I => \U712_CHIP_RAM.N_264_cascade_\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__4725\,
            I => \U712_CHIP_RAM.N_36_cascade_\
        );

    \I__639\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4718\
        );

    \I__638\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4715\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4718\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__4715\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1\
        );

    \I__635\ : CascadeMux
    port map (
            O => \N__4710\,
            I => \U712_CHIP_RAM.N_342_cascade_\
        );

    \I__634\ : InMux
    port map (
            O => \N__4707\,
            I => \N__4703\
        );

    \I__633\ : InMux
    port map (
            O => \N__4706\,
            I => \N__4700\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__4703\,
            I => \U712_CHIP_RAM.N_381\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4700\,
            I => \U712_CHIP_RAM.N_381\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__4695\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\
        );

    \I__629\ : InMux
    port map (
            O => \N__4692\,
            I => \N__4689\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__4689\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_0\
        );

    \I__627\ : CascadeMux
    port map (
            O => \N__4686\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_1_cascade_\
        );

    \I__626\ : InMux
    port map (
            O => \N__4683\,
            I => \N__4680\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4680\,
            I => \N__4677\
        );

    \I__624\ : Sp12to4
    port map (
            O => \N__4677\,
            I => \N__4674\
        );

    \I__623\ : Span12Mux_v
    port map (
            O => \N__4674\,
            I => \N__4671\
        );

    \I__622\ : Span12Mux_h
    port map (
            O => \N__4671\,
            I => \N__4668\
        );

    \I__621\ : Odrv12
    port map (
            O => \N__4668\,
            I => \A_c_8\
        );

    \I__620\ : InMux
    port map (
            O => \N__4665\,
            I => \N__4662\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4662\,
            I => \N__4659\
        );

    \I__618\ : Span4Mux_v
    port map (
            O => \N__4659\,
            I => \N__4656\
        );

    \I__617\ : Span4Mux_v
    port map (
            O => \N__4656\,
            I => \N__4653\
        );

    \I__616\ : Sp12to4
    port map (
            O => \N__4653\,
            I => \N__4650\
        );

    \I__615\ : Odrv12
    port map (
            O => \N__4650\,
            I => \A_c_15\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__4647\,
            I => \N__4644\
        );

    \I__613\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4640\
        );

    \I__612\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4637\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__4640\,
            I => \U712_CHIP_RAM.N_270_4\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__4637\,
            I => \U712_CHIP_RAM.N_270_4\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__4632\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_i_0_3_cascade_\
        );

    \I__608\ : InMux
    port map (
            O => \N__4629\,
            I => \N__4626\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__4626\,
            I => \U712_REG_SM.N_289\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__4623\,
            I => \U712_REG_SM.N_289_cascade_\
        );

    \I__605\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4608\
        );

    \I__604\ : InMux
    port map (
            O => \N__4619\,
            I => \N__4608\
        );

    \I__603\ : InMux
    port map (
            O => \N__4618\,
            I => \N__4608\
        );

    \I__602\ : InMux
    port map (
            O => \N__4617\,
            I => \N__4608\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__4608\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__600\ : InMux
    port map (
            O => \N__4605\,
            I => \N__4602\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4602\,
            I => \N__4597\
        );

    \I__598\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4594\
        );

    \I__597\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4591\
        );

    \I__596\ : Span4Mux_h
    port map (
            O => \N__4597\,
            I => \N__4583\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4594\,
            I => \N__4583\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__4591\,
            I => \N__4583\
        );

    \I__593\ : InMux
    port map (
            O => \N__4590\,
            I => \N__4580\
        );

    \I__592\ : Span4Mux_v
    port map (
            O => \N__4583\,
            I => \N__4577\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4580\,
            I => \N__4574\
        );

    \I__590\ : Sp12to4
    port map (
            O => \N__4577\,
            I => \N__4571\
        );

    \I__589\ : Span4Mux_v
    port map (
            O => \N__4574\,
            I => \N__4568\
        );

    \I__588\ : Span12Mux_h
    port map (
            O => \N__4571\,
            I => \N__4565\
        );

    \I__587\ : Span4Mux_h
    port map (
            O => \N__4568\,
            I => \N__4562\
        );

    \I__586\ : Span12Mux_v
    port map (
            O => \N__4565\,
            I => \N__4559\
        );

    \I__585\ : Span4Mux_h
    port map (
            O => \N__4562\,
            I => \N__4556\
        );

    \I__584\ : Odrv12
    port map (
            O => \N__4559\,
            I => \RnW_c\
        );

    \I__583\ : Odrv4
    port map (
            O => \N__4556\,
            I => \RnW_c\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__4551\,
            I => \U712_CHIP_RAM.N_261_cascade_\
        );

    \I__581\ : IoInMux
    port map (
            O => \N__4548\,
            I => \N__4545\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4545\,
            I => \N__4542\
        );

    \I__579\ : IoSpan4Mux
    port map (
            O => \N__4542\,
            I => \N__4539\
        );

    \I__578\ : Sp12to4
    port map (
            O => \N__4539\,
            I => \N__4536\
        );

    \I__577\ : Span12Mux_s7_h
    port map (
            O => \N__4536\,
            I => \N__4533\
        );

    \I__576\ : Span12Mux_h
    port map (
            O => \N__4533\,
            I => \N__4529\
        );

    \I__575\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4526\
        );

    \I__574\ : Odrv12
    port map (
            O => \N__4529\,
            I => \CLK_EN_c\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4526\,
            I => \CLK_EN_c\
        );

    \I__572\ : InMux
    port map (
            O => \N__4521\,
            I => \N__4518\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4518\,
            I => \U712_CHIP_RAM.N_260\
        );

    \I__570\ : CascadeMux
    port map (
            O => \N__4515\,
            I => \N__4512\
        );

    \I__569\ : InMux
    port map (
            O => \N__4512\,
            I => \N__4508\
        );

    \I__568\ : InMux
    port map (
            O => \N__4511\,
            I => \N__4505\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4508\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4505\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__565\ : InMux
    port map (
            O => \N__4500\,
            I => \N__4488\
        );

    \I__564\ : InMux
    port map (
            O => \N__4499\,
            I => \N__4488\
        );

    \I__563\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4488\
        );

    \I__562\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4488\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__4488\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__560\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4482\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4482\,
            I => \N__4478\
        );

    \I__558\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4475\
        );

    \I__557\ : Span4Mux_v
    port map (
            O => \N__4478\,
            I => \N__4472\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4475\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__555\ : Odrv4
    port map (
            O => \N__4472\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__554\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4464\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4464\,
            I => \N__4461\
        );

    \I__552\ : Odrv4
    port map (
            O => \N__4461\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__4458\,
            I => \N__4455\
        );

    \I__550\ : InMux
    port map (
            O => \N__4455\,
            I => \N__4452\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4452\,
            I => \N__4448\
        );

    \I__548\ : InMux
    port map (
            O => \N__4451\,
            I => \N__4445\
        );

    \I__547\ : Span4Mux_v
    port map (
            O => \N__4448\,
            I => \N__4442\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__4445\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__4442\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__544\ : InMux
    port map (
            O => \N__4437\,
            I => \N__4434\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4434\,
            I => \N__4431\
        );

    \I__542\ : Odrv12
    port map (
            O => \N__4431\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__4428\,
            I => \N__4425\
        );

    \I__540\ : InMux
    port map (
            O => \N__4425\,
            I => \N__4422\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4422\,
            I => \N__4419\
        );

    \I__538\ : Span4Mux_h
    port map (
            O => \N__4419\,
            I => \N__4415\
        );

    \I__537\ : IoInMux
    port map (
            O => \N__4418\,
            I => \N__4412\
        );

    \I__536\ : Sp12to4
    port map (
            O => \N__4415\,
            I => \N__4409\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4412\,
            I => \N__4406\
        );

    \I__534\ : Span12Mux_v
    port map (
            O => \N__4409\,
            I => \N__4403\
        );

    \I__533\ : IoSpan4Mux
    port map (
            O => \N__4406\,
            I => \N__4400\
        );

    \I__532\ : Odrv12
    port map (
            O => \N__4403\,
            I => \RAMENn_c\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__4400\,
            I => \RAMENn_c\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__4395\,
            I => \N__4392\
        );

    \I__529\ : InMux
    port map (
            O => \N__4392\,
            I => \N__4388\
        );

    \I__528\ : InMux
    port map (
            O => \N__4391\,
            I => \N__4385\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4388\,
            I => \REG_TACK\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4385\,
            I => \REG_TACK\
        );

    \I__525\ : InMux
    port map (
            O => \N__4380\,
            I => \N__4377\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4377\,
            I => \U712_REG_SM.N_225\
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__4374\,
            I => \U712_REG_SM.N_225_cascade_\
        );

    \I__522\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4368\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4368\,
            I => \U712_REG_SM.N_292\
        );

    \I__520\ : InMux
    port map (
            O => \N__4365\,
            I => \N__4362\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4362\,
            I => \U712_REG_SM.REG_TACK_RNOZ0Z_0\
        );

    \I__518\ : CascadeMux
    port map (
            O => \N__4359\,
            I => \U712_CHIP_RAM.N_332_cascade_\
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__4356\,
            I => \N__4353\
        );

    \I__516\ : InMux
    port map (
            O => \N__4353\,
            I => \N__4350\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4350\,
            I => \U712_CHIP_RAM.A_m_2_20\
        );

    \I__514\ : InMux
    port map (
            O => \N__4347\,
            I => \N__4344\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__512\ : Span4Mux_v
    port map (
            O => \N__4341\,
            I => \N__4338\
        );

    \I__511\ : Sp12to4
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__510\ : Span12Mux_h
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__509\ : Span12Mux_v
    port map (
            O => \N__4332\,
            I => \N__4329\
        );

    \I__508\ : Odrv12
    port map (
            O => \N__4329\,
            I => \A_c_20\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__4326\,
            I => \U712_CHIP_RAM.A_m_2_20_cascade_\
        );

    \I__506\ : CascadeMux
    port map (
            O => \N__4323\,
            I => \U712_CHIP_RAM.BANK0_esr_RNOZ0Z_1_cascade_\
        );

    \I__505\ : IoInMux
    port map (
            O => \N__4320\,
            I => \N__4317\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__4317\,
            I => \N__4314\
        );

    \I__503\ : Span4Mux_s3_v
    port map (
            O => \N__4314\,
            I => \N__4311\
        );

    \I__502\ : Span4Mux_v
    port map (
            O => \N__4311\,
            I => \N__4308\
        );

    \I__501\ : Span4Mux_v
    port map (
            O => \N__4308\,
            I => \N__4305\
        );

    \I__500\ : Span4Mux_h
    port map (
            O => \N__4305\,
            I => \N__4302\
        );

    \I__499\ : Odrv4
    port map (
            O => \N__4302\,
            I => \BANK0_c\
        );

    \I__498\ : CEMux
    port map (
            O => \N__4299\,
            I => \N__4296\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4296\,
            I => \N__4293\
        );

    \I__496\ : Odrv4
    port map (
            O => \N__4293\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_10_0_0\
        );

    \I__495\ : InMux
    port map (
            O => \N__4290\,
            I => \N__4287\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__4287\,
            I => \N__4284\
        );

    \I__493\ : Odrv4
    port map (
            O => \N__4284\,
            I => \U712_CHIP_RAM.CPU_TACK_e_1\
        );

    \I__492\ : InMux
    port map (
            O => \N__4281\,
            I => \N__4277\
        );

    \I__491\ : InMux
    port map (
            O => \N__4280\,
            I => \N__4274\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4277\,
            I => \CPU_TACKm\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4274\,
            I => \CPU_TACKm\
        );

    \I__488\ : IoInMux
    port map (
            O => \N__4269\,
            I => \N__4266\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4266\,
            I => \N__4263\
        );

    \I__486\ : IoSpan4Mux
    port map (
            O => \N__4263\,
            I => \N__4260\
        );

    \I__485\ : Span4Mux_s0_h
    port map (
            O => \N__4260\,
            I => \N__4257\
        );

    \I__484\ : Sp12to4
    port map (
            O => \N__4257\,
            I => \N__4254\
        );

    \I__483\ : Span12Mux_s11_h
    port map (
            O => \N__4254\,
            I => \N__4250\
        );

    \I__482\ : InMux
    port map (
            O => \N__4253\,
            I => \N__4247\
        );

    \I__481\ : Odrv12
    port map (
            O => \N__4250\,
            I => \TACK_OUTn\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4247\,
            I => \TACK_OUTn\
        );

    \I__479\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4237\
        );

    \I__478\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4234\
        );

    \I__477\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4231\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4237\,
            I => \N__4228\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__4234\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4231\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__473\ : Odrv4
    port map (
            O => \N__4228\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__4221\,
            I => \N__4217\
        );

    \I__471\ : InMux
    port map (
            O => \N__4220\,
            I => \N__4214\
        );

    \I__470\ : InMux
    port map (
            O => \N__4217\,
            I => \N__4210\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4214\,
            I => \N__4207\
        );

    \I__468\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4204\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4210\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__466\ : Odrv4
    port map (
            O => \N__4207\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4204\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__464\ : InMux
    port map (
            O => \N__4197\,
            I => \N__4194\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4194\,
            I => \U712_CHIP_RAM.N_243\
        );

    \I__462\ : InMux
    port map (
            O => \N__4191\,
            I => \N__4188\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4188\,
            I => \N__4185\
        );

    \I__460\ : Span12Mux_v
    port map (
            O => \N__4185\,
            I => \N__4182\
        );

    \I__459\ : Odrv12
    port map (
            O => \N__4182\,
            I => \A_c_13\
        );

    \I__458\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4176\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__4176\,
            I => \N__4173\
        );

    \I__456\ : Span4Mux_h
    port map (
            O => \N__4173\,
            I => \N__4170\
        );

    \I__455\ : Sp12to4
    port map (
            O => \N__4170\,
            I => \N__4167\
        );

    \I__454\ : Span12Mux_v
    port map (
            O => \N__4167\,
            I => \N__4164\
        );

    \I__453\ : Odrv12
    port map (
            O => \N__4164\,
            I => \A_c_6\
        );

    \I__452\ : InMux
    port map (
            O => \N__4161\,
            I => \N__4158\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__4158\,
            I => \N__4155\
        );

    \I__450\ : Span4Mux_h
    port map (
            O => \N__4155\,
            I => \N__4152\
        );

    \I__449\ : Sp12to4
    port map (
            O => \N__4152\,
            I => \N__4149\
        );

    \I__448\ : Span12Mux_v
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__447\ : Odrv12
    port map (
            O => \N__4146\,
            I => \A_c_18\
        );

    \I__446\ : InMux
    port map (
            O => \N__4143\,
            I => \N__4140\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4140\,
            I => \N__4137\
        );

    \I__444\ : Span4Mux_v
    port map (
            O => \N__4137\,
            I => \N__4134\
        );

    \I__443\ : Span4Mux_v
    port map (
            O => \N__4134\,
            I => \N__4131\
        );

    \I__442\ : Sp12to4
    port map (
            O => \N__4131\,
            I => \N__4128\
        );

    \I__441\ : Span12Mux_h
    port map (
            O => \N__4128\,
            I => \N__4125\
        );

    \I__440\ : Odrv12
    port map (
            O => \N__4125\,
            I => \A_c_16\
        );

    \I__439\ : IoInMux
    port map (
            O => \N__4122\,
            I => \N__4119\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__4119\,
            I => \N__4116\
        );

    \I__437\ : Span12Mux_s4_v
    port map (
            O => \N__4116\,
            I => \N__4113\
        );

    \I__436\ : Odrv12
    port map (
            O => \N__4113\,
            I => \N_187_i\
        );

    \I__435\ : CascadeMux
    port map (
            O => \N__4110\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_0_a3_0_cascade_\
        );

    \I__434\ : CascadeMux
    port map (
            O => \N__4107\,
            I => \N__4104\
        );

    \I__433\ : InMux
    port map (
            O => \N__4104\,
            I => \N__4101\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4101\,
            I => \N__4097\
        );

    \I__431\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4094\
        );

    \I__430\ : Span4Mux_h
    port map (
            O => \N__4097\,
            I => \N__4091\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4094\,
            I => \U712_CHIP_RAM.N_273\
        );

    \I__428\ : Odrv4
    port map (
            O => \N__4091\,
            I => \U712_CHIP_RAM.N_273\
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__4086\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1_cascade_\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__4083\,
            I => \U712_CHIP_RAM.N_328_cascade_\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__4080\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__4077\,
            I => \U712_CYCLE_TERM.N_223_i_0_en_cascade_\
        );

    \I__423\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4071\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__4071\,
            I => \N__4068\
        );

    \I__421\ : Odrv4
    port map (
            O => \N__4068\,
            I => \TACK_EN_i_ess\
        );

    \I__420\ : CEMux
    port map (
            O => \N__4065\,
            I => \N__4062\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__4062\,
            I => \N__4059\
        );

    \I__418\ : Span4Mux_v
    port map (
            O => \N__4059\,
            I => \N__4056\
        );

    \I__417\ : Span4Mux_h
    port map (
            O => \N__4056\,
            I => \N__4053\
        );

    \I__416\ : Odrv4
    port map (
            O => \N__4053\,
            I => \U712_CYCLE_TERM.N_223_i_0_en_0\
        );

    \I__415\ : InMux
    port map (
            O => \N__4050\,
            I => \N__4047\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__4047\,
            I => \N__4043\
        );

    \I__413\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4040\
        );

    \I__412\ : Span4Mux_v
    port map (
            O => \N__4043\,
            I => \N__4034\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__4040\,
            I => \N__4034\
        );

    \I__410\ : InMux
    port map (
            O => \N__4039\,
            I => \N__4031\
        );

    \I__409\ : Span4Mux_h
    port map (
            O => \N__4034\,
            I => \N__4028\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__4031\,
            I => \N__4025\
        );

    \I__407\ : Sp12to4
    port map (
            O => \N__4028\,
            I => \N__4022\
        );

    \I__406\ : Span4Mux_v
    port map (
            O => \N__4025\,
            I => \N__4019\
        );

    \I__405\ : Span12Mux_v
    port map (
            O => \N__4022\,
            I => \N__4016\
        );

    \I__404\ : IoSpan4Mux
    port map (
            O => \N__4019\,
            I => \N__4013\
        );

    \I__403\ : Odrv12
    port map (
            O => \N__4016\,
            I => \AWEn_c\
        );

    \I__402\ : Odrv4
    port map (
            O => \N__4013\,
            I => \AWEn_c\
        );

    \I__401\ : IoInMux
    port map (
            O => \N__4008\,
            I => \N__4005\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__4005\,
            I => \N__4002\
        );

    \I__399\ : IoSpan4Mux
    port map (
            O => \N__4002\,
            I => \N__3999\
        );

    \I__398\ : Span4Mux_s3_h
    port map (
            O => \N__3999\,
            I => \N__3996\
        );

    \I__397\ : Sp12to4
    port map (
            O => \N__3996\,
            I => \N__3993\
        );

    \I__396\ : Span12Mux_s6_v
    port map (
            O => \N__3993\,
            I => \N__3990\
        );

    \I__395\ : Span12Mux_h
    port map (
            O => \N__3990\,
            I => \N__3987\
        );

    \I__394\ : Odrv12
    port map (
            O => \N__3987\,
            I => \N_242\
        );

    \I__393\ : InMux
    port map (
            O => \N__3984\,
            I => \N__3980\
        );

    \I__392\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3977\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__3980\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3977\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__389\ : InMux
    port map (
            O => \N__3972\,
            I => \N__3968\
        );

    \I__388\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3965\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3968\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__3965\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__385\ : CascadeMux
    port map (
            O => \N__3960\,
            I => \N__3956\
        );

    \I__384\ : InMux
    port map (
            O => \N__3959\,
            I => \N__3953\
        );

    \I__383\ : InMux
    port map (
            O => \N__3956\,
            I => \N__3950\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3953\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__3950\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__380\ : InMux
    port map (
            O => \N__3945\,
            I => \N__3941\
        );

    \I__379\ : InMux
    port map (
            O => \N__3944\,
            I => \N__3938\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__3941\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__3938\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__376\ : CascadeMux
    port map (
            O => \N__3933\,
            I => \U712_CHIP_RAM.N_381_cascade_\
        );

    \I__375\ : IoInMux
    port map (
            O => \N__3930\,
            I => \N__3927\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3927\,
            I => \N__3924\
        );

    \I__373\ : Span12Mux_s9_v
    port map (
            O => \N__3924\,
            I => \N__3921\
        );

    \I__372\ : Odrv12
    port map (
            O => \N__3921\,
            I => \VBENn_c\
        );

    \I__371\ : InMux
    port map (
            O => \N__3918\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__370\ : InMux
    port map (
            O => \N__3915\,
            I => \N__3911\
        );

    \I__369\ : InMux
    port map (
            O => \N__3914\,
            I => \N__3908\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3911\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__3908\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__366\ : InMux
    port map (
            O => \N__3903\,
            I => \N__3899\
        );

    \I__365\ : InMux
    port map (
            O => \N__3902\,
            I => \N__3896\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3899\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3896\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__362\ : IoInMux
    port map (
            O => \N__3891\,
            I => \N__3888\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__3888\,
            I => \N__3884\
        );

    \I__360\ : CascadeMux
    port map (
            O => \N__3887\,
            I => \N__3881\
        );

    \I__359\ : Span12Mux_s7_v
    port map (
            O => \N__3884\,
            I => \N__3878\
        );

    \I__358\ : InMux
    port map (
            O => \N__3881\,
            I => \N__3875\
        );

    \I__357\ : Odrv12
    port map (
            O => \N__3878\,
            I => \DBDIR_c\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__3875\,
            I => \DBDIR_c\
        );

    \I__355\ : CascadeMux
    port map (
            O => \N__3870\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0_cascade_\
        );

    \I__354\ : InMux
    port map (
            O => \N__3867\,
            I => \N__3862\
        );

    \I__353\ : InMux
    port map (
            O => \N__3866\,
            I => \N__3857\
        );

    \I__352\ : InMux
    port map (
            O => \N__3865\,
            I => \N__3857\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3862\,
            I => \N__3854\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__3857\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_a3_0_0\
        );

    \I__349\ : Odrv4
    port map (
            O => \N__3854\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_a3_0_0\
        );

    \I__348\ : IoInMux
    port map (
            O => \N__3849\,
            I => \N__3846\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__3846\,
            I => \N__3843\
        );

    \I__346\ : Span4Mux_s2_v
    port map (
            O => \N__3843\,
            I => \N__3840\
        );

    \I__345\ : Span4Mux_v
    port map (
            O => \N__3840\,
            I => \N__3837\
        );

    \I__344\ : Span4Mux_h
    port map (
            O => \N__3837\,
            I => \N__3834\
        );

    \I__343\ : Odrv4
    port map (
            O => \N__3834\,
            I => \CLK80_PLL_i_i\
        );

    \I__342\ : IoInMux
    port map (
            O => \N__3831\,
            I => \N__3828\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__3828\,
            I => \N__3825\
        );

    \I__340\ : Span4Mux_s2_h
    port map (
            O => \N__3825\,
            I => \N__3822\
        );

    \I__339\ : Sp12to4
    port map (
            O => \N__3822\,
            I => \N__3819\
        );

    \I__338\ : Span12Mux_v
    port map (
            O => \N__3819\,
            I => \N__3816\
        );

    \I__337\ : Odrv12
    port map (
            O => \N__3816\,
            I => \N_1012_i\
        );

    \I__336\ : InMux
    port map (
            O => \N__3813\,
            I => \bfn_7_5_0_\
        );

    \I__335\ : InMux
    port map (
            O => \N__3810\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__334\ : InMux
    port map (
            O => \N__3807\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__333\ : InMux
    port map (
            O => \N__3804\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__332\ : InMux
    port map (
            O => \N__3801\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__331\ : InMux
    port map (
            O => \N__3798\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__330\ : InMux
    port map (
            O => \N__3795\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__329\ : IoInMux
    port map (
            O => \N__3792\,
            I => \N__3789\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__3789\,
            I => \N__3786\
        );

    \I__327\ : IoSpan4Mux
    port map (
            O => \N__3786\,
            I => \N__3783\
        );

    \I__326\ : Span4Mux_s2_v
    port map (
            O => \N__3783\,
            I => \N__3780\
        );

    \I__325\ : Sp12to4
    port map (
            O => \N__3780\,
            I => \N__3777\
        );

    \I__324\ : Span12Mux_v
    port map (
            O => \N__3777\,
            I => \N__3774\
        );

    \I__323\ : Odrv12
    port map (
            O => \N__3774\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__7733\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__7734\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__7731\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__7732\
        );

    \IN_MUX_bfv_10_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_8_0_\
        );

    \IN_MUX_bfv_7_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_5_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7560\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5153\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5123\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8736\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4074\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_1012_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3945\,
            in2 => \_gnd_net_\,
            in3 => \N__3813\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_7_5_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__5274\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3972\,
            in2 => \_gnd_net_\,
            in3 => \N__3810\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__5274\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3984\,
            in2 => \_gnd_net_\,
            in3 => \N__3807\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__5274\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4481\,
            in2 => \_gnd_net_\,
            in3 => \N__3804\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__5274\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3959\,
            in2 => \_gnd_net_\,
            in3 => \N__3801\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__5274\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3903\,
            in2 => \_gnd_net_\,
            in3 => \N__3798\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__5274\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3915\,
            in2 => \_gnd_net_\,
            in3 => \N__3795\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__5274\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4451\,
            in2 => \_gnd_net_\,
            in3 => \N__3918\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7730\,
            ce => 'H',
            sr => \N__5274\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100101111"
        )
    port map (
            in0 => \N__9615\,
            in1 => \N__7349\,
            in2 => \N__8456\,
            in3 => \N__7275\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3914\,
            in2 => \_gnd_net_\,
            in3 => \N__3902\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__4100\,
            in1 => \N__9619\,
            in2 => \N__4356\,
            in3 => \N__6135\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8719\,
            ce => 'H',
            sr => \N__10115\
        );

    \U712_CHIP_RAM.DBDIR_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111010011110000"
        )
    port map (
            in0 => \N__4050\,
            in1 => \N__3867\,
            in2 => \N__3887\,
            in3 => \N__4917\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8719\,
            ce => 'H',
            sr => \N__10115\
        );

    \U712_CHIP_RAM.DMA_CYCLE_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__4915\,
            in1 => \N__9476\,
            in2 => \N__4107\,
            in3 => \N__3866\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8723\,
            ce => 'H',
            sr => \N__10109\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__3865\,
            in1 => \N__4743\,
            in2 => \_gnd_net_\,
            in3 => \N__4914\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101011111010"
        )
    port map (
            in0 => \N__9358\,
            in1 => \N__5813\,
            in2 => \N__3870\,
            in3 => \N__8040\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8723\,
            ce => 'H',
            sr => \N__10109\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6250\,
            in2 => \_gnd_net_\,
            in3 => \N__6118\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__6251\,
            in1 => \N__4046\,
            in2 => \_gnd_net_\,
            in3 => \N__4605\,
            lcout => \U712_CHIP_RAM.N_243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4280\,
            in2 => \_gnd_net_\,
            in3 => \N__4391\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__7698\,
            in1 => \N__4213\,
            in2 => \N__4080\,
            in3 => \N__4511\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_223_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10139\,
            in1 => \_gnd_net_\,
            in2 => \N__4077\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_223_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__4220\,
            in1 => \N__7697\,
            in2 => \_gnd_net_\,
            in3 => \N__4241\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8730\,
            ce => \N__4065\,
            sr => \N__10096\
        );

    \U712_BUFFERS.DRDDIR_i_m2_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__4590\,
            in1 => \N__4039\,
            in2 => \_gnd_net_\,
            in3 => \N__9523\,
            lcout => \N_242\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__3983\,
            in1 => \N__3971\,
            in2 => \N__3960\,
            in3 => \N__3944\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4JG83_2_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5814\,
            in1 => \N__5696\,
            in2 => \_gnd_net_\,
            in3 => \N__6168\,
            lcout => \U712_CHIP_RAM.N_381\,
            ltout => \U712_CHIP_RAM.N_381_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__6169\,
            in1 => \N__4643\,
            in2 => \N__3933\,
            in3 => \N__5916\,
            lcout => \U712_CHIP_RAM.CPU_TACK_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a3_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8523\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9620\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__4191\,
            in1 => \_gnd_net_\,
            in2 => \N__8403\,
            in3 => \N__4179\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4161\,
            in1 => \N__4143\,
            in2 => \_gnd_net_\,
            in3 => \N__8364\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_187_i_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110001"
        )
    port map (
            in0 => \N__9621\,
            in1 => \N__8766\,
            in2 => \N__9860\,
            in3 => \N__10207\,
            lcout => \N_187_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000101000000"
        )
    port map (
            in0 => \N__5815\,
            in1 => \N__5697\,
            in2 => \N__6015\,
            in3 => \N__4783\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_6_0_0_0_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6133\,
            in1 => \N__5915\,
            in2 => \N__4110\,
            in3 => \N__5382\,
            lcout => \U712_CHIP_RAM.N_273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNI4ICS5_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__4907\,
            in1 => \N__6289\,
            in2 => \N__6258\,
            in3 => \N__4857\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__4742\,
            in1 => \N__10140\,
            in2 => \N__4086\,
            in3 => \N__6136\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI85LA2_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6007\,
            in2 => \_gnd_net_\,
            in3 => \N__5375\,
            lcout => \U712_CHIP_RAM.N_328\,
            ltout => \U712_CHIP_RAM.N_328_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5774\,
            in1 => \N__5913\,
            in2 => \N__4083\,
            in3 => \N__5666\,
            lcout => \U712_CHIP_RAM.N_332\,
            ltout => \U712_CHIP_RAM.N_332_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNI4ICS5_0_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6256\,
            in1 => \N__6288\,
            in2 => \N__4359\,
            in3 => \N__4856\,
            lcout => \U712_CHIP_RAM.A_m_2_20\,
            ltout => \U712_CHIP_RAM.A_m_2_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4347\,
            in2 => \N__4326\,
            in3 => \N__9129\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.BANK0_esr_RNOZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__6257\,
            in1 => \N__4916\,
            in2 => \N__4323\,
            in3 => \N__7137\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8715\,
            ce => \N__4299\,
            sr => \N__10110\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__6705\,
            in1 => \N__4240\,
            in2 => \N__4515\,
            in3 => \N__4497\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8720\,
            ce => 'H',
            sr => \N__10100\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010111000"
        )
    port map (
            in0 => \N__4281\,
            in1 => \N__4797\,
            in2 => \N__9660\,
            in3 => \N__4290\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8720\,
            ce => 'H',
            sr => \N__10100\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110100010"
        )
    port map (
            in0 => \N__4253\,
            in1 => \N__4499\,
            in2 => \N__7914\,
            in3 => \N__6736\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8720\,
            ce => 'H',
            sr => \N__10100\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101010110000"
        )
    port map (
            in0 => \N__4500\,
            in1 => \N__4242\,
            in2 => \N__4221\,
            in3 => \N__7912\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8720\,
            ce => 'H',
            sr => \N__10100\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001011110000"
        )
    port map (
            in0 => \N__6142\,
            in1 => \N__4197\,
            in2 => \N__4785\,
            in3 => \N__4721\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8720\,
            ce => 'H',
            sr => \N__10100\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6719\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8720\,
            ce => 'H',
            sr => \N__10100\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6737\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8720\,
            ce => 'H',
            sr => \N__10100\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4498\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7908\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8720\,
            ce => 'H',
            sr => \N__10100\
        );

    \U712_CHIP_RAM.REFRESH_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__4485\,
            in1 => \N__4467\,
            in2 => \N__4458\,
            in3 => \N__4437\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8724\,
            ce => 'H',
            sr => \N__10097\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__5054\,
            in1 => \N__9639\,
            in2 => \N__4428\,
            in3 => \N__4869\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8724\,
            ce => 'H',
            sr => \N__10097\
        );

    \U712_REG_SM.REG_TACK_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__4365\,
            in1 => \N__4371\,
            in2 => \N__4395\,
            in3 => \N__4380\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8727\,
            ce => 'H',
            sr => \N__10091\
        );

    \U712_REG_SM.STATE_COUNT_RNI4BRH_3_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4618\,
            in1 => \N__6550\,
            in2 => \_gnd_net_\,
            in3 => \N__6693\,
            lcout => \U712_REG_SM.N_225\,
            ltout => \U712_REG_SM.N_225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100010001"
        )
    port map (
            in0 => \N__7614\,
            in1 => \N__4629\,
            in2 => \N__4374\,
            in3 => \N__6498\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8731\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6692\,
            in1 => \N__6549\,
            in2 => \_gnd_net_\,
            in3 => \N__5191\,
            lcout => \U712_REG_SM.N_292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__5597\,
            in1 => \N__4601\,
            in2 => \N__6662\,
            in3 => \N__4617\,
            lcout => \U712_REG_SM.REG_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__4619\,
            in1 => \N__7617\,
            in2 => \_gnd_net_\,
            in3 => \N__6694\,
            lcout => OPEN,
            ltout => \U712_REG_SM.STATE_COUNT_srsts_i_i_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__6695\,
            in1 => \N__5192\,
            in2 => \N__4632\,
            in3 => \N__4961\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8731\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIEMV42_4_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6657\,
            in1 => \N__7616\,
            in2 => \_gnd_net_\,
            in3 => \N__5596\,
            lcout => \U712_REG_SM.N_289\,
            ltout => \U712_REG_SM.N_289_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__7615\,
            in1 => \N__5193\,
            in2 => \N__4623\,
            in3 => \N__4620\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8731\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011101"
        )
    port map (
            in0 => \N__4600\,
            in1 => \N__6653\,
            in2 => \_gnd_net_\,
            in3 => \N__6588\,
            lcout => \U712_REG_SM.DS_EN_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5905\,
            in1 => \N__4784\,
            in2 => \N__6150\,
            in3 => \N__4707\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_261_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4532\,
            in2 => \N__4551\,
            in3 => \N__4521\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8710\,
            ce => 'H',
            sr => \N__10116\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6012\,
            in1 => \N__6188\,
            in2 => \N__6149\,
            in3 => \N__5388\,
            lcout => \U712_CHIP_RAM.N_260\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIS6PC1_2_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5904\,
            in1 => \N__5816\,
            in2 => \_gnd_net_\,
            in3 => \N__5701\,
            lcout => \U712_CHIP_RAM.N_342\,
            ltout => \U712_CHIP_RAM.N_342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__5817\,
            in1 => \N__5706\,
            in2 => \N__4710\,
            in3 => \N__6011\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__5414\,
            in1 => \_gnd_net_\,
            in2 => \N__4647\,
            in3 => \N__6170\,
            lcout => \U712_CHIP_RAM.N_284\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI2B8VE_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__5337\,
            in1 => \N__4706\,
            in2 => \N__4836\,
            in3 => \N__4791\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_sbtinv_1_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4695\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__4692\,
            in1 => \N__5699\,
            in2 => \N__6013\,
            in3 => \N__6117\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__8821\,
            in1 => \N__5431\,
            in2 => \N__4686\,
            in3 => \N__5442\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4683\,
            in1 => \N__4665\,
            in2 => \_gnd_net_\,
            in3 => \N__8369\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100111111"
        )
    port map (
            in0 => \N__4782\,
            in1 => \N__5700\,
            in2 => \N__6134\,
            in3 => \N__5903\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER44_4_0_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNILL8G1_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5811\,
            in1 => \N__5698\,
            in2 => \N__5914\,
            in3 => \N__4781\,
            lcout => \U712_CHIP_RAM.N_270_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_1_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__7692\,
            in1 => \N__6300\,
            in2 => \N__5613\,
            in3 => \N__5454\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8713\,
            ce => \N__4815\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5468\,
            in1 => \N__5483\,
            in2 => \N__5502\,
            in3 => \N__6338\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_1_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5788\,
            in2 => \N__4809\,
            in3 => \N__5979\,
            lcout => \U712_CHIP_RAM.N_211\,
            ltout => \U712_CHIP_RAM.N_211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4806\,
            in2 => \N__4800\,
            in3 => \N__4932\,
            lcout => \U712_CHIP_RAM.N_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL6NI4_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5787\,
            in1 => \N__7693\,
            in2 => \N__5387\,
            in3 => \N__4947\,
            lcout => \U712_CHIP_RAM.N_266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001010000000"
        )
    port map (
            in0 => \N__5781\,
            in1 => \N__5670\,
            in2 => \N__6000\,
            in3 => \N__4766\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5869\,
            in1 => \N__6110\,
            in2 => \N__4746\,
            in3 => \N__5377\,
            lcout => \U712_CHIP_RAM.N_264\,
            ltout => \U712_CHIP_RAM.N_264_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHUFGC_0_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__7662\,
            in1 => \N__4938\,
            in2 => \N__4728\,
            in3 => \N__4919\,
            lcout => \U712_CHIP_RAM.N_36\,
            ltout => \U712_CHIP_RAM.N_36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__5410\,
            in1 => \N__5517\,
            in2 => \N__4725\,
            in3 => \N__4722\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8716\,
            ce => \N__6327\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_1_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000100000"
        )
    port map (
            in0 => \N__6109\,
            in1 => \N__5669\,
            in2 => \N__5999\,
            in3 => \N__5868\,
            lcout => \U712_CHIP_RAM.N_209\,
            ltout => \U712_CHIP_RAM.N_209_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_0_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5782\,
            in2 => \N__4941\,
            in3 => \N__5378\,
            lcout => \U712_CHIP_RAM.N_263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__6201\,
            in1 => \N__6369\,
            in2 => \N__4926\,
            in3 => \N__5529\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8716\,
            ce => \N__6327\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100011"
        )
    port map (
            in0 => \N__5671\,
            in1 => \N__5783\,
            in2 => \N__5899\,
            in3 => \N__5978\,
            lcout => \U712_CHIP_RAM.N_246\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNILCLN6_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__4855\,
            in1 => \N__4824\,
            in2 => \N__5415\,
            in3 => \N__4918\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_SYNC_RNI5J861_1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100111111"
        )
    port map (
            in0 => \N__5069\,
            in1 => \N__4868\,
            in2 => \N__4994\,
            in3 => \N__5088\,
            lcout => \U712_CHIP_RAM.N_203\,
            ltout => \U712_CHIP_RAM.N_203_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIH0703_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7661\,
            in1 => \N__4823\,
            in2 => \N__4839\,
            in3 => \N__6083\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__9513\,
            in1 => \N__5001\,
            in2 => \N__6242\,
            in3 => \N__7119\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8721\,
            ce => 'H',
            sr => \N__10092\
        );

    \U712_CHIP_RAM.REFRESH_RNIRILU_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6276\,
            in2 => \_gnd_net_\,
            in3 => \N__6226\,
            lcout => \U712_CHIP_RAM.N_341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_SYNC_1_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5070\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8721\,
            ce => 'H',
            sr => \N__10092\
        );

    \U712_CHIP_RAM.REFRESH_SYNC_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5082\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9162\,
            lcout => \U712_CHIP_RAM.REFRESH_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8721\,
            ce => 'H',
            sr => \N__10092\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001101"
        )
    port map (
            in0 => \N__5061\,
            in1 => \N__5178\,
            in2 => \N__5025\,
            in3 => \N__8512\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8725\,
            ce => 'H',
            sr => \N__10086\
        );

    \DBR_SYNC_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7811\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8725\,
            ce => 'H',
            sr => \N__10086\
        );

    \DBR_SYNC_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4977\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8725\,
            ce => 'H',
            sr => \N__10086\
        );

    \U712_CHIP_RAM.CAS_SYNC_2_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8538\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8725\,
            ce => 'H',
            sr => \N__10086\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__6696\,
            in1 => \N__7612\,
            in2 => \N__4962\,
            in3 => \N__7085\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8728\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI07K21_1_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__6586\,
            in1 => \N__6623\,
            in2 => \N__4995\,
            in3 => \N__4976\,
            lcout => OPEN,
            ltout => \U712_REG_SM.STATE_COUNT_srsts_i_i_0_o2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI35EO1_1_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__5582\,
            in1 => \_gnd_net_\,
            in2 => \N__4965\,
            in3 => \N__5560\,
            lcout => \U712_REG_SM.N_245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIAS4F1_0_1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__6585\,
            in1 => \N__5559\,
            in2 => \N__6627\,
            in3 => \N__5580\,
            lcout => \U712_REG_SM.N_215\,
            ltout => \U712_REG_SM.N_215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNITO6S1_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5177\,
            in2 => \N__5166\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.N_228\,
            ltout => \U712_REG_SM.N_228_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111110111"
        )
    port map (
            in0 => \N__7613\,
            in1 => \N__6479\,
            in2 => \N__5163\,
            in3 => \N__6554\,
            lcout => OPEN,
            ltout => \U712_REG_SM.STATE_COUNT_srsts_i_i_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__6624\,
            in1 => \N__6587\,
            in2 => \N__5160\,
            in3 => \N__7749\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8728\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNIAS4F1_1_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__6584\,
            in1 => \N__5558\,
            in2 => \N__6626\,
            in3 => \N__5581\,
            lcout => \U712_REG_SM.N_210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5157\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8732\,
            ce => 'H',
            sr => \N__10081\
        );

    \U712_REG_SM.C1_SYNC_1_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5562\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8732\,
            ce => 'H',
            sr => \N__10081\
        );

    \U712_REG_SM.C3_SYNC_1_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6591\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8732\,
            ce => 'H',
            sr => \N__10081\
        );

    \U712_REG_SM.C3_SYNC_0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5124\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8732\,
            ce => 'H',
            sr => \N__10081\
        );

    \U712_REG_SM.REG_CYCLE_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6464\,
            in1 => \N__7696\,
            in2 => \_gnd_net_\,
            in3 => \N__7789\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8893\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_0_3_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8813\,
            in1 => \N__7530\,
            in2 => \N__8269\,
            in3 => \N__8396\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5262\,
            in1 => \N__5241\,
            in2 => \_gnd_net_\,
            in3 => \N__8397\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5229\,
            in1 => \N__9688\,
            in2 => \_gnd_net_\,
            in3 => \N__8577\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__7336\,
            in1 => \_gnd_net_\,
            in2 => \N__5208\,
            in3 => \N__8398\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNITDMK_3_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111101"
        )
    port map (
            in0 => \N__8270\,
            in1 => \N__7532\,
            in2 => \N__8399\,
            in3 => \N__8814\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI9CFE_0_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__7533\,
            in1 => \N__8360\,
            in2 => \_gnd_net_\,
            in3 => \N__8271\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101101110"
        )
    port map (
            in0 => \N__5705\,
            in1 => \N__6132\,
            in2 => \N__6014\,
            in3 => \N__5906\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5386\,
            in1 => \N__7694\,
            in2 => \N__5205\,
            in3 => \N__5812\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001011"
        )
    port map (
            in0 => \N__8272\,
            in1 => \N__5432\,
            in2 => \N__5202\,
            in3 => \N__5199\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9683\,
            in1 => \N__5280\,
            in2 => \N__8430\,
            in3 => \N__7941\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIISK15_2_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__7695\,
            in1 => \N__5535\,
            in2 => \_gnd_net_\,
            in3 => \N__5453\,
            lcout => \U712_CHIP_RAM.N_64_1\,
            ltout => \U712_CHIP_RAM.N_64_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111011000"
        )
    port map (
            in0 => \N__5433\,
            in1 => \N__7540\,
            in2 => \N__5418\,
            in3 => \N__5328\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8711\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7685\,
            in2 => \_gnd_net_\,
            in3 => \N__6106\,
            lcout => \U712_CHIP_RAM.N_340\,
            ltout => \U712_CHIP_RAM.N_340_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOGP34_3_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5886\,
            in1 => \N__5321\,
            in2 => \N__5391\,
            in3 => \N__5376\,
            lcout => \U712_CHIP_RAM.N_267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5890\,
            in1 => \N__5790\,
            in2 => \_gnd_net_\,
            in3 => \N__5971\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_281_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__5322\,
            in1 => \_gnd_net_\,
            in2 => \N__5331\,
            in3 => \N__6108\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_102_i_a2_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5667\,
            in2 => \_gnd_net_\,
            in3 => \N__5970\,
            lcout => \U712_CHIP_RAM.N_207_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5313\,
            in1 => \N__5295\,
            in2 => \_gnd_net_\,
            in3 => \N__8368\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNINN5O1_2_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100011100"
        )
    port map (
            in0 => \N__6107\,
            in1 => \N__5789\,
            in2 => \N__5907\,
            in3 => \N__5668\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_141_i_a2_0_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5794\,
            in2 => \_gnd_net_\,
            in3 => \N__5523\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \bfn_10_8_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6370\,
            in1 => \N__5981\,
            in2 => \_gnd_net_\,
            in3 => \N__5520\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__8714\,
            ce => \N__6323\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5695\,
            in2 => \_gnd_net_\,
            in3 => \N__5508\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6371\,
            in1 => \N__5894\,
            in2 => \_gnd_net_\,
            in3 => \N__5505\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__8714\,
            ce => \N__6323\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6366\,
            in1 => \N__5501\,
            in2 => \_gnd_net_\,
            in3 => \N__5487\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__8714\,
            ce => \N__6323\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6372\,
            in1 => \N__5484\,
            in2 => \_gnd_net_\,
            in3 => \N__5472\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__8714\,
            ce => \N__6323\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__6367\,
            in1 => \N__5469\,
            in2 => \_gnd_net_\,
            in3 => \N__5457\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__8714\,
            ce => \N__6323\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__6339\,
            in1 => \N__6368\,
            in2 => \_gnd_net_\,
            in3 => \N__6342\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8714\,
            ce => \N__6323\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_0_1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100000000"
        )
    port map (
            in0 => \N__5793\,
            in1 => \N__6290\,
            in2 => \N__6252\,
            in3 => \N__6091\,
            lcout => \U712_CHIP_RAM.N_285\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010001010"
        )
    port map (
            in0 => \N__7663\,
            in1 => \N__6291\,
            in2 => \N__6122\,
            in3 => \N__6241\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_0_a3_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__6195\,
            in1 => \N__6095\,
            in2 => \_gnd_net_\,
            in3 => \N__6177\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8717\,
            ce => 'H',
            sr => \N__10087\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_2_1_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000010001"
        )
    port map (
            in0 => \N__5791\,
            in1 => \N__6090\,
            in2 => \_gnd_net_\,
            in3 => \N__5980\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_2_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNO_1_1_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110110"
        )
    port map (
            in0 => \N__5898\,
            in1 => \N__5792\,
            in2 => \N__5709\,
            in3 => \N__5694\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_62_i_a2_2_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIOC3L1_4_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__6658\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5598\,
            lcout => \U712_REG_SM.ASn_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_3_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111101110"
        )
    port map (
            in0 => \N__6690\,
            in1 => \N__6622\,
            in2 => \_gnd_net_\,
            in3 => \N__6589\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_248_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_2_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110101"
        )
    port map (
            in0 => \N__6547\,
            in1 => \N__5583\,
            in2 => \N__5565\,
            in3 => \N__5561\,
            lcout => \U712_REG_SM.un1_ASn_0_sqmuxa_1_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__6691\,
            in1 => \N__6548\,
            in2 => \N__6663\,
            in3 => \N__7747\,
            lcout => \U712_REG_SM.N_300\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIBMB91_1_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__6625\,
            in1 => \N__6590\,
            in2 => \N__6555\,
            in3 => \N__7746\,
            lcout => \U712_REG_SM.N_226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001011"
        )
    port map (
            in0 => \N__10307\,
            in1 => \N__6522\,
            in2 => \N__6516\,
            in3 => \N__6504\,
            lcout => \DS_ENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8729\,
            ce => 'H',
            sr => \N__10078\
        );

    \U712_REG_SM.REGENn_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110101011111010"
        )
    port map (
            in0 => \N__7098\,
            in1 => \N__6497\,
            in2 => \N__6460\,
            in3 => \N__6486\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8729\,
            ce => 'H',
            sr => \N__10078\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__7203\,
            in1 => \N__8121\,
            in2 => \N__7359\,
            in3 => \N__6432\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8701\,
            ce => \N__7385\,
            sr => \N__10111\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIJNI41_3_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10138\,
            in2 => \_gnd_net_\,
            in3 => \N__6411\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9705\,
            in1 => \N__6405\,
            in2 => \N__8457\,
            in3 => \N__7929\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7293\,
            in1 => \N__6399\,
            in2 => \_gnd_net_\,
            in3 => \N__6777\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8706\,
            ce => \N__7386\,
            sr => \N__10098\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7531\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8255\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6819\,
            in1 => \N__6744\,
            in2 => \_gnd_net_\,
            in3 => \N__6885\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8706\,
            ce => \N__7386\,
            sr => \N__10098\
        );

    \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5_1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8405\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9640\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_e_0_RNIR4H5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6858\,
            in1 => \N__6840\,
            in2 => \_gnd_net_\,
            in3 => \N__8404\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__7467\,
            in1 => \N__8132\,
            in2 => \N__9684\,
            in3 => \N__6767\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6813\,
            in1 => \N__6795\,
            in2 => \_gnd_net_\,
            in3 => \N__8406\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8407\,
            in1 => \N__9641\,
            in2 => \N__6780\,
            in3 => \N__7953\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011111111"
        )
    port map (
            in0 => \N__8133\,
            in1 => \N__9642\,
            in2 => \N__6771\,
            in3 => \N__7468\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6738\,
            in2 => \_gnd_net_\,
            in3 => \N__6720\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__7055\,
            in1 => \N__7097\,
            in2 => \_gnd_net_\,
            in3 => \N__7086\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8722\,
            ce => 'H',
            sr => \N__10079\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7550\,
            in1 => \N__8459\,
            in2 => \N__8835\,
            in3 => \N__8279\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8697\,
            ce => \N__7407\,
            sr => \N__10108\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__7204\,
            in1 => \N__7284\,
            in2 => \N__7356\,
            in3 => \N__6900\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8700\,
            ce => \N__7387\,
            sr => \N__10095\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__6996\,
            in1 => \N__7481\,
            in2 => \N__9722\,
            in3 => \N__9174\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8700\,
            ce => \N__7387\,
            sr => \N__10095\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__7205\,
            in1 => \N__9234\,
            in2 => \N__7357\,
            in3 => \N__6960\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8700\,
            ce => \N__7387\,
            sr => \N__10095\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__8103\,
            in1 => \N__7348\,
            in2 => \N__7209\,
            in3 => \N__7254\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8700\,
            ce => \N__7387\,
            sr => \N__10095\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9696\,
            in1 => \N__6906\,
            in2 => \N__8460\,
            in3 => \N__7992\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9697\,
            in1 => \N__6894\,
            in2 => \N__8461\,
            in3 => \N__8619\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9698\,
            in1 => \N__7248\,
            in2 => \N__8462\,
            in3 => \N__7146\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9646\,
            in1 => \N__7239\,
            in2 => \N__8458\,
            in3 => \N__8625\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__7191\,
            in1 => \N__7346\,
            in2 => \N__7227\,
            in3 => \N__8109\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8705\,
            ce => \N__7403\,
            sr => \N__10085\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__7192\,
            in1 => \N__7347\,
            in2 => \N__8094\,
            in3 => \N__7173\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8705\,
            ce => \N__7403\,
            sr => \N__10085\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8961\,
            in1 => \N__9125\,
            in2 => \_gnd_net_\,
            in3 => \N__9222\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__8561\,
            sr => \N__10083\
        );

    \U712_CHIP_RAM.DMA_A20_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__9099\,
            in1 => \N__7104\,
            in2 => \N__8960\,
            in3 => \N__7133\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10080\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8534\,
            in2 => \_gnd_net_\,
            in3 => \N__8750\,
            lcout => \U712_CHIP_RAM.un5_DMA_CYCLE_START_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS10_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7804\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8901\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10\,
            ltout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_ctle_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7917\,
            in3 => \N__10137\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_RNI8MQ3_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7913\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__10136\,
            in1 => \N__7812\,
            in2 => \_gnd_net_\,
            in3 => \N__7748\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7657\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RASn_LC_13_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7551\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8698\,
            ce => 'H',
            sr => \N__10117\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__7482\,
            in1 => \N__7449\,
            in2 => \N__9723\,
            in3 => \N__8913\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8703\,
            ce => \N__7396\,
            sr => \N__10101\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011110000"
        )
    port map (
            in0 => \N__9695\,
            in1 => \N__7265\,
            in2 => \N__7358\,
            in3 => \N__8443\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9100\,
            in1 => \N__8027\,
            in2 => \_gnd_net_\,
            in3 => \N__8082\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8895\,
            ce => \N__8866\,
            sr => \N__10093\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8028\,
            in1 => \N__9101\,
            in2 => \_gnd_net_\,
            in3 => \N__7982\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8895\,
            ce => \N__8866\,
            sr => \N__10093\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__7983\,
            in1 => \N__9276\,
            in2 => \N__9122\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8895\,
            ce => \N__8866\,
            sr => \N__10093\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__8208\,
            in1 => \_gnd_net_\,
            in2 => \N__9123\,
            in3 => \N__9330\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8895\,
            ce => \N__8866\,
            sr => \N__10093\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__8172\,
            in1 => \_gnd_net_\,
            in2 => \N__9124\,
            in3 => \N__8609\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8895\,
            ce => \N__8866\,
            sr => \N__10093\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8610\,
            in1 => \N__9221\,
            in2 => \_gnd_net_\,
            in3 => \N__9111\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8895\,
            ce => \N__8866\,
            sr => \N__10093\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8081\,
            in1 => \N__9084\,
            in2 => \_gnd_net_\,
            in3 => \N__8020\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__8565\,
            sr => \N__10088\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__8021\,
            in1 => \_gnd_net_\,
            in2 => \N__9118\,
            in3 => \N__7980\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__8565\,
            sr => \N__10088\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7981\,
            in1 => \N__9088\,
            in2 => \_gnd_net_\,
            in3 => \N__9271\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__8565\,
            sr => \N__10088\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9272\,
            in1 => \_gnd_net_\,
            in2 => \N__9119\,
            in3 => \N__9328\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__8565\,
            sr => \N__10088\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9329\,
            in1 => \N__9092\,
            in2 => \_gnd_net_\,
            in3 => \N__8205\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__8565\,
            sr => \N__10088\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__8168\,
            in1 => \_gnd_net_\,
            in2 => \N__9120\,
            in3 => \N__8206\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__8565\,
            sr => \N__10088\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__9220\,
            in1 => \_gnd_net_\,
            in2 => \N__9121\,
            in3 => \N__8608\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__8565\,
            sr => \N__10088\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8167\,
            in1 => \N__9040\,
            in2 => \_gnd_net_\,
            in3 => \N__8607\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__8557\,
            sr => \N__10084\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8751\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8718\,
            ce => 'H',
            sr => \N__10082\
        );

    \U712_BUFFERS.un1_DRDENn_0_a3_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9522\,
            in2 => \_gnd_net_\,
            in3 => \N__8519\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_14_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8466\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8699\,
            ce => 'H',
            sr => \N__10119\
        );

    \U712_CHIP_RAM.WEn_LC_14_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8280\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8702\,
            ce => 'H',
            sr => \N__10118\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8207\,
            in1 => \N__9076\,
            in2 => \_gnd_net_\,
            in3 => \N__8166\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8897\,
            ce => \N__8870\,
            sr => \N__10099\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9324\,
            in1 => \N__9041\,
            in2 => \_gnd_net_\,
            in3 => \N__9257\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8896\,
            ce => \N__8871\,
            sr => \N__10094\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9210\,
            in1 => \_gnd_net_\,
            in2 => \N__9083\,
            in3 => \N__8947\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8896\,
            ce => \N__8871\,
            sr => \N__10094\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9158\,
            in1 => \N__9014\,
            in2 => \_gnd_net_\,
            in3 => \N__8946\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8894\,
            ce => \N__8856\,
            sr => \N__10089\
        );

    \U712_CHIP_RAM.CRCSn_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8834\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8704\,
            ce => 'H',
            sr => \N__10120\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_a3_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__10292\,
            in1 => \_gnd_net_\,
            in2 => \N__9770\,
            in3 => \N__9725\,
            lcout => \U712_BYTE_ENABLE.N_313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a3_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__9724\,
            in1 => \N__9762\,
            in2 => \N__9875\,
            in3 => \N__10291\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_315_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__9374\,
            in1 => \N__9987\,
            in2 => \N__8769\,
            in3 => \N__9514\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9449\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9982\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__8726\,
            ce => 'H',
            sr => \N__10090\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__9392\,
            in1 => \N__9945\,
            in2 => \N__9986\,
            in3 => \N__9528\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a3_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__10286\,
            in1 => \N__9766\,
            in2 => \N__9876\,
            in3 => \N__9718\,
            lcout => \U712_BYTE_ENABLE.N_311\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_0_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__9939\,
            in1 => \N__9450\,
            in2 => \N__9524\,
            in3 => \N__9375\,
            lcout => \U712_BYTE_ENABLE.un1_CLMBEn_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__10200\,
            in1 => \N__10274\,
            in2 => \_gnd_net_\,
            in3 => \N__10319\,
            lcout => \N_170\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_174_i_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101000101"
        )
    port map (
            in0 => \N__9915\,
            in1 => \N__9879\,
            in2 => \N__9726\,
            in3 => \N__10231\,
            lcout => \N_174_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_172_i_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000110011"
        )
    port map (
            in0 => \N__9877\,
            in1 => \N__9336\,
            in2 => \N__10232\,
            in3 => \N__9647\,
            lcout => \N_172_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_176_i_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000110011"
        )
    port map (
            in0 => \N__9878\,
            in1 => \N__9801\,
            in2 => \N__10233\,
            in3 => \N__9648\,
            lcout => \N_176_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_a3_0_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__9774\,
            in1 => \N__10296\,
            in2 => \_gnd_net_\,
            in3 => \N__9709\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_309_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110000"
        )
    port map (
            in0 => \N__9518\,
            in1 => \N__9442\,
            in2 => \N__9399\,
            in3 => \N__9385\,
            lcout => \U712_BYTE_ENABLE.un1_CUUBEn_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_UDSn_i_0_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__10320\,
            in1 => \N__10287\,
            in2 => \_gnd_net_\,
            in3 => \N__10216\,
            lcout => \N_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

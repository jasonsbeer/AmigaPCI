// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 8 2025 19:54:41

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    DRA,
    CMA,
    DA,
    A,
    DBRn,
    RAMENn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    TCIn,
    TBIn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    input [9:0] DRA;
    output [10:0] CMA;
    output [2:0] DA;
    input [20:0] A;
    input DBRn;
    output RAMENn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    output TCIn;
    output TBIn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__12194;
    wire N__12193;
    wire N__12192;
    wire N__12185;
    wire N__12184;
    wire N__12183;
    wire N__12176;
    wire N__12175;
    wire N__12174;
    wire N__12167;
    wire N__12166;
    wire N__12165;
    wire N__12158;
    wire N__12157;
    wire N__12156;
    wire N__12149;
    wire N__12148;
    wire N__12147;
    wire N__12140;
    wire N__12139;
    wire N__12138;
    wire N__12131;
    wire N__12130;
    wire N__12129;
    wire N__12122;
    wire N__12121;
    wire N__12120;
    wire N__12113;
    wire N__12112;
    wire N__12111;
    wire N__12104;
    wire N__12103;
    wire N__12102;
    wire N__12095;
    wire N__12094;
    wire N__12093;
    wire N__12086;
    wire N__12085;
    wire N__12084;
    wire N__12077;
    wire N__12076;
    wire N__12075;
    wire N__12068;
    wire N__12067;
    wire N__12066;
    wire N__12059;
    wire N__12058;
    wire N__12057;
    wire N__12050;
    wire N__12049;
    wire N__12048;
    wire N__12041;
    wire N__12040;
    wire N__12039;
    wire N__12032;
    wire N__12031;
    wire N__12030;
    wire N__12023;
    wire N__12022;
    wire N__12021;
    wire N__12014;
    wire N__12013;
    wire N__12012;
    wire N__12005;
    wire N__12004;
    wire N__12003;
    wire N__11996;
    wire N__11995;
    wire N__11994;
    wire N__11987;
    wire N__11986;
    wire N__11985;
    wire N__11978;
    wire N__11977;
    wire N__11976;
    wire N__11969;
    wire N__11968;
    wire N__11967;
    wire N__11960;
    wire N__11959;
    wire N__11958;
    wire N__11951;
    wire N__11950;
    wire N__11949;
    wire N__11942;
    wire N__11941;
    wire N__11940;
    wire N__11933;
    wire N__11932;
    wire N__11931;
    wire N__11924;
    wire N__11923;
    wire N__11922;
    wire N__11915;
    wire N__11914;
    wire N__11913;
    wire N__11906;
    wire N__11905;
    wire N__11904;
    wire N__11897;
    wire N__11896;
    wire N__11895;
    wire N__11888;
    wire N__11887;
    wire N__11886;
    wire N__11879;
    wire N__11878;
    wire N__11877;
    wire N__11870;
    wire N__11869;
    wire N__11868;
    wire N__11861;
    wire N__11860;
    wire N__11859;
    wire N__11852;
    wire N__11851;
    wire N__11850;
    wire N__11843;
    wire N__11842;
    wire N__11841;
    wire N__11834;
    wire N__11833;
    wire N__11832;
    wire N__11825;
    wire N__11824;
    wire N__11823;
    wire N__11816;
    wire N__11815;
    wire N__11814;
    wire N__11807;
    wire N__11806;
    wire N__11805;
    wire N__11798;
    wire N__11797;
    wire N__11796;
    wire N__11789;
    wire N__11788;
    wire N__11787;
    wire N__11780;
    wire N__11779;
    wire N__11778;
    wire N__11771;
    wire N__11770;
    wire N__11769;
    wire N__11762;
    wire N__11761;
    wire N__11760;
    wire N__11753;
    wire N__11752;
    wire N__11751;
    wire N__11744;
    wire N__11743;
    wire N__11742;
    wire N__11735;
    wire N__11734;
    wire N__11733;
    wire N__11726;
    wire N__11725;
    wire N__11724;
    wire N__11717;
    wire N__11716;
    wire N__11715;
    wire N__11708;
    wire N__11707;
    wire N__11706;
    wire N__11699;
    wire N__11698;
    wire N__11697;
    wire N__11690;
    wire N__11689;
    wire N__11688;
    wire N__11681;
    wire N__11680;
    wire N__11679;
    wire N__11672;
    wire N__11671;
    wire N__11670;
    wire N__11663;
    wire N__11662;
    wire N__11661;
    wire N__11654;
    wire N__11653;
    wire N__11652;
    wire N__11645;
    wire N__11644;
    wire N__11643;
    wire N__11636;
    wire N__11635;
    wire N__11634;
    wire N__11627;
    wire N__11626;
    wire N__11625;
    wire N__11618;
    wire N__11617;
    wire N__11616;
    wire N__11609;
    wire N__11608;
    wire N__11607;
    wire N__11600;
    wire N__11599;
    wire N__11598;
    wire N__11591;
    wire N__11590;
    wire N__11589;
    wire N__11582;
    wire N__11581;
    wire N__11580;
    wire N__11573;
    wire N__11572;
    wire N__11571;
    wire N__11564;
    wire N__11563;
    wire N__11562;
    wire N__11555;
    wire N__11554;
    wire N__11553;
    wire N__11546;
    wire N__11545;
    wire N__11544;
    wire N__11537;
    wire N__11536;
    wire N__11535;
    wire N__11528;
    wire N__11527;
    wire N__11526;
    wire N__11519;
    wire N__11518;
    wire N__11517;
    wire N__11510;
    wire N__11509;
    wire N__11508;
    wire N__11501;
    wire N__11500;
    wire N__11499;
    wire N__11492;
    wire N__11491;
    wire N__11490;
    wire N__11483;
    wire N__11482;
    wire N__11481;
    wire N__11474;
    wire N__11473;
    wire N__11472;
    wire N__11465;
    wire N__11464;
    wire N__11463;
    wire N__11456;
    wire N__11455;
    wire N__11454;
    wire N__11447;
    wire N__11446;
    wire N__11445;
    wire N__11438;
    wire N__11437;
    wire N__11436;
    wire N__11429;
    wire N__11428;
    wire N__11427;
    wire N__11420;
    wire N__11419;
    wire N__11418;
    wire N__11411;
    wire N__11410;
    wire N__11409;
    wire N__11402;
    wire N__11401;
    wire N__11400;
    wire N__11393;
    wire N__11392;
    wire N__11391;
    wire N__11384;
    wire N__11383;
    wire N__11382;
    wire N__11375;
    wire N__11374;
    wire N__11373;
    wire N__11366;
    wire N__11365;
    wire N__11364;
    wire N__11357;
    wire N__11356;
    wire N__11355;
    wire N__11348;
    wire N__11347;
    wire N__11346;
    wire N__11329;
    wire N__11326;
    wire N__11325;
    wire N__11324;
    wire N__11321;
    wire N__11320;
    wire N__11317;
    wire N__11316;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11304;
    wire N__11301;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11289;
    wire N__11286;
    wire N__11283;
    wire N__11280;
    wire N__11275;
    wire N__11270;
    wire N__11267;
    wire N__11262;
    wire N__11257;
    wire N__11256;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11245;
    wire N__11242;
    wire N__11237;
    wire N__11234;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11224;
    wire N__11219;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11201;
    wire N__11196;
    wire N__11193;
    wire N__11190;
    wire N__11187;
    wire N__11184;
    wire N__11179;
    wire N__11176;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11157;
    wire N__11156;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11146;
    wire N__11143;
    wire N__11138;
    wire N__11133;
    wire N__11130;
    wire N__11127;
    wire N__11122;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11110;
    wire N__11107;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11095;
    wire N__11092;
    wire N__11089;
    wire N__11088;
    wire N__11087;
    wire N__11086;
    wire N__11085;
    wire N__11084;
    wire N__11083;
    wire N__11076;
    wire N__11071;
    wire N__11066;
    wire N__11065;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11053;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11026;
    wire N__11023;
    wire N__11020;
    wire N__11019;
    wire N__11018;
    wire N__11013;
    wire N__11012;
    wire N__11011;
    wire N__11010;
    wire N__11007;
    wire N__11006;
    wire N__11005;
    wire N__11002;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10966;
    wire N__10961;
    wire N__10958;
    wire N__10953;
    wire N__10950;
    wire N__10947;
    wire N__10942;
    wire N__10941;
    wire N__10940;
    wire N__10937;
    wire N__10936;
    wire N__10933;
    wire N__10930;
    wire N__10929;
    wire N__10928;
    wire N__10927;
    wire N__10924;
    wire N__10917;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10902;
    wire N__10897;
    wire N__10894;
    wire N__10885;
    wire N__10882;
    wire N__10879;
    wire N__10876;
    wire N__10873;
    wire N__10870;
    wire N__10869;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10858;
    wire N__10857;
    wire N__10854;
    wire N__10851;
    wire N__10844;
    wire N__10843;
    wire N__10842;
    wire N__10841;
    wire N__10836;
    wire N__10833;
    wire N__10828;
    wire N__10825;
    wire N__10822;
    wire N__10815;
    wire N__10812;
    wire N__10809;
    wire N__10804;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10789;
    wire N__10786;
    wire N__10785;
    wire N__10782;
    wire N__10779;
    wire N__10778;
    wire N__10773;
    wire N__10770;
    wire N__10769;
    wire N__10764;
    wire N__10761;
    wire N__10758;
    wire N__10755;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10731;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10720;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10701;
    wire N__10698;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10684;
    wire N__10681;
    wire N__10678;
    wire N__10675;
    wire N__10674;
    wire N__10673;
    wire N__10668;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10641;
    wire N__10638;
    wire N__10635;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10617;
    wire N__10616;
    wire N__10615;
    wire N__10614;
    wire N__10613;
    wire N__10606;
    wire N__10603;
    wire N__10600;
    wire N__10599;
    wire N__10598;
    wire N__10597;
    wire N__10596;
    wire N__10595;
    wire N__10594;
    wire N__10593;
    wire N__10592;
    wire N__10591;
    wire N__10588;
    wire N__10587;
    wire N__10584;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10569;
    wire N__10562;
    wire N__10559;
    wire N__10556;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10535;
    wire N__10532;
    wire N__10531;
    wire N__10530;
    wire N__10527;
    wire N__10522;
    wire N__10521;
    wire N__10518;
    wire N__10515;
    wire N__10512;
    wire N__10509;
    wire N__10506;
    wire N__10503;
    wire N__10498;
    wire N__10493;
    wire N__10490;
    wire N__10485;
    wire N__10480;
    wire N__10475;
    wire N__10468;
    wire N__10465;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10446;
    wire N__10443;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10404;
    wire N__10403;
    wire N__10398;
    wire N__10395;
    wire N__10392;
    wire N__10389;
    wire N__10386;
    wire N__10383;
    wire N__10380;
    wire N__10377;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10363;
    wire N__10360;
    wire N__10357;
    wire N__10356;
    wire N__10355;
    wire N__10354;
    wire N__10353;
    wire N__10352;
    wire N__10351;
    wire N__10350;
    wire N__10333;
    wire N__10330;
    wire N__10327;
    wire N__10326;
    wire N__10325;
    wire N__10324;
    wire N__10323;
    wire N__10322;
    wire N__10321;
    wire N__10320;
    wire N__10319;
    wire N__10318;
    wire N__10317;
    wire N__10316;
    wire N__10315;
    wire N__10314;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10278;
    wire N__10277;
    wire N__10276;
    wire N__10275;
    wire N__10272;
    wire N__10269;
    wire N__10266;
    wire N__10261;
    wire N__10260;
    wire N__10259;
    wire N__10258;
    wire N__10257;
    wire N__10256;
    wire N__10255;
    wire N__10254;
    wire N__10253;
    wire N__10252;
    wire N__10251;
    wire N__10250;
    wire N__10247;
    wire N__10246;
    wire N__10245;
    wire N__10244;
    wire N__10243;
    wire N__10240;
    wire N__10239;
    wire N__10238;
    wire N__10237;
    wire N__10236;
    wire N__10235;
    wire N__10234;
    wire N__10233;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10225;
    wire N__10224;
    wire N__10223;
    wire N__10222;
    wire N__10221;
    wire N__10220;
    wire N__10219;
    wire N__10218;
    wire N__10217;
    wire N__10216;
    wire N__10215;
    wire N__10214;
    wire N__10213;
    wire N__10132;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10119;
    wire N__10116;
    wire N__10113;
    wire N__10110;
    wire N__10107;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10090;
    wire N__10087;
    wire N__10084;
    wire N__10081;
    wire N__10080;
    wire N__10077;
    wire N__10074;
    wire N__10069;
    wire N__10068;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10050;
    wire N__10045;
    wire N__10042;
    wire N__10039;
    wire N__10038;
    wire N__10033;
    wire N__10030;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10020;
    wire N__10019;
    wire N__10018;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10002;
    wire N__9999;
    wire N__9996;
    wire N__9993;
    wire N__9990;
    wire N__9987;
    wire N__9984;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9967;
    wire N__9964;
    wire N__9961;
    wire N__9958;
    wire N__9955;
    wire N__9954;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9946;
    wire N__9943;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9925;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9913;
    wire N__9910;
    wire N__9909;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9880;
    wire N__9877;
    wire N__9874;
    wire N__9871;
    wire N__9868;
    wire N__9865;
    wire N__9862;
    wire N__9859;
    wire N__9856;
    wire N__9853;
    wire N__9850;
    wire N__9849;
    wire N__9846;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9835;
    wire N__9834;
    wire N__9831;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9809;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9796;
    wire N__9787;
    wire N__9784;
    wire N__9783;
    wire N__9782;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9774;
    wire N__9771;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9743;
    wire N__9740;
    wire N__9739;
    wire N__9738;
    wire N__9735;
    wire N__9732;
    wire N__9729;
    wire N__9726;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9707;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9670;
    wire N__9667;
    wire N__9666;
    wire N__9665;
    wire N__9664;
    wire N__9663;
    wire N__9660;
    wire N__9659;
    wire N__9658;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9648;
    wire N__9645;
    wire N__9644;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9636;
    wire N__9635;
    wire N__9634;
    wire N__9633;
    wire N__9630;
    wire N__9629;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9621;
    wire N__9620;
    wire N__9617;
    wire N__9616;
    wire N__9613;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9592;
    wire N__9589;
    wire N__9586;
    wire N__9585;
    wire N__9580;
    wire N__9579;
    wire N__9578;
    wire N__9577;
    wire N__9572;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9556;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9535;
    wire N__9532;
    wire N__9527;
    wire N__9520;
    wire N__9513;
    wire N__9506;
    wire N__9501;
    wire N__9490;
    wire N__9487;
    wire N__9484;
    wire N__9481;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9469;
    wire N__9466;
    wire N__9463;
    wire N__9460;
    wire N__9457;
    wire N__9456;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9448;
    wire N__9445;
    wire N__9440;
    wire N__9437;
    wire N__9430;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9412;
    wire N__9409;
    wire N__9408;
    wire N__9407;
    wire N__9402;
    wire N__9399;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9389;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9339;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9313;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9292;
    wire N__9289;
    wire N__9286;
    wire N__9285;
    wire N__9282;
    wire N__9279;
    wire N__9274;
    wire N__9271;
    wire N__9270;
    wire N__9267;
    wire N__9264;
    wire N__9261;
    wire N__9256;
    wire N__9253;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9202;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9161;
    wire N__9160;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9148;
    wire N__9147;
    wire N__9144;
    wire N__9141;
    wire N__9138;
    wire N__9133;
    wire N__9130;
    wire N__9123;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9094;
    wire N__9091;
    wire N__9088;
    wire N__9087;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9076;
    wire N__9075;
    wire N__9074;
    wire N__9073;
    wire N__9072;
    wire N__9071;
    wire N__9070;
    wire N__9069;
    wire N__9068;
    wire N__9065;
    wire N__9062;
    wire N__9059;
    wire N__9052;
    wire N__9051;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9039;
    wire N__9036;
    wire N__9035;
    wire N__9032;
    wire N__9023;
    wire N__9022;
    wire N__9021;
    wire N__9016;
    wire N__9011;
    wire N__9006;
    wire N__9005;
    wire N__9004;
    wire N__9003;
    wire N__9002;
    wire N__9001;
    wire N__8998;
    wire N__8997;
    wire N__8996;
    wire N__8991;
    wire N__8988;
    wire N__8985;
    wire N__8982;
    wire N__8977;
    wire N__8970;
    wire N__8967;
    wire N__8964;
    wire N__8961;
    wire N__8956;
    wire N__8951;
    wire N__8942;
    wire N__8929;
    wire N__8928;
    wire N__8927;
    wire N__8926;
    wire N__8923;
    wire N__8922;
    wire N__8921;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8905;
    wire N__8902;
    wire N__8893;
    wire N__8892;
    wire N__8891;
    wire N__8890;
    wire N__8889;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8875;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8856;
    wire N__8851;
    wire N__8848;
    wire N__8845;
    wire N__8842;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8800;
    wire N__8799;
    wire N__8798;
    wire N__8797;
    wire N__8796;
    wire N__8795;
    wire N__8794;
    wire N__8793;
    wire N__8792;
    wire N__8791;
    wire N__8790;
    wire N__8789;
    wire N__8788;
    wire N__8787;
    wire N__8786;
    wire N__8785;
    wire N__8784;
    wire N__8783;
    wire N__8782;
    wire N__8781;
    wire N__8780;
    wire N__8779;
    wire N__8778;
    wire N__8777;
    wire N__8776;
    wire N__8775;
    wire N__8774;
    wire N__8773;
    wire N__8770;
    wire N__8769;
    wire N__8768;
    wire N__8767;
    wire N__8766;
    wire N__8765;
    wire N__8764;
    wire N__8763;
    wire N__8762;
    wire N__8761;
    wire N__8760;
    wire N__8759;
    wire N__8680;
    wire N__8677;
    wire N__8676;
    wire N__8675;
    wire N__8674;
    wire N__8671;
    wire N__8668;
    wire N__8667;
    wire N__8664;
    wire N__8663;
    wire N__8660;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8638;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8608;
    wire N__8605;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8584;
    wire N__8581;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8569;
    wire N__8566;
    wire N__8563;
    wire N__8560;
    wire N__8557;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8536;
    wire N__8533;
    wire N__8530;
    wire N__8527;
    wire N__8524;
    wire N__8523;
    wire N__8520;
    wire N__8517;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8503;
    wire N__8500;
    wire N__8497;
    wire N__8494;
    wire N__8491;
    wire N__8488;
    wire N__8485;
    wire N__8482;
    wire N__8479;
    wire N__8476;
    wire N__8473;
    wire N__8470;
    wire N__8467;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8431;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8354;
    wire N__8353;
    wire N__8352;
    wire N__8347;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8331;
    wire N__8328;
    wire N__8325;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8298;
    wire N__8297;
    wire N__8296;
    wire N__8295;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8259;
    wire N__8254;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8233;
    wire N__8230;
    wire N__8227;
    wire N__8224;
    wire N__8221;
    wire N__8218;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8185;
    wire N__8184;
    wire N__8183;
    wire N__8182;
    wire N__8179;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8163;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8141;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8094;
    wire N__8089;
    wire N__8088;
    wire N__8085;
    wire N__8082;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8070;
    wire N__8069;
    wire N__8066;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8050;
    wire N__8049;
    wire N__8046;
    wire N__8043;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8031;
    wire N__8030;
    wire N__8029;
    wire N__8028;
    wire N__8027;
    wire N__8026;
    wire N__8025;
    wire N__8024;
    wire N__8023;
    wire N__8022;
    wire N__8015;
    wire N__8008;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__8000;
    wire N__7999;
    wire N__7996;
    wire N__7991;
    wire N__7990;
    wire N__7989;
    wire N__7988;
    wire N__7987;
    wire N__7986;
    wire N__7985;
    wire N__7984;
    wire N__7979;
    wire N__7976;
    wire N__7975;
    wire N__7972;
    wire N__7969;
    wire N__7964;
    wire N__7963;
    wire N__7962;
    wire N__7961;
    wire N__7960;
    wire N__7959;
    wire N__7954;
    wire N__7951;
    wire N__7950;
    wire N__7949;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7933;
    wire N__7928;
    wire N__7925;
    wire N__7924;
    wire N__7917;
    wire N__7908;
    wire N__7905;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7885;
    wire N__7880;
    wire N__7877;
    wire N__7872;
    wire N__7865;
    wire N__7862;
    wire N__7857;
    wire N__7854;
    wire N__7847;
    wire N__7844;
    wire N__7839;
    wire N__7836;
    wire N__7833;
    wire N__7828;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7813;
    wire N__7810;
    wire N__7807;
    wire N__7804;
    wire N__7803;
    wire N__7802;
    wire N__7801;
    wire N__7800;
    wire N__7797;
    wire N__7796;
    wire N__7795;
    wire N__7794;
    wire N__7793;
    wire N__7792;
    wire N__7791;
    wire N__7790;
    wire N__7787;
    wire N__7784;
    wire N__7783;
    wire N__7782;
    wire N__7779;
    wire N__7776;
    wire N__7773;
    wire N__7768;
    wire N__7765;
    wire N__7760;
    wire N__7753;
    wire N__7746;
    wire N__7729;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7710;
    wire N__7707;
    wire N__7704;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7681;
    wire N__7678;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7666;
    wire N__7665;
    wire N__7662;
    wire N__7659;
    wire N__7656;
    wire N__7653;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7642;
    wire N__7639;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7621;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7599;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7586;
    wire N__7585;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7567;
    wire N__7564;
    wire N__7561;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7516;
    wire N__7513;
    wire N__7510;
    wire N__7507;
    wire N__7504;
    wire N__7501;
    wire N__7498;
    wire N__7495;
    wire N__7492;
    wire N__7489;
    wire N__7486;
    wire N__7483;
    wire N__7480;
    wire N__7477;
    wire N__7474;
    wire N__7471;
    wire N__7468;
    wire N__7465;
    wire N__7462;
    wire N__7459;
    wire N__7456;
    wire N__7453;
    wire N__7450;
    wire N__7447;
    wire N__7444;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7411;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7401;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7389;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7372;
    wire N__7371;
    wire N__7370;
    wire N__7367;
    wire N__7362;
    wire N__7357;
    wire N__7354;
    wire N__7351;
    wire N__7350;
    wire N__7349;
    wire N__7348;
    wire N__7345;
    wire N__7338;
    wire N__7333;
    wire N__7332;
    wire N__7329;
    wire N__7326;
    wire N__7321;
    wire N__7320;
    wire N__7317;
    wire N__7316;
    wire N__7315;
    wire N__7314;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7302;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7290;
    wire N__7287;
    wire N__7284;
    wire N__7273;
    wire N__7272;
    wire N__7269;
    wire N__7268;
    wire N__7267;
    wire N__7266;
    wire N__7265;
    wire N__7264;
    wire N__7261;
    wire N__7256;
    wire N__7247;
    wire N__7240;
    wire N__7237;
    wire N__7236;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7219;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7188;
    wire N__7185;
    wire N__7180;
    wire N__7179;
    wire N__7178;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7168;
    wire N__7167;
    wire N__7162;
    wire N__7161;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7144;
    wire N__7143;
    wire N__7140;
    wire N__7133;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7084;
    wire N__7081;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7042;
    wire N__7041;
    wire N__7038;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7006;
    wire N__7003;
    wire N__7002;
    wire N__6999;
    wire N__6998;
    wire N__6997;
    wire N__6994;
    wire N__6987;
    wire N__6982;
    wire N__6979;
    wire N__6978;
    wire N__6977;
    wire N__6976;
    wire N__6973;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6957;
    wire N__6954;
    wire N__6949;
    wire N__6948;
    wire N__6947;
    wire N__6946;
    wire N__6941;
    wire N__6936;
    wire N__6931;
    wire N__6928;
    wire N__6927;
    wire N__6924;
    wire N__6921;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6898;
    wire N__6895;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6883;
    wire N__6880;
    wire N__6877;
    wire N__6876;
    wire N__6873;
    wire N__6870;
    wire N__6865;
    wire N__6864;
    wire N__6863;
    wire N__6862;
    wire N__6861;
    wire N__6860;
    wire N__6859;
    wire N__6858;
    wire N__6841;
    wire N__6838;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6823;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6813;
    wire N__6810;
    wire N__6807;
    wire N__6804;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6769;
    wire N__6766;
    wire N__6763;
    wire N__6762;
    wire N__6761;
    wire N__6760;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6752;
    wire N__6751;
    wire N__6748;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6740;
    wire N__6739;
    wire N__6738;
    wire N__6737;
    wire N__6736;
    wire N__6731;
    wire N__6728;
    wire N__6721;
    wire N__6718;
    wire N__6715;
    wire N__6710;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6694;
    wire N__6689;
    wire N__6686;
    wire N__6681;
    wire N__6670;
    wire N__6669;
    wire N__6666;
    wire N__6665;
    wire N__6662;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6654;
    wire N__6653;
    wire N__6652;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6636;
    wire N__6633;
    wire N__6628;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6600;
    wire N__6597;
    wire N__6596;
    wire N__6595;
    wire N__6594;
    wire N__6593;
    wire N__6588;
    wire N__6581;
    wire N__6580;
    wire N__6579;
    wire N__6578;
    wire N__6577;
    wire N__6574;
    wire N__6573;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6552;
    wire N__6549;
    wire N__6538;
    wire N__6537;
    wire N__6536;
    wire N__6535;
    wire N__6534;
    wire N__6531;
    wire N__6530;
    wire N__6529;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6512;
    wire N__6509;
    wire N__6508;
    wire N__6507;
    wire N__6506;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6496;
    wire N__6493;
    wire N__6490;
    wire N__6479;
    wire N__6476;
    wire N__6463;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6441;
    wire N__6438;
    wire N__6435;
    wire N__6432;
    wire N__6431;
    wire N__6426;
    wire N__6423;
    wire N__6418;
    wire N__6417;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6372;
    wire N__6369;
    wire N__6366;
    wire N__6361;
    wire N__6358;
    wire N__6357;
    wire N__6354;
    wire N__6351;
    wire N__6346;
    wire N__6343;
    wire N__6342;
    wire N__6339;
    wire N__6336;
    wire N__6331;
    wire N__6328;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6316;
    wire N__6313;
    wire N__6312;
    wire N__6309;
    wire N__6306;
    wire N__6303;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6288;
    wire N__6287;
    wire N__6286;
    wire N__6283;
    wire N__6276;
    wire N__6275;
    wire N__6274;
    wire N__6269;
    wire N__6264;
    wire N__6259;
    wire N__6256;
    wire N__6255;
    wire N__6254;
    wire N__6253;
    wire N__6252;
    wire N__6249;
    wire N__6242;
    wire N__6241;
    wire N__6240;
    wire N__6237;
    wire N__6232;
    wire N__6227;
    wire N__6220;
    wire N__6219;
    wire N__6218;
    wire N__6213;
    wire N__6210;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6169;
    wire N__6166;
    wire N__6163;
    wire N__6160;
    wire N__6157;
    wire N__6154;
    wire N__6151;
    wire N__6150;
    wire N__6147;
    wire N__6146;
    wire N__6145;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6125;
    wire N__6118;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6108;
    wire N__6107;
    wire N__6106;
    wire N__6105;
    wire N__6104;
    wire N__6103;
    wire N__6098;
    wire N__6097;
    wire N__6094;
    wire N__6093;
    wire N__6090;
    wire N__6089;
    wire N__6088;
    wire N__6087;
    wire N__6086;
    wire N__6083;
    wire N__6082;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6063;
    wire N__6062;
    wire N__6061;
    wire N__6056;
    wire N__6053;
    wire N__6052;
    wire N__6049;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6032;
    wire N__6029;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6009;
    wire N__5998;
    wire N__5983;
    wire N__5982;
    wire N__5979;
    wire N__5978;
    wire N__5977;
    wire N__5976;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5968;
    wire N__5965;
    wire N__5964;
    wire N__5963;
    wire N__5962;
    wire N__5959;
    wire N__5958;
    wire N__5955;
    wire N__5954;
    wire N__5953;
    wire N__5952;
    wire N__5949;
    wire N__5948;
    wire N__5943;
    wire N__5942;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5928;
    wire N__5927;
    wire N__5926;
    wire N__5925;
    wire N__5922;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5895;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5879;
    wire N__5874;
    wire N__5851;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5839;
    wire N__5836;
    wire N__5835;
    wire N__5834;
    wire N__5831;
    wire N__5830;
    wire N__5829;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5817;
    wire N__5814;
    wire N__5809;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5788;
    wire N__5785;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5775;
    wire N__5772;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5730;
    wire N__5727;
    wire N__5724;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5706;
    wire N__5703;
    wire N__5700;
    wire N__5695;
    wire N__5692;
    wire N__5689;
    wire N__5686;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5676;
    wire N__5673;
    wire N__5670;
    wire N__5665;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5650;
    wire N__5647;
    wire N__5646;
    wire N__5645;
    wire N__5644;
    wire N__5641;
    wire N__5638;
    wire N__5633;
    wire N__5630;
    wire N__5625;
    wire N__5620;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5598;
    wire N__5595;
    wire N__5592;
    wire N__5589;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5554;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5541;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5524;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5448;
    wire N__5447;
    wire N__5446;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5432;
    wire N__5431;
    wire N__5430;
    wire N__5427;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5404;
    wire N__5403;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5386;
    wire N__5379;
    wire N__5376;
    wire N__5373;
    wire N__5370;
    wire N__5353;
    wire N__5350;
    wire N__5349;
    wire N__5348;
    wire N__5347;
    wire N__5346;
    wire N__5343;
    wire N__5342;
    wire N__5341;
    wire N__5340;
    wire N__5337;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5295;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5224;
    wire N__5221;
    wire N__5218;
    wire N__5215;
    wire N__5212;
    wire N__5209;
    wire N__5206;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5198;
    wire N__5195;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5181;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5163;
    wire N__5162;
    wire N__5159;
    wire N__5158;
    wire N__5157;
    wire N__5154;
    wire N__5151;
    wire N__5150;
    wire N__5149;
    wire N__5146;
    wire N__5141;
    wire N__5140;
    wire N__5139;
    wire N__5134;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5104;
    wire N__5103;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5089;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5026;
    wire N__5023;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5010;
    wire N__5005;
    wire N__5004;
    wire N__5003;
    wire N__5002;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4981;
    wire N__4980;
    wire N__4975;
    wire N__4974;
    wire N__4973;
    wire N__4972;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4956;
    wire N__4953;
    wire N__4942;
    wire N__4939;
    wire N__4936;
    wire N__4933;
    wire N__4930;
    wire N__4927;
    wire N__4924;
    wire N__4921;
    wire N__4918;
    wire N__4915;
    wire N__4912;
    wire N__4909;
    wire N__4906;
    wire N__4903;
    wire N__4900;
    wire N__4899;
    wire N__4898;
    wire N__4897;
    wire N__4896;
    wire N__4895;
    wire N__4894;
    wire N__4893;
    wire N__4884;
    wire N__4879;
    wire N__4874;
    wire N__4867;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4854;
    wire N__4851;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4824;
    wire N__4823;
    wire N__4822;
    wire N__4821;
    wire N__4820;
    wire N__4819;
    wire N__4816;
    wire N__4815;
    wire N__4814;
    wire N__4813;
    wire N__4812;
    wire N__4811;
    wire N__4810;
    wire N__4809;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4797;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4778;
    wire N__4775;
    wire N__4768;
    wire N__4747;
    wire N__4744;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4704;
    wire N__4703;
    wire N__4702;
    wire N__4701;
    wire N__4698;
    wire N__4695;
    wire N__4692;
    wire N__4687;
    wire N__4678;
    wire N__4675;
    wire N__4672;
    wire N__4669;
    wire N__4666;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4645;
    wire N__4642;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4630;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4596;
    wire N__4593;
    wire N__4590;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4573;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4561;
    wire N__4558;
    wire N__4555;
    wire N__4552;
    wire N__4549;
    wire N__4546;
    wire N__4543;
    wire N__4542;
    wire N__4539;
    wire N__4536;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4486;
    wire N__4483;
    wire N__4482;
    wire N__4479;
    wire N__4476;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4453;
    wire N__4450;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4420;
    wire N__4417;
    wire N__4414;
    wire N__4411;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4384;
    wire N__4381;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4369;
    wire N__4366;
    wire N__4363;
    wire N__4360;
    wire N__4357;
    wire N__4354;
    wire N__4351;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4300;
    wire N__4297;
    wire N__4294;
    wire N__4291;
    wire N__4288;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4273;
    wire N__4270;
    wire N__4267;
    wire N__4264;
    wire N__4261;
    wire N__4258;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4222;
    wire N__4219;
    wire N__4216;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4195;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4183;
    wire N__4180;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4141;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4123;
    wire N__4120;
    wire N__4117;
    wire N__4114;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire U712_CYCLE_TERM_TBIn_0_i;
    wire CLK80_PLL_i_i;
    wire DBRn_c_i_0;
    wire CLK_EN_c;
    wire DBRn_c;
    wire DBR_SYNCZ0Z_0;
    wire A_c_18;
    wire A_c_16;
    wire A_c_6;
    wire A_c_13;
    wire A_c_14;
    wire A_c_7;
    wire \U712_CHIP_RAM.N_543_cascade_ ;
    wire \U712_CHIP_RAM.N_322_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0_0 ;
    wire \U712_CHIP_RAM.CLK_EN_6_0_a3_0_a2_1 ;
    wire \U712_CHIP_RAM.N_599_cascade_ ;
    wire \U712_CHIP_RAM.CLK_EN_6_0 ;
    wire \U712_CHIP_RAM.N_504_cascade_ ;
    wire \U712_CHIP_RAM.N_404 ;
    wire \U712_CHIP_RAM.N_404_cascade_ ;
    wire A_c_5;
    wire A_c_12;
    wire \U712_CHIP_RAM.N_591 ;
    wire VBENn_c;
    wire A_c_8;
    wire A_c_15;
    wire \U712_CHIP_RAM.N_578_cascade_ ;
    wire \U712_CHIP_RAM.N_545 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER18_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_cascade_ ;
    wire \U712_CHIP_RAM.N_552 ;
    wire bfn_8_7_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.N_554_cascade_ ;
    wire BANK0_c;
    wire \U712_CHIP_RAM.N_588 ;
    wire \U712_CHIP_RAM.N_553_cascade_ ;
    wire \U712_CHIP_RAM.N_437_cascade_ ;
    wire \U712_CHIP_RAM.N_414 ;
    wire \U712_CHIP_RAM.N_507 ;
    wire \U712_CHIP_RAM.N_507_cascade_ ;
    wire \U712_CHIP_RAM.N_506 ;
    wire \U712_CHIP_RAM.N_696 ;
    wire \U712_CHIP_RAM.N_534 ;
    wire \U712_CHIP_RAM.N_442_cascade_ ;
    wire \U712_CHIP_RAM.BANK0_RNOZ0Z_3 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.BANK0_RNOZ0Z_1 ;
    wire A_c_20;
    wire \U712_CHIP_RAM.BANK0_RNOZ0Z_2 ;
    wire \U712_CHIP_RAM.N_605_cascade_ ;
    wire \U712_CHIP_RAM.N_605 ;
    wire \U712_CHIP_RAM.N_697_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2_cascade_ ;
    wire \U712_CHIP_RAM.N_539 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_697 ;
    wire \U712_CHIP_RAM.N_551 ;
    wire \U712_CHIP_RAM.N_580 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire \U712_CHIP_RAM.N_505 ;
    wire \U712_CHIP_RAM.N_437 ;
    wire \U712_CHIP_RAM.N_587 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.N_70 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire REGSPACEn_c;
    wire \U712_REG_SM.N_513_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1 ;
    wire \U712_CHIP_RAM.N_589 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ;
    wire \U712_REG_SM.N_694_cascade_ ;
    wire \U712_REG_SM.N_522_cascade_ ;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ;
    wire \U712_REG_SM.N_429_cascade_ ;
    wire \U712_REG_SM.N_511_cascade_ ;
    wire \U712_REG_SM.N_694 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ;
    wire \U712_CHIP_RAM.N_700 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0_a2_0_1 ;
    wire \U712_CHIP_RAM.N_578 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.N_405 ;
    wire \U712_CHIP_RAM.N_699 ;
    wire \U712_CHIP_RAM.N_597_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_ ;
    wire LATCH_CLK_c;
    wire \U712_CHIP_RAM.N_528 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_REG_SM.N_482_cascade_ ;
    wire RAMENn_c;
    wire \U712_CHIP_RAM.N_527 ;
    wire TSn_c;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_553 ;
    wire \U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.N_597 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_ ;
    wire \U712_CHIP_RAM.N_537 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_703 ;
    wire \U712_CHIP_RAM.N_530_cascade_ ;
    wire \U712_CHIP_RAM.N_600 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0 ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.BANK0_0_sqmuxa_1 ;
    wire DBDIR_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ;
    wire \U712_CHIP_RAM.DBENn_8_0 ;
    wire \U712_REG_SM.START_RSTZ0 ;
    wire \U712_REG_SM.STATE_COUNT_srsts_i_i_i_a2_0_0_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_2 ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_0 ;
    wire \U712_REG_SM.START_RST_0_sqmuxa ;
    wire \U712_REG_SM.un1_STATE_COUNT_4_i_i_0_0 ;
    wire \U712_REG_SM.DS_EN_RNOZ0Z_0 ;
    wire \U712_REG_SM.N_515 ;
    wire \U712_REG_SM.N_443 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire ASn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire RESETn_c_i;
    wire N_549;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_11_5_0_;
    wire \U712_CHIP_RAM.REFRESH5lto1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH5lto2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire C1_c_g;
    wire A_c_2;
    wire A_c_9;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.REFRESH_RST_cascade_ ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_595 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0 ;
    wire \U712_CYCLE_TERM.TACK_EN_RNOZ0Z_0_cascade_ ;
    wire \U712_CYCLE_TERM.N_598_cascade_ ;
    wire \U712_REG_SM.N_422 ;
    wire \U712_REG_SM.N_514 ;
    wire REG_TACK;
    wire CPU_TACKm;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.N_571_cascade_ ;
    wire \U712_REG_SM.N_480 ;
    wire \U712_REG_SM.REG_TACK_RNOZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_REG_SM.N_407 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire RnW_c;
    wire WRITE_CYCLEm;
    wire N_483;
    wire CMA_c_10;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.un1_CMA28_0_i ;
    wire \U712_CHIP_RAM.N_412_cascade_ ;
    wire A_c_3;
    wire \U712_CHIP_RAM.N_478 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_ ;
    wire CMA_c_0;
    wire CMA_c_2;
    wire A_c_4;
    wire A_c_11;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CLK40_PLL_i;
    wire CLK40_PLL_i_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.N_598 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ1Z_2 ;
    wire \U712_CYCLE_TERM.N_440 ;
    wire \U712_CYCLE_TERM.un13_0 ;
    wire RESETn_c;
    wire \U712_CYCLE_TERM.N_566 ;
    wire \U712_CYCLE_TERM.un13_0_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.N_93 ;
    wire A_c_10;
    wire \U712_CHIP_RAM.N_455 ;
    wire TACK_OUTn;
    wire \U712_CYCLE_TERM.RAM_CYCLEZ0 ;
    wire TACK_EN;
    wire U712_CYCLE_TERM_TCIn_0_i;
    wire CONSTANT_ONE_NET;
    wire \U712_BYTE_ENABLE.N_563_cascade_ ;
    wire N_56_i;
    wire WEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire A_c_17;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CMA_5_i_0_8 ;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire N_58_i;
    wire \U712_BYTE_ENABLE.N_410 ;
    wire \U712_BYTE_ENABLE.N_559 ;
    wire N_129_i;
    wire CASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire RASn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ;
    wire \U712_CHIP_RAM.N_412 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_ ;
    wire CMA_c_4;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ;
    wire un1_UDSn_i_0_0;
    wire DS_ENm;
    wire un1_LDSn_i_0_0;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire DRA_c_1;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire N_57_i;
    wire DBENn_c;
    wire DMA_CYCLEm;
    wire N_59_i;
    wire \U712_BYTE_ENABLE.N_557 ;
    wire CPU_CYCLEm;
    wire \U712_BYTE_ENABLE.N_561 ;
    wire \U712_BYTE_ENABLE.N_397_i ;
    wire N_130_i;
    wire N_127_i;
    wire A_c_0;
    wire A_c_1;
    wire SIZ_c_0;
    wire SIZ_c_1;
    wire N_128_i;
    wire DRA_c_6;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire AGNUS_REV_c;
    wire RAS0n_c;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire REG_CYCLEm;
    wire CASLn_c;
    wire CASUn_c;
    wire DRDENn_c;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__4102),
            .RESETB(N__7546),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__12194),
            .DIN(N__12193),
            .DOUT(N__12192),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__12194),
            .PADOUT(N__12193),
            .PADIN(N__12192),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9849),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__12185),
            .DIN(N__12184),
            .DOUT(N__12183),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__12185),
            .PADOUT(N__12184),
            .PADIN(N__12183),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__12176),
            .DIN(N__12175),
            .DOUT(N__12174),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__12176),
            .PADOUT(N__12175),
            .PADIN(N__12174),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9187),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__12167),
            .DIN(N__12166),
            .DOUT(N__12165),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__12167),
            .PADOUT(N__12166),
            .PADIN(N__12165),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7099),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__12158),
            .DIN(N__12157),
            .DOUT(N__12156),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__12158),
            .PADOUT(N__12157),
            .PADIN(N__12156),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__12149),
            .DIN(N__12148),
            .DOUT(N__12147),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__12149),
            .PADOUT(N__12148),
            .PADIN(N__12147),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__12140),
            .DIN(N__12139),
            .DOUT(N__12138),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__12140),
            .PADOUT(N__12139),
            .PADIN(N__12138),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__12131),
            .DIN(N__12130),
            .DOUT(N__12129),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__12131),
            .PADOUT(N__12130),
            .PADIN(N__12129),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__12122),
            .DIN(N__12121),
            .DOUT(N__12120),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__12122),
            .PADOUT(N__12121),
            .PADIN(N__12120),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__12113),
            .DIN(N__12112),
            .DOUT(N__12111),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__12113),
            .PADOUT(N__12112),
            .PADIN(N__12111),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__12104),
            .DIN(N__12103),
            .DOUT(N__12102),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__12104),
            .PADOUT(N__12103),
            .PADIN(N__12102),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8542),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__12095),
            .DIN(N__12094),
            .DOUT(N__12093),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__12095),
            .PADOUT(N__12094),
            .PADIN(N__12093),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9202),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__12086),
            .DIN(N__12085),
            .DOUT(N__12084),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__12086),
            .PADOUT(N__12085),
            .PADIN(N__12084),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__12077),
            .DIN(N__12076),
            .DOUT(N__12075),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__12077),
            .PADOUT(N__12076),
            .PADIN(N__12075),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5607),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__12068),
            .DIN(N__12067),
            .DOUT(N__12066),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__12068),
            .PADOUT(N__12067),
            .PADIN(N__12066),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__12059),
            .DIN(N__12058),
            .DOUT(N__12057),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__12059),
            .PADOUT(N__12058),
            .PADIN(N__12057),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__12050),
            .DIN(N__12049),
            .DOUT(N__12048),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__12050),
            .PADOUT(N__12049),
            .PADIN(N__12048),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4348),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__12041),
            .DIN(N__12040),
            .DOUT(N__12039),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__12041),
            .PADOUT(N__12040),
            .PADIN(N__12039),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__12032),
            .DIN(N__12031),
            .DOUT(N__12030),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__12032),
            .PADOUT(N__12031),
            .PADIN(N__12030),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__12023),
            .DIN(N__12022),
            .DOUT(N__12021),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__12023),
            .PADOUT(N__12022),
            .PADIN(N__12021),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7465),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__12014),
            .DIN(N__12013),
            .DOUT(N__12012),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__12014),
            .PADOUT(N__12013),
            .PADIN(N__12012),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__12005),
            .DIN(N__12004),
            .DOUT(N__12003),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__12005),
            .PADOUT(N__12004),
            .PADIN(N__12003),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8320),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11996),
            .DIN(N__11995),
            .DOUT(N__11994),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11996),
            .PADOUT(N__11995),
            .PADIN(N__11994),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__11987),
            .DIN(N__11986),
            .DOUT(N__11985),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__11987),
            .PADOUT(N__11986),
            .PADIN(N__11985),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10798),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__11978),
            .DIN(N__11977),
            .DOUT(N__11976),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__11978),
            .PADOUT(N__11977),
            .PADIN(N__11976),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11969),
            .DIN(N__11968),
            .DOUT(N__11967),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11969),
            .PADOUT(N__11968),
            .PADIN(N__11967),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__11960),
            .DIN(N__11959),
            .DOUT(N__11958),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__11960),
            .PADOUT(N__11959),
            .PADIN(N__11958),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMENn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11951),
            .DIN(N__11950),
            .DOUT(N__11949),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11951),
            .PADOUT(N__11950),
            .PADIN(N__11949),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__11942),
            .DIN(N__11941),
            .DOUT(N__11940),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__11942),
            .PADOUT(N__11941),
            .PADIN(N__11940),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__11933),
            .DIN(N__11932),
            .DOUT(N__11931),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__11933),
            .PADOUT(N__11932),
            .PADIN(N__11931),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6391),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__11924),
            .DIN(N__11923),
            .DOUT(N__11922),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__11924),
            .PADOUT(N__11923),
            .PADIN(N__11922),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11915),
            .DIN(N__11914),
            .DOUT(N__11913),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11915),
            .PADOUT(N__11914),
            .PADIN(N__11913),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11906),
            .DIN(N__11905),
            .DOUT(N__11904),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11906),
            .PADOUT(N__11905),
            .PADIN(N__11904),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11897),
            .DIN(N__11896),
            .DOUT(N__11895),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11897),
            .PADOUT(N__11896),
            .PADIN(N__11895),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuf_iopad (
            .OE(N__11888),
            .DIN(N__11887),
            .DOUT(N__11886),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TCIn_obuf_preio (
            .PADOEN(N__11888),
            .PADOUT(N__11887),
            .PADIN(N__11886),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7567),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__11879),
            .DIN(N__11878),
            .DOUT(N__11877),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__11879),
            .PADOUT(N__11878),
            .PADIN(N__11877),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__11870),
            .DIN(N__11869),
            .DOUT(N__11868),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__11870),
            .PADOUT(N__11869),
            .PADIN(N__11868),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9118),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__11861),
            .DIN(N__11860),
            .DOUT(N__11859),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__11861),
            .PADOUT(N__11860),
            .PADIN(N__11859),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4612),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__11852),
            .DIN(N__11851),
            .DOUT(N__11850),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__11852),
            .PADOUT(N__11851),
            .PADIN(N__11850),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__11843),
            .DIN(N__11842),
            .DOUT(N__11841),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__11843),
            .PADOUT(N__11842),
            .PADIN(N__11841),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6463),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_0_iopad (
            .OE(N__11834),
            .DIN(N__11833),
            .DOUT(N__11832),
            .PACKAGEPIN(DA[0]));
    defparam DA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_0_preio (
            .PADOEN(N__11834),
            .PADOUT(N__11833),
            .PADIN(N__11832),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6814),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11825),
            .DIN(N__11824),
            .DOUT(N__11823),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11825),
            .PADOUT(N__11824),
            .PADIN(N__11823),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8464),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11816),
            .DIN(N__11815),
            .DOUT(N__11814),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11816),
            .PADOUT(N__11815),
            .PADIN(N__11814),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11807),
            .DIN(N__11806),
            .DOUT(N__11805),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11807),
            .PADOUT(N__11806),
            .PADIN(N__11805),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11798),
            .DIN(N__11797),
            .DOUT(N__11796),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11798),
            .PADOUT(N__11797),
            .PADIN(N__11796),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__11789),
            .DIN(N__11788),
            .DOUT(N__11787),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__11789),
            .PADOUT(N__11788),
            .PADIN(N__11787),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__11780),
            .DIN(N__11779),
            .DOUT(N__11778),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__11780),
            .PADOUT(N__11779),
            .PADIN(N__11778),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7075),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11771),
            .DIN(N__11770),
            .DOUT(N__11769),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11771),
            .PADOUT(N__11770),
            .PADIN(N__11769),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11762),
            .DIN(N__11761),
            .DOUT(N__11760),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11762),
            .PADOUT(N__11761),
            .PADIN(N__11760),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8141),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__11753),
            .DIN(N__11752),
            .DOUT(N__11751),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__11753),
            .PADOUT(N__11752),
            .PADIN(N__11751),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8824),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11744),
            .DIN(N__11743),
            .DOUT(N__11742),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11744),
            .PADOUT(N__11743),
            .PADIN(N__11742),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11179),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11735),
            .DIN(N__11734),
            .DOUT(N__11733),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11735),
            .PADOUT(N__11734),
            .PADIN(N__11733),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8404),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11726),
            .DIN(N__11725),
            .DOUT(N__11724),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11726),
            .PADOUT(N__11725),
            .PADIN(N__11724),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8491),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__11717),
            .DIN(N__11716),
            .DOUT(N__11715),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__11717),
            .PADOUT(N__11716),
            .PADIN(N__11715),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6462),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11708),
            .DIN(N__11707),
            .DOUT(N__11706),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11708),
            .PADOUT(N__11707),
            .PADIN(N__11706),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__11699),
            .DIN(N__11698),
            .DOUT(N__11697),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__11699),
            .PADOUT(N__11698),
            .PADIN(N__11697),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__11690),
            .DIN(N__11689),
            .DOUT(N__11688),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__11690),
            .PADOUT(N__11689),
            .PADIN(N__11688),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9868),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__11681),
            .DIN(N__11680),
            .DOUT(N__11679),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__11681),
            .PADOUT(N__11680),
            .PADIN(N__11679),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8383),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__11672),
            .DIN(N__11671),
            .DOUT(N__11670),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__11672),
            .PADOUT(N__11671),
            .PADIN(N__11670),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5743),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__11663),
            .DIN(N__11662),
            .DOUT(N__11661),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__11663),
            .PADOUT(N__11662),
            .PADIN(N__11661),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9256),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__11654),
            .DIN(N__11653),
            .DOUT(N__11652),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__11654),
            .PADOUT(N__11653),
            .PADIN(N__11652),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11645),
            .DIN(N__11644),
            .DOUT(N__11643),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11645),
            .PADOUT(N__11644),
            .PADIN(N__11643),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_2_iopad (
            .OE(N__11636),
            .DIN(N__11635),
            .DOUT(N__11634),
            .PACKAGEPIN(DA[2]));
    defparam DA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_2_preio (
            .PADOEN(N__11636),
            .PADOUT(N__11635),
            .PADIN(N__11634),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7414),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11627),
            .DIN(N__11626),
            .DOUT(N__11625),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11627),
            .PADOUT(N__11626),
            .PADIN(N__11625),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11618),
            .DIN(N__11617),
            .DOUT(N__11616),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11618),
            .PADOUT(N__11617),
            .PADIN(N__11616),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__11609),
            .DIN(N__11608),
            .DOUT(N__11607),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__11609),
            .PADOUT(N__11608),
            .PADIN(N__11607),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7063),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__11600),
            .DIN(N__11599),
            .DOUT(N__11598),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__11600),
            .PADOUT(N__11599),
            .PADIN(N__11598),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11122),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__11591),
            .DIN(N__11590),
            .DOUT(N__11589),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__11591),
            .PADOUT(N__11590),
            .PADIN(N__11589),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__11582),
            .DIN(N__11581),
            .DOUT(N__11580),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__11582),
            .PADOUT(N__11581),
            .PADIN(N__11580),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9694),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__11573),
            .DIN(N__11572),
            .DOUT(N__11571),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__11573),
            .PADOUT(N__11572),
            .PADIN(N__11571),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7609),
            .DIN0(),
            .DOUT0(N__7666),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__11564),
            .DIN(N__11563),
            .DOUT(N__11562),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__11564),
            .PADOUT(N__11563),
            .PADIN(N__11562),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7453),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__11555),
            .DIN(N__11554),
            .DOUT(N__11553),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__11555),
            .PADOUT(N__11554),
            .PADIN(N__11553),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11546),
            .DIN(N__11545),
            .DOUT(N__11544),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11546),
            .PADOUT(N__11545),
            .PADIN(N__11544),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__11537),
            .DIN(N__11536),
            .DOUT(N__11535),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__11537),
            .PADOUT(N__11536),
            .PADIN(N__11535),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8569),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuf_iopad (
            .OE(N__11528),
            .DIN(N__11527),
            .DOUT(N__11526),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TBIn_obuf_preio (
            .PADOEN(N__11528),
            .PADOUT(N__11527),
            .PADIN(N__11526),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4273),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__11519),
            .DIN(N__11518),
            .DOUT(N__11517),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__11519),
            .PADOUT(N__11518),
            .PADIN(N__11517),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__11510),
            .DIN(N__11509),
            .DOUT(N__11508),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__11510),
            .PADOUT(N__11509),
            .PADIN(N__11508),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_1_iopad (
            .OE(N__11501),
            .DIN(N__11500),
            .DOUT(N__11499),
            .PACKAGEPIN(DA[1]));
    defparam DA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_1_preio (
            .PADOEN(N__11501),
            .PADOUT(N__11500),
            .PADIN(N__11499),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7717),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11492),
            .DIN(N__11491),
            .DOUT(N__11490),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11492),
            .PADOUT(N__11491),
            .PADIN(N__11490),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11483),
            .DIN(N__11482),
            .DOUT(N__11481),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11483),
            .PADOUT(N__11482),
            .PADIN(N__11481),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__11474),
            .DIN(N__11473),
            .DOUT(N__11472),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__11474),
            .PADOUT(N__11473),
            .PADIN(N__11472),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8215),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__11465),
            .DIN(N__11464),
            .DOUT(N__11463),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__11465),
            .PADOUT(N__11464),
            .PADIN(N__11463),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9358),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__11456),
            .DIN(N__11455),
            .DOUT(N__11454),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__11456),
            .PADOUT(N__11455),
            .PADIN(N__11454),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11107),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__11447),
            .DIN(N__11446),
            .DOUT(N__11445),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__11447),
            .PADOUT(N__11446),
            .PADIN(N__11445),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4216),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__11438),
            .DIN(N__11437),
            .DOUT(N__11436),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__11438),
            .PADOUT(N__11437),
            .PADIN(N__11436),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11429),
            .DIN(N__11428),
            .DOUT(N__11427),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11429),
            .PADOUT(N__11428),
            .PADIN(N__11427),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__11420),
            .DIN(N__11419),
            .DOUT(N__11418),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__11420),
            .PADOUT(N__11419),
            .PADIN(N__11418),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8611),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__11411),
            .DIN(N__11410),
            .DOUT(N__11409),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__11411),
            .PADOUT(N__11410),
            .PADIN(N__11409),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__11402),
            .DIN(N__11401),
            .DOUT(N__11400),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__11402),
            .PADOUT(N__11401),
            .PADIN(N__11400),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__11393),
            .DIN(N__11392),
            .DOUT(N__11391),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__11393),
            .PADOUT(N__11392),
            .PADIN(N__11391),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5692),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__11384),
            .DIN(N__11383),
            .DOUT(N__11382),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__11384),
            .PADOUT(N__11383),
            .PADIN(N__11382),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9313),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11375),
            .DIN(N__11374),
            .DOUT(N__11373),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11375),
            .PADOUT(N__11374),
            .PADIN(N__11373),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8149),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11366),
            .DIN(N__11365),
            .DOUT(N__11364),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11366),
            .PADOUT(N__11365),
            .PADIN(N__11364),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11357),
            .DIN(N__11356),
            .DOUT(N__11355),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11357),
            .PADOUT(N__11356),
            .PADIN(N__11355),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8148),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11348),
            .DIN(N__11347),
            .DOUT(N__11346),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11348),
            .PADOUT(N__11347),
            .PADIN(N__11346),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4252),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2768 (
            .O(N__11329),
            .I(N__11326));
    LocalMux I__2767 (
            .O(N__11326),
            .I(N__11321));
    InMux I__2766 (
            .O(N__11325),
            .I(N__11317));
    InMux I__2765 (
            .O(N__11324),
            .I(N__11313));
    Span4Mux_v I__2764 (
            .O(N__11321),
            .I(N__11310));
    InMux I__2763 (
            .O(N__11320),
            .I(N__11307));
    LocalMux I__2762 (
            .O(N__11317),
            .I(N__11304));
    InMux I__2761 (
            .O(N__11316),
            .I(N__11301));
    LocalMux I__2760 (
            .O(N__11313),
            .I(N__11297));
    Span4Mux_v I__2759 (
            .O(N__11310),
            .I(N__11294));
    LocalMux I__2758 (
            .O(N__11307),
            .I(N__11289));
    Sp12to4 I__2757 (
            .O(N__11304),
            .I(N__11289));
    LocalMux I__2756 (
            .O(N__11301),
            .I(N__11286));
    InMux I__2755 (
            .O(N__11300),
            .I(N__11283));
    Span12Mux_h I__2754 (
            .O(N__11297),
            .I(N__11280));
    Sp12to4 I__2753 (
            .O(N__11294),
            .I(N__11275));
    Span12Mux_v I__2752 (
            .O(N__11289),
            .I(N__11275));
    Span12Mux_h I__2751 (
            .O(N__11286),
            .I(N__11270));
    LocalMux I__2750 (
            .O(N__11283),
            .I(N__11270));
    Span12Mux_v I__2749 (
            .O(N__11280),
            .I(N__11267));
    Span12Mux_h I__2748 (
            .O(N__11275),
            .I(N__11262));
    Span12Mux_v I__2747 (
            .O(N__11270),
            .I(N__11262));
    Odrv12 I__2746 (
            .O(N__11267),
            .I(CASLn_c));
    Odrv12 I__2745 (
            .O(N__11262),
            .I(CASLn_c));
    InMux I__2744 (
            .O(N__11257),
            .I(N__11252));
    InMux I__2743 (
            .O(N__11256),
            .I(N__11249));
    InMux I__2742 (
            .O(N__11255),
            .I(N__11246));
    LocalMux I__2741 (
            .O(N__11252),
            .I(N__11242));
    LocalMux I__2740 (
            .O(N__11249),
            .I(N__11237));
    LocalMux I__2739 (
            .O(N__11246),
            .I(N__11237));
    InMux I__2738 (
            .O(N__11245),
            .I(N__11234));
    Span4Mux_v I__2737 (
            .O(N__11242),
            .I(N__11231));
    Span4Mux_h I__2736 (
            .O(N__11237),
            .I(N__11228));
    LocalMux I__2735 (
            .O(N__11234),
            .I(N__11225));
    Span4Mux_v I__2734 (
            .O(N__11231),
            .I(N__11219));
    Span4Mux_h I__2733 (
            .O(N__11228),
            .I(N__11219));
    Span4Mux_v I__2732 (
            .O(N__11225),
            .I(N__11215));
    InMux I__2731 (
            .O(N__11224),
            .I(N__11212));
    Span4Mux_h I__2730 (
            .O(N__11219),
            .I(N__11209));
    InMux I__2729 (
            .O(N__11218),
            .I(N__11206));
    Sp12to4 I__2728 (
            .O(N__11215),
            .I(N__11201));
    LocalMux I__2727 (
            .O(N__11212),
            .I(N__11201));
    Span4Mux_h I__2726 (
            .O(N__11209),
            .I(N__11196));
    LocalMux I__2725 (
            .O(N__11206),
            .I(N__11196));
    Span12Mux_h I__2724 (
            .O(N__11201),
            .I(N__11193));
    Span4Mux_h I__2723 (
            .O(N__11196),
            .I(N__11190));
    Span12Mux_v I__2722 (
            .O(N__11193),
            .I(N__11187));
    Span4Mux_v I__2721 (
            .O(N__11190),
            .I(N__11184));
    Odrv12 I__2720 (
            .O(N__11187),
            .I(CASUn_c));
    Odrv4 I__2719 (
            .O(N__11184),
            .I(CASUn_c));
    IoInMux I__2718 (
            .O(N__11179),
            .I(N__11176));
    LocalMux I__2717 (
            .O(N__11176),
            .I(N__11173));
    Span12Mux_s7_v I__2716 (
            .O(N__11173),
            .I(N__11170));
    Odrv12 I__2715 (
            .O(N__11170),
            .I(DRDENn_c));
    InMux I__2714 (
            .O(N__11167),
            .I(N__11164));
    LocalMux I__2713 (
            .O(N__11164),
            .I(N__11161));
    Odrv4 I__2712 (
            .O(N__11161),
            .I(\U712_BYTE_ENABLE.N_561 ));
    InMux I__2711 (
            .O(N__11158),
            .I(N__11152));
    InMux I__2710 (
            .O(N__11157),
            .I(N__11149));
    CascadeMux I__2709 (
            .O(N__11156),
            .I(N__11146));
    CascadeMux I__2708 (
            .O(N__11155),
            .I(N__11143));
    LocalMux I__2707 (
            .O(N__11152),
            .I(N__11138));
    LocalMux I__2706 (
            .O(N__11149),
            .I(N__11138));
    InMux I__2705 (
            .O(N__11146),
            .I(N__11133));
    InMux I__2704 (
            .O(N__11143),
            .I(N__11133));
    Span4Mux_v I__2703 (
            .O(N__11138),
            .I(N__11130));
    LocalMux I__2702 (
            .O(N__11133),
            .I(N__11127));
    Odrv4 I__2701 (
            .O(N__11130),
            .I(\U712_BYTE_ENABLE.N_397_i ));
    Odrv4 I__2700 (
            .O(N__11127),
            .I(\U712_BYTE_ENABLE.N_397_i ));
    IoInMux I__2699 (
            .O(N__11122),
            .I(N__11119));
    LocalMux I__2698 (
            .O(N__11119),
            .I(N__11116));
    Span4Mux_s0_v I__2697 (
            .O(N__11116),
            .I(N__11113));
    Span4Mux_v I__2696 (
            .O(N__11113),
            .I(N__11110));
    Odrv4 I__2695 (
            .O(N__11110),
            .I(N_130_i));
    IoInMux I__2694 (
            .O(N__11107),
            .I(N__11104));
    LocalMux I__2693 (
            .O(N__11104),
            .I(N__11101));
    IoSpan4Mux I__2692 (
            .O(N__11101),
            .I(N__11098));
    Span4Mux_s2_v I__2691 (
            .O(N__11098),
            .I(N__11095));
    Span4Mux_v I__2690 (
            .O(N__11095),
            .I(N__11092));
    Odrv4 I__2689 (
            .O(N__11092),
            .I(N_127_i));
    InMux I__2688 (
            .O(N__11089),
            .I(N__11076));
    InMux I__2687 (
            .O(N__11088),
            .I(N__11076));
    InMux I__2686 (
            .O(N__11087),
            .I(N__11076));
    InMux I__2685 (
            .O(N__11086),
            .I(N__11071));
    InMux I__2684 (
            .O(N__11085),
            .I(N__11071));
    InMux I__2683 (
            .O(N__11084),
            .I(N__11066));
    InMux I__2682 (
            .O(N__11083),
            .I(N__11066));
    LocalMux I__2681 (
            .O(N__11076),
            .I(N__11060));
    LocalMux I__2680 (
            .O(N__11071),
            .I(N__11060));
    LocalMux I__2679 (
            .O(N__11066),
            .I(N__11057));
    InMux I__2678 (
            .O(N__11065),
            .I(N__11054));
    Span4Mux_v I__2677 (
            .O(N__11060),
            .I(N__11048));
    Span4Mux_v I__2676 (
            .O(N__11057),
            .I(N__11048));
    LocalMux I__2675 (
            .O(N__11054),
            .I(N__11045));
    InMux I__2674 (
            .O(N__11053),
            .I(N__11042));
    Span4Mux_h I__2673 (
            .O(N__11048),
            .I(N__11039));
    Span4Mux_v I__2672 (
            .O(N__11045),
            .I(N__11036));
    LocalMux I__2671 (
            .O(N__11042),
            .I(N__11033));
    Sp12to4 I__2670 (
            .O(N__11039),
            .I(N__11026));
    Sp12to4 I__2669 (
            .O(N__11036),
            .I(N__11026));
    Span12Mux_v I__2668 (
            .O(N__11033),
            .I(N__11026));
    Span12Mux_h I__2667 (
            .O(N__11026),
            .I(N__11023));
    Odrv12 I__2666 (
            .O(N__11023),
            .I(A_c_0));
    InMux I__2665 (
            .O(N__11020),
            .I(N__11013));
    InMux I__2664 (
            .O(N__11019),
            .I(N__11013));
    InMux I__2663 (
            .O(N__11018),
            .I(N__11007));
    LocalMux I__2662 (
            .O(N__11013),
            .I(N__11002));
    InMux I__2661 (
            .O(N__11012),
            .I(N__10995));
    InMux I__2660 (
            .O(N__11011),
            .I(N__10995));
    InMux I__2659 (
            .O(N__11010),
            .I(N__10995));
    LocalMux I__2658 (
            .O(N__11007),
            .I(N__10992));
    InMux I__2657 (
            .O(N__11006),
            .I(N__10989));
    InMux I__2656 (
            .O(N__11005),
            .I(N__10986));
    Span4Mux_v I__2655 (
            .O(N__11002),
            .I(N__10983));
    LocalMux I__2654 (
            .O(N__10995),
            .I(N__10980));
    Span4Mux_v I__2653 (
            .O(N__10992),
            .I(N__10977));
    LocalMux I__2652 (
            .O(N__10989),
            .I(N__10974));
    LocalMux I__2651 (
            .O(N__10986),
            .I(N__10971));
    Span4Mux_v I__2650 (
            .O(N__10983),
            .I(N__10966));
    Span4Mux_v I__2649 (
            .O(N__10980),
            .I(N__10966));
    Span4Mux_v I__2648 (
            .O(N__10977),
            .I(N__10961));
    Span4Mux_v I__2647 (
            .O(N__10974),
            .I(N__10961));
    Span12Mux_v I__2646 (
            .O(N__10971),
            .I(N__10958));
    Sp12to4 I__2645 (
            .O(N__10966),
            .I(N__10953));
    Sp12to4 I__2644 (
            .O(N__10961),
            .I(N__10953));
    Span12Mux_h I__2643 (
            .O(N__10958),
            .I(N__10950));
    Span12Mux_h I__2642 (
            .O(N__10953),
            .I(N__10947));
    Odrv12 I__2641 (
            .O(N__10950),
            .I(A_c_1));
    Odrv12 I__2640 (
            .O(N__10947),
            .I(A_c_1));
    InMux I__2639 (
            .O(N__10942),
            .I(N__10937));
    CascadeMux I__2638 (
            .O(N__10941),
            .I(N__10933));
    CascadeMux I__2637 (
            .O(N__10940),
            .I(N__10930));
    LocalMux I__2636 (
            .O(N__10937),
            .I(N__10924));
    InMux I__2635 (
            .O(N__10936),
            .I(N__10917));
    InMux I__2634 (
            .O(N__10933),
            .I(N__10917));
    InMux I__2633 (
            .O(N__10930),
            .I(N__10917));
    CascadeMux I__2632 (
            .O(N__10929),
            .I(N__10914));
    CascadeMux I__2631 (
            .O(N__10928),
            .I(N__10911));
    CascadeMux I__2630 (
            .O(N__10927),
            .I(N__10908));
    Span4Mux_h I__2629 (
            .O(N__10924),
            .I(N__10905));
    LocalMux I__2628 (
            .O(N__10917),
            .I(N__10902));
    InMux I__2627 (
            .O(N__10914),
            .I(N__10897));
    InMux I__2626 (
            .O(N__10911),
            .I(N__10897));
    InMux I__2625 (
            .O(N__10908),
            .I(N__10894));
    Span4Mux_v I__2624 (
            .O(N__10905),
            .I(N__10885));
    Span4Mux_h I__2623 (
            .O(N__10902),
            .I(N__10885));
    LocalMux I__2622 (
            .O(N__10897),
            .I(N__10885));
    LocalMux I__2621 (
            .O(N__10894),
            .I(N__10885));
    Span4Mux_h I__2620 (
            .O(N__10885),
            .I(N__10882));
    Span4Mux_v I__2619 (
            .O(N__10882),
            .I(N__10879));
    Sp12to4 I__2618 (
            .O(N__10879),
            .I(N__10876));
    Span12Mux_h I__2617 (
            .O(N__10876),
            .I(N__10873));
    Odrv12 I__2616 (
            .O(N__10873),
            .I(SIZ_c_0));
    InMux I__2615 (
            .O(N__10870),
            .I(N__10865));
    InMux I__2614 (
            .O(N__10869),
            .I(N__10862));
    CascadeMux I__2613 (
            .O(N__10868),
            .I(N__10859));
    LocalMux I__2612 (
            .O(N__10865),
            .I(N__10854));
    LocalMux I__2611 (
            .O(N__10862),
            .I(N__10851));
    InMux I__2610 (
            .O(N__10859),
            .I(N__10844));
    InMux I__2609 (
            .O(N__10858),
            .I(N__10844));
    InMux I__2608 (
            .O(N__10857),
            .I(N__10844));
    Span4Mux_h I__2607 (
            .O(N__10854),
            .I(N__10836));
    Span4Mux_v I__2606 (
            .O(N__10851),
            .I(N__10836));
    LocalMux I__2605 (
            .O(N__10844),
            .I(N__10833));
    InMux I__2604 (
            .O(N__10843),
            .I(N__10828));
    InMux I__2603 (
            .O(N__10842),
            .I(N__10828));
    InMux I__2602 (
            .O(N__10841),
            .I(N__10825));
    Span4Mux_v I__2601 (
            .O(N__10836),
            .I(N__10822));
    Span4Mux_h I__2600 (
            .O(N__10833),
            .I(N__10815));
    LocalMux I__2599 (
            .O(N__10828),
            .I(N__10815));
    LocalMux I__2598 (
            .O(N__10825),
            .I(N__10815));
    Span4Mux_v I__2597 (
            .O(N__10822),
            .I(N__10812));
    Sp12to4 I__2596 (
            .O(N__10815),
            .I(N__10809));
    Sp12to4 I__2595 (
            .O(N__10812),
            .I(N__10804));
    Span12Mux_v I__2594 (
            .O(N__10809),
            .I(N__10804));
    Span12Mux_h I__2593 (
            .O(N__10804),
            .I(N__10801));
    Odrv12 I__2592 (
            .O(N__10801),
            .I(SIZ_c_1));
    IoInMux I__2591 (
            .O(N__10798),
            .I(N__10795));
    LocalMux I__2590 (
            .O(N__10795),
            .I(N__10792));
    Span4Mux_s3_v I__2589 (
            .O(N__10792),
            .I(N__10789));
    Odrv4 I__2588 (
            .O(N__10789),
            .I(N_128_i));
    InMux I__2587 (
            .O(N__10786),
            .I(N__10782));
    InMux I__2586 (
            .O(N__10785),
            .I(N__10779));
    LocalMux I__2585 (
            .O(N__10782),
            .I(N__10773));
    LocalMux I__2584 (
            .O(N__10779),
            .I(N__10773));
    InMux I__2583 (
            .O(N__10778),
            .I(N__10770));
    Span4Mux_h I__2582 (
            .O(N__10773),
            .I(N__10764));
    LocalMux I__2581 (
            .O(N__10770),
            .I(N__10764));
    InMux I__2580 (
            .O(N__10769),
            .I(N__10761));
    Span4Mux_v I__2579 (
            .O(N__10764),
            .I(N__10758));
    LocalMux I__2578 (
            .O(N__10761),
            .I(N__10755));
    Span4Mux_v I__2577 (
            .O(N__10758),
            .I(N__10752));
    Span4Mux_h I__2576 (
            .O(N__10755),
            .I(N__10749));
    Span4Mux_h I__2575 (
            .O(N__10752),
            .I(N__10746));
    Sp12to4 I__2574 (
            .O(N__10749),
            .I(N__10743));
    Sp12to4 I__2573 (
            .O(N__10746),
            .I(N__10738));
    Span12Mux_v I__2572 (
            .O(N__10743),
            .I(N__10738));
    Odrv12 I__2571 (
            .O(N__10738),
            .I(DRA_c_6));
    InMux I__2570 (
            .O(N__10735),
            .I(N__10732));
    LocalMux I__2569 (
            .O(N__10732),
            .I(N__10727));
    InMux I__2568 (
            .O(N__10731),
            .I(N__10724));
    InMux I__2567 (
            .O(N__10730),
            .I(N__10721));
    Span4Mux_h I__2566 (
            .O(N__10727),
            .I(N__10715));
    LocalMux I__2565 (
            .O(N__10724),
            .I(N__10715));
    LocalMux I__2564 (
            .O(N__10721),
            .I(N__10712));
    InMux I__2563 (
            .O(N__10720),
            .I(N__10709));
    Span4Mux_v I__2562 (
            .O(N__10715),
            .I(N__10706));
    Sp12to4 I__2561 (
            .O(N__10712),
            .I(N__10701));
    LocalMux I__2560 (
            .O(N__10709),
            .I(N__10701));
    Sp12to4 I__2559 (
            .O(N__10706),
            .I(N__10698));
    Span12Mux_v I__2558 (
            .O(N__10701),
            .I(N__10695));
    Span12Mux_h I__2557 (
            .O(N__10698),
            .I(N__10692));
    Span12Mux_h I__2556 (
            .O(N__10695),
            .I(N__10689));
    Odrv12 I__2555 (
            .O(N__10692),
            .I(DRA_c_7));
    Odrv12 I__2554 (
            .O(N__10689),
            .I(DRA_c_7));
    InMux I__2553 (
            .O(N__10684),
            .I(N__10681));
    LocalMux I__2552 (
            .O(N__10681),
            .I(N__10678));
    Odrv4 I__2551 (
            .O(N__10678),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2550 (
            .O(N__10675),
            .I(N__10668));
    InMux I__2549 (
            .O(N__10674),
            .I(N__10668));
    InMux I__2548 (
            .O(N__10673),
            .I(N__10664));
    LocalMux I__2547 (
            .O(N__10668),
            .I(N__10661));
    InMux I__2546 (
            .O(N__10667),
            .I(N__10658));
    LocalMux I__2545 (
            .O(N__10664),
            .I(N__10655));
    Span4Mux_v I__2544 (
            .O(N__10661),
            .I(N__10652));
    LocalMux I__2543 (
            .O(N__10658),
            .I(N__10649));
    Span12Mux_v I__2542 (
            .O(N__10655),
            .I(N__10646));
    Span4Mux_h I__2541 (
            .O(N__10652),
            .I(N__10641));
    Span4Mux_v I__2540 (
            .O(N__10649),
            .I(N__10641));
    Span12Mux_h I__2539 (
            .O(N__10646),
            .I(N__10638));
    Sp12to4 I__2538 (
            .O(N__10641),
            .I(N__10635));
    Odrv12 I__2537 (
            .O(N__10638),
            .I(DRA_c_8));
    Odrv12 I__2536 (
            .O(N__10635),
            .I(DRA_c_8));
    InMux I__2535 (
            .O(N__10630),
            .I(N__10627));
    LocalMux I__2534 (
            .O(N__10627),
            .I(N__10624));
    Span4Mux_v I__2533 (
            .O(N__10624),
            .I(N__10621));
    Odrv4 I__2532 (
            .O(N__10621),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2531 (
            .O(N__10618),
            .I(N__10606));
    InMux I__2530 (
            .O(N__10617),
            .I(N__10606));
    InMux I__2529 (
            .O(N__10616),
            .I(N__10606));
    InMux I__2528 (
            .O(N__10615),
            .I(N__10603));
    InMux I__2527 (
            .O(N__10614),
            .I(N__10600));
    InMux I__2526 (
            .O(N__10613),
            .I(N__10588));
    LocalMux I__2525 (
            .O(N__10606),
            .I(N__10584));
    LocalMux I__2524 (
            .O(N__10603),
            .I(N__10579));
    LocalMux I__2523 (
            .O(N__10600),
            .I(N__10579));
    InMux I__2522 (
            .O(N__10599),
            .I(N__10576));
    InMux I__2521 (
            .O(N__10598),
            .I(N__10573));
    InMux I__2520 (
            .O(N__10597),
            .I(N__10570));
    InMux I__2519 (
            .O(N__10596),
            .I(N__10562));
    InMux I__2518 (
            .O(N__10595),
            .I(N__10562));
    InMux I__2517 (
            .O(N__10594),
            .I(N__10562));
    InMux I__2516 (
            .O(N__10593),
            .I(N__10559));
    InMux I__2515 (
            .O(N__10592),
            .I(N__10556));
    CascadeMux I__2514 (
            .O(N__10591),
            .I(N__10552));
    LocalMux I__2513 (
            .O(N__10588),
            .I(N__10549));
    InMux I__2512 (
            .O(N__10587),
            .I(N__10546));
    Span4Mux_v I__2511 (
            .O(N__10584),
            .I(N__10535));
    Span4Mux_v I__2510 (
            .O(N__10579),
            .I(N__10535));
    LocalMux I__2509 (
            .O(N__10576),
            .I(N__10535));
    LocalMux I__2508 (
            .O(N__10573),
            .I(N__10535));
    LocalMux I__2507 (
            .O(N__10570),
            .I(N__10535));
    InMux I__2506 (
            .O(N__10569),
            .I(N__10532));
    LocalMux I__2505 (
            .O(N__10562),
            .I(N__10527));
    LocalMux I__2504 (
            .O(N__10559),
            .I(N__10522));
    LocalMux I__2503 (
            .O(N__10556),
            .I(N__10522));
    InMux I__2502 (
            .O(N__10555),
            .I(N__10518));
    InMux I__2501 (
            .O(N__10552),
            .I(N__10515));
    Span4Mux_v I__2500 (
            .O(N__10549),
            .I(N__10512));
    LocalMux I__2499 (
            .O(N__10546),
            .I(N__10509));
    Span4Mux_v I__2498 (
            .O(N__10535),
            .I(N__10506));
    LocalMux I__2497 (
            .O(N__10532),
            .I(N__10503));
    InMux I__2496 (
            .O(N__10531),
            .I(N__10498));
    InMux I__2495 (
            .O(N__10530),
            .I(N__10498));
    Span4Mux_h I__2494 (
            .O(N__10527),
            .I(N__10493));
    Span4Mux_v I__2493 (
            .O(N__10522),
            .I(N__10493));
    InMux I__2492 (
            .O(N__10521),
            .I(N__10490));
    LocalMux I__2491 (
            .O(N__10518),
            .I(N__10485));
    LocalMux I__2490 (
            .O(N__10515),
            .I(N__10485));
    Span4Mux_h I__2489 (
            .O(N__10512),
            .I(N__10480));
    Span4Mux_v I__2488 (
            .O(N__10509),
            .I(N__10480));
    Span4Mux_h I__2487 (
            .O(N__10506),
            .I(N__10475));
    Span4Mux_v I__2486 (
            .O(N__10503),
            .I(N__10475));
    LocalMux I__2485 (
            .O(N__10498),
            .I(N__10468));
    Sp12to4 I__2484 (
            .O(N__10493),
            .I(N__10468));
    LocalMux I__2483 (
            .O(N__10490),
            .I(N__10468));
    Sp12to4 I__2482 (
            .O(N__10485),
            .I(N__10465));
    Sp12to4 I__2481 (
            .O(N__10480),
            .I(N__10460));
    Sp12to4 I__2480 (
            .O(N__10475),
            .I(N__10460));
    Span12Mux_h I__2479 (
            .O(N__10468),
            .I(N__10457));
    Span12Mux_v I__2478 (
            .O(N__10465),
            .I(N__10454));
    Span12Mux_h I__2477 (
            .O(N__10460),
            .I(N__10451));
    Span12Mux_v I__2476 (
            .O(N__10457),
            .I(N__10446));
    Span12Mux_h I__2475 (
            .O(N__10454),
            .I(N__10446));
    Span12Mux_v I__2474 (
            .O(N__10451),
            .I(N__10443));
    Odrv12 I__2473 (
            .O(N__10446),
            .I(AGNUS_REV_c));
    Odrv12 I__2472 (
            .O(N__10443),
            .I(AGNUS_REV_c));
    InMux I__2471 (
            .O(N__10438),
            .I(N__10435));
    LocalMux I__2470 (
            .O(N__10435),
            .I(N__10432));
    Odrv12 I__2469 (
            .O(N__10432),
            .I(RAS0n_c));
    InMux I__2468 (
            .O(N__10429),
            .I(N__10425));
    InMux I__2467 (
            .O(N__10428),
            .I(N__10422));
    LocalMux I__2466 (
            .O(N__10425),
            .I(N__10418));
    LocalMux I__2465 (
            .O(N__10422),
            .I(N__10415));
    InMux I__2464 (
            .O(N__10421),
            .I(N__10412));
    Span4Mux_v I__2463 (
            .O(N__10418),
            .I(N__10409));
    Span4Mux_v I__2462 (
            .O(N__10415),
            .I(N__10404));
    LocalMux I__2461 (
            .O(N__10412),
            .I(N__10404));
    Span4Mux_v I__2460 (
            .O(N__10409),
            .I(N__10398));
    Span4Mux_v I__2459 (
            .O(N__10404),
            .I(N__10398));
    InMux I__2458 (
            .O(N__10403),
            .I(N__10395));
    Sp12to4 I__2457 (
            .O(N__10398),
            .I(N__10392));
    LocalMux I__2456 (
            .O(N__10395),
            .I(N__10389));
    Span12Mux_h I__2455 (
            .O(N__10392),
            .I(N__10386));
    Span12Mux_v I__2454 (
            .O(N__10389),
            .I(N__10383));
    Span12Mux_v I__2453 (
            .O(N__10386),
            .I(N__10380));
    Span12Mux_v I__2452 (
            .O(N__10383),
            .I(N__10377));
    Odrv12 I__2451 (
            .O(N__10380),
            .I(DRA_c_9));
    Odrv12 I__2450 (
            .O(N__10377),
            .I(DRA_c_9));
    InMux I__2449 (
            .O(N__10372),
            .I(N__10369));
    LocalMux I__2448 (
            .O(N__10369),
            .I(N__10366));
    Span4Mux_h I__2447 (
            .O(N__10366),
            .I(N__10363));
    Span4Mux_h I__2446 (
            .O(N__10363),
            .I(N__10360));
    Odrv4 I__2445 (
            .O(N__10360),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    ClkMux I__2444 (
            .O(N__10357),
            .I(N__10333));
    ClkMux I__2443 (
            .O(N__10356),
            .I(N__10333));
    ClkMux I__2442 (
            .O(N__10355),
            .I(N__10333));
    ClkMux I__2441 (
            .O(N__10354),
            .I(N__10333));
    ClkMux I__2440 (
            .O(N__10353),
            .I(N__10333));
    ClkMux I__2439 (
            .O(N__10352),
            .I(N__10333));
    ClkMux I__2438 (
            .O(N__10351),
            .I(N__10333));
    ClkMux I__2437 (
            .O(N__10350),
            .I(N__10333));
    GlobalMux I__2436 (
            .O(N__10333),
            .I(N__10330));
    gio2CtrlBuf I__2435 (
            .O(N__10330),
            .I(C3_c_g));
    CEMux I__2434 (
            .O(N__10327),
            .I(N__10285));
    CEMux I__2433 (
            .O(N__10326),
            .I(N__10285));
    CEMux I__2432 (
            .O(N__10325),
            .I(N__10285));
    CEMux I__2431 (
            .O(N__10324),
            .I(N__10285));
    CEMux I__2430 (
            .O(N__10323),
            .I(N__10285));
    CEMux I__2429 (
            .O(N__10322),
            .I(N__10285));
    CEMux I__2428 (
            .O(N__10321),
            .I(N__10285));
    CEMux I__2427 (
            .O(N__10320),
            .I(N__10285));
    CEMux I__2426 (
            .O(N__10319),
            .I(N__10285));
    CEMux I__2425 (
            .O(N__10318),
            .I(N__10285));
    CEMux I__2424 (
            .O(N__10317),
            .I(N__10285));
    CEMux I__2423 (
            .O(N__10316),
            .I(N__10285));
    CEMux I__2422 (
            .O(N__10315),
            .I(N__10285));
    CEMux I__2421 (
            .O(N__10314),
            .I(N__10285));
    GlobalMux I__2420 (
            .O(N__10285),
            .I(N__10282));
    gio2CtrlBuf I__2419 (
            .O(N__10282),
            .I(DBRn_c_i_0_g));
    InMux I__2418 (
            .O(N__10279),
            .I(N__10272));
    InMux I__2417 (
            .O(N__10278),
            .I(N__10269));
    InMux I__2416 (
            .O(N__10277),
            .I(N__10266));
    InMux I__2415 (
            .O(N__10276),
            .I(N__10261));
    InMux I__2414 (
            .O(N__10275),
            .I(N__10261));
    LocalMux I__2413 (
            .O(N__10272),
            .I(N__10247));
    LocalMux I__2412 (
            .O(N__10269),
            .I(N__10240));
    LocalMux I__2411 (
            .O(N__10266),
            .I(N__10229));
    LocalMux I__2410 (
            .O(N__10261),
            .I(N__10226));
    SRMux I__2409 (
            .O(N__10260),
            .I(N__10132));
    SRMux I__2408 (
            .O(N__10259),
            .I(N__10132));
    SRMux I__2407 (
            .O(N__10258),
            .I(N__10132));
    SRMux I__2406 (
            .O(N__10257),
            .I(N__10132));
    SRMux I__2405 (
            .O(N__10256),
            .I(N__10132));
    SRMux I__2404 (
            .O(N__10255),
            .I(N__10132));
    SRMux I__2403 (
            .O(N__10254),
            .I(N__10132));
    SRMux I__2402 (
            .O(N__10253),
            .I(N__10132));
    SRMux I__2401 (
            .O(N__10252),
            .I(N__10132));
    SRMux I__2400 (
            .O(N__10251),
            .I(N__10132));
    SRMux I__2399 (
            .O(N__10250),
            .I(N__10132));
    Glb2LocalMux I__2398 (
            .O(N__10247),
            .I(N__10132));
    SRMux I__2397 (
            .O(N__10246),
            .I(N__10132));
    SRMux I__2396 (
            .O(N__10245),
            .I(N__10132));
    SRMux I__2395 (
            .O(N__10244),
            .I(N__10132));
    SRMux I__2394 (
            .O(N__10243),
            .I(N__10132));
    Glb2LocalMux I__2393 (
            .O(N__10240),
            .I(N__10132));
    SRMux I__2392 (
            .O(N__10239),
            .I(N__10132));
    SRMux I__2391 (
            .O(N__10238),
            .I(N__10132));
    SRMux I__2390 (
            .O(N__10237),
            .I(N__10132));
    SRMux I__2389 (
            .O(N__10236),
            .I(N__10132));
    SRMux I__2388 (
            .O(N__10235),
            .I(N__10132));
    SRMux I__2387 (
            .O(N__10234),
            .I(N__10132));
    SRMux I__2386 (
            .O(N__10233),
            .I(N__10132));
    SRMux I__2385 (
            .O(N__10232),
            .I(N__10132));
    Glb2LocalMux I__2384 (
            .O(N__10229),
            .I(N__10132));
    Glb2LocalMux I__2383 (
            .O(N__10226),
            .I(N__10132));
    SRMux I__2382 (
            .O(N__10225),
            .I(N__10132));
    SRMux I__2381 (
            .O(N__10224),
            .I(N__10132));
    SRMux I__2380 (
            .O(N__10223),
            .I(N__10132));
    SRMux I__2379 (
            .O(N__10222),
            .I(N__10132));
    SRMux I__2378 (
            .O(N__10221),
            .I(N__10132));
    SRMux I__2377 (
            .O(N__10220),
            .I(N__10132));
    SRMux I__2376 (
            .O(N__10219),
            .I(N__10132));
    SRMux I__2375 (
            .O(N__10218),
            .I(N__10132));
    SRMux I__2374 (
            .O(N__10217),
            .I(N__10132));
    SRMux I__2373 (
            .O(N__10216),
            .I(N__10132));
    SRMux I__2372 (
            .O(N__10215),
            .I(N__10132));
    SRMux I__2371 (
            .O(N__10214),
            .I(N__10132));
    SRMux I__2370 (
            .O(N__10213),
            .I(N__10132));
    GlobalMux I__2369 (
            .O(N__10132),
            .I(N__10129));
    gio2CtrlBuf I__2368 (
            .O(N__10129),
            .I(RESETn_c_i_g));
    InMux I__2367 (
            .O(N__10126),
            .I(N__10123));
    LocalMux I__2366 (
            .O(N__10123),
            .I(N__10120));
    Sp12to4 I__2365 (
            .O(N__10120),
            .I(N__10116));
    InMux I__2364 (
            .O(N__10119),
            .I(N__10113));
    Span12Mux_v I__2363 (
            .O(N__10116),
            .I(N__10110));
    LocalMux I__2362 (
            .O(N__10113),
            .I(N__10107));
    Span12Mux_h I__2361 (
            .O(N__10110),
            .I(N__10103));
    Span4Mux_v I__2360 (
            .O(N__10107),
            .I(N__10100));
    InMux I__2359 (
            .O(N__10106),
            .I(N__10097));
    Odrv12 I__2358 (
            .O(N__10103),
            .I(REG_CYCLEm));
    Odrv4 I__2357 (
            .O(N__10100),
            .I(REG_CYCLEm));
    LocalMux I__2356 (
            .O(N__10097),
            .I(REG_CYCLEm));
    InMux I__2355 (
            .O(N__10090),
            .I(N__10087));
    LocalMux I__2354 (
            .O(N__10087),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2353 (
            .O(N__10084),
            .I(N__10081));
    LocalMux I__2352 (
            .O(N__10081),
            .I(N__10077));
    InMux I__2351 (
            .O(N__10080),
            .I(N__10074));
    Span4Mux_h I__2350 (
            .O(N__10077),
            .I(N__10069));
    LocalMux I__2349 (
            .O(N__10074),
            .I(N__10069));
    Span4Mux_v I__2348 (
            .O(N__10069),
            .I(N__10064));
    InMux I__2347 (
            .O(N__10068),
            .I(N__10061));
    InMux I__2346 (
            .O(N__10067),
            .I(N__10058));
    Span4Mux_v I__2345 (
            .O(N__10064),
            .I(N__10055));
    LocalMux I__2344 (
            .O(N__10061),
            .I(N__10050));
    LocalMux I__2343 (
            .O(N__10058),
            .I(N__10050));
    Sp12to4 I__2342 (
            .O(N__10055),
            .I(N__10045));
    Span12Mux_v I__2341 (
            .O(N__10050),
            .I(N__10045));
    Span12Mux_h I__2340 (
            .O(N__10045),
            .I(N__10042));
    Odrv12 I__2339 (
            .O(N__10042),
            .I(DRA_c_5));
    InMux I__2338 (
            .O(N__10039),
            .I(N__10033));
    InMux I__2337 (
            .O(N__10038),
            .I(N__10033));
    LocalMux I__2336 (
            .O(N__10033),
            .I(N__10030));
    Span4Mux_v I__2335 (
            .O(N__10030),
            .I(N__10027));
    Odrv4 I__2334 (
            .O(N__10027),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    CascadeMux I__2333 (
            .O(N__10024),
            .I(N__10021));
    InMux I__2332 (
            .O(N__10021),
            .I(N__10013));
    InMux I__2331 (
            .O(N__10020),
            .I(N__10013));
    InMux I__2330 (
            .O(N__10019),
            .I(N__10010));
    InMux I__2329 (
            .O(N__10018),
            .I(N__10007));
    LocalMux I__2328 (
            .O(N__10013),
            .I(N__10002));
    LocalMux I__2327 (
            .O(N__10010),
            .I(N__10002));
    LocalMux I__2326 (
            .O(N__10007),
            .I(N__9999));
    Span4Mux_v I__2325 (
            .O(N__10002),
            .I(N__9996));
    Sp12to4 I__2324 (
            .O(N__9999),
            .I(N__9993));
    Sp12to4 I__2323 (
            .O(N__9996),
            .I(N__9990));
    Span12Mux_v I__2322 (
            .O(N__9993),
            .I(N__9987));
    Span12Mux_h I__2321 (
            .O(N__9990),
            .I(N__9984));
    Span12Mux_h I__2320 (
            .O(N__9987),
            .I(N__9979));
    Span12Mux_v I__2319 (
            .O(N__9984),
            .I(N__9979));
    Odrv12 I__2318 (
            .O(N__9979),
            .I(DRA_c_2));
    InMux I__2317 (
            .O(N__9976),
            .I(N__9973));
    LocalMux I__2316 (
            .O(N__9973),
            .I(N__9970));
    Odrv4 I__2315 (
            .O(N__9970),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2314 (
            .O(N__9967),
            .I(N__9964));
    LocalMux I__2313 (
            .O(N__9964),
            .I(N__9961));
    Span4Mux_h I__2312 (
            .O(N__9961),
            .I(N__9958));
    Odrv4 I__2311 (
            .O(N__9958),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__2310 (
            .O(N__9955),
            .I(N__9950));
    InMux I__2309 (
            .O(N__9954),
            .I(N__9947));
    InMux I__2308 (
            .O(N__9953),
            .I(N__9943));
    LocalMux I__2307 (
            .O(N__9950),
            .I(N__9938));
    LocalMux I__2306 (
            .O(N__9947),
            .I(N__9938));
    InMux I__2305 (
            .O(N__9946),
            .I(N__9935));
    LocalMux I__2304 (
            .O(N__9943),
            .I(N__9932));
    Span4Mux_v I__2303 (
            .O(N__9938),
            .I(N__9925));
    LocalMux I__2302 (
            .O(N__9935),
            .I(N__9925));
    Span4Mux_v I__2301 (
            .O(N__9932),
            .I(N__9925));
    Sp12to4 I__2300 (
            .O(N__9925),
            .I(N__9922));
    Span12Mux_h I__2299 (
            .O(N__9922),
            .I(N__9919));
    Span12Mux_v I__2298 (
            .O(N__9919),
            .I(N__9916));
    Odrv12 I__2297 (
            .O(N__9916),
            .I(DRA_c_1));
    InMux I__2296 (
            .O(N__9913),
            .I(N__9910));
    LocalMux I__2295 (
            .O(N__9910),
            .I(N__9906));
    InMux I__2294 (
            .O(N__9909),
            .I(N__9903));
    Sp12to4 I__2293 (
            .O(N__9906),
            .I(N__9900));
    LocalMux I__2292 (
            .O(N__9903),
            .I(N__9897));
    Span12Mux_v I__2291 (
            .O(N__9900),
            .I(N__9894));
    Span12Mux_h I__2290 (
            .O(N__9897),
            .I(N__9891));
    Span12Mux_h I__2289 (
            .O(N__9894),
            .I(N__9888));
    Span12Mux_v I__2288 (
            .O(N__9891),
            .I(N__9885));
    Odrv12 I__2287 (
            .O(N__9888),
            .I(DRA_c_0));
    Odrv12 I__2286 (
            .O(N__9885),
            .I(DRA_c_0));
    InMux I__2285 (
            .O(N__9880),
            .I(N__9877));
    LocalMux I__2284 (
            .O(N__9877),
            .I(N__9874));
    Span4Mux_h I__2283 (
            .O(N__9874),
            .I(N__9871));
    Odrv4 I__2282 (
            .O(N__9871),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    IoInMux I__2281 (
            .O(N__9868),
            .I(N__9865));
    LocalMux I__2280 (
            .O(N__9865),
            .I(N__9862));
    Sp12to4 I__2279 (
            .O(N__9862),
            .I(N__9859));
    Span12Mux_h I__2278 (
            .O(N__9859),
            .I(N__9856));
    Span12Mux_v I__2277 (
            .O(N__9856),
            .I(N__9853));
    Odrv12 I__2276 (
            .O(N__9853),
            .I(N_57_i));
    CascadeMux I__2275 (
            .O(N__9850),
            .I(N__9846));
    IoInMux I__2274 (
            .O(N__9849),
            .I(N__9842));
    InMux I__2273 (
            .O(N__9846),
            .I(N__9839));
    InMux I__2272 (
            .O(N__9845),
            .I(N__9836));
    LocalMux I__2271 (
            .O(N__9842),
            .I(N__9831));
    LocalMux I__2270 (
            .O(N__9839),
            .I(N__9826));
    LocalMux I__2269 (
            .O(N__9836),
            .I(N__9826));
    InMux I__2268 (
            .O(N__9835),
            .I(N__9823));
    InMux I__2267 (
            .O(N__9834),
            .I(N__9820));
    Span12Mux_s2_v I__2266 (
            .O(N__9831),
            .I(N__9817));
    Span4Mux_v I__2265 (
            .O(N__9826),
            .I(N__9814));
    LocalMux I__2264 (
            .O(N__9823),
            .I(N__9809));
    LocalMux I__2263 (
            .O(N__9820),
            .I(N__9809));
    Span12Mux_v I__2262 (
            .O(N__9817),
            .I(N__9805));
    Span4Mux_h I__2261 (
            .O(N__9814),
            .I(N__9802));
    Span4Mux_v I__2260 (
            .O(N__9809),
            .I(N__9799));
    InMux I__2259 (
            .O(N__9808),
            .I(N__9796));
    Odrv12 I__2258 (
            .O(N__9805),
            .I(DBENn_c));
    Odrv4 I__2257 (
            .O(N__9802),
            .I(DBENn_c));
    Odrv4 I__2256 (
            .O(N__9799),
            .I(DBENn_c));
    LocalMux I__2255 (
            .O(N__9796),
            .I(DBENn_c));
    CascadeMux I__2254 (
            .O(N__9787),
            .I(N__9784));
    InMux I__2253 (
            .O(N__9784),
            .I(N__9778));
    InMux I__2252 (
            .O(N__9783),
            .I(N__9775));
    InMux I__2251 (
            .O(N__9782),
            .I(N__9771));
    InMux I__2250 (
            .O(N__9781),
            .I(N__9767));
    LocalMux I__2249 (
            .O(N__9778),
            .I(N__9764));
    LocalMux I__2248 (
            .O(N__9775),
            .I(N__9761));
    InMux I__2247 (
            .O(N__9774),
            .I(N__9758));
    LocalMux I__2246 (
            .O(N__9771),
            .I(N__9754));
    InMux I__2245 (
            .O(N__9770),
            .I(N__9751));
    LocalMux I__2244 (
            .O(N__9767),
            .I(N__9748));
    Span4Mux_h I__2243 (
            .O(N__9764),
            .I(N__9743));
    Span4Mux_v I__2242 (
            .O(N__9761),
            .I(N__9743));
    LocalMux I__2241 (
            .O(N__9758),
            .I(N__9740));
    InMux I__2240 (
            .O(N__9757),
            .I(N__9735));
    Span4Mux_v I__2239 (
            .O(N__9754),
            .I(N__9732));
    LocalMux I__2238 (
            .O(N__9751),
            .I(N__9729));
    Span4Mux_v I__2237 (
            .O(N__9748),
            .I(N__9726));
    Span4Mux_v I__2236 (
            .O(N__9743),
            .I(N__9721));
    Span4Mux_v I__2235 (
            .O(N__9740),
            .I(N__9721));
    InMux I__2234 (
            .O(N__9739),
            .I(N__9718));
    InMux I__2233 (
            .O(N__9738),
            .I(N__9715));
    LocalMux I__2232 (
            .O(N__9735),
            .I(N__9712));
    Span4Mux_h I__2231 (
            .O(N__9732),
            .I(N__9707));
    Span4Mux_h I__2230 (
            .O(N__9729),
            .I(N__9707));
    Odrv4 I__2229 (
            .O(N__9726),
            .I(DMA_CYCLEm));
    Odrv4 I__2228 (
            .O(N__9721),
            .I(DMA_CYCLEm));
    LocalMux I__2227 (
            .O(N__9718),
            .I(DMA_CYCLEm));
    LocalMux I__2226 (
            .O(N__9715),
            .I(DMA_CYCLEm));
    Odrv12 I__2225 (
            .O(N__9712),
            .I(DMA_CYCLEm));
    Odrv4 I__2224 (
            .O(N__9707),
            .I(DMA_CYCLEm));
    IoInMux I__2223 (
            .O(N__9694),
            .I(N__9691));
    LocalMux I__2222 (
            .O(N__9691),
            .I(N__9688));
    Span4Mux_s2_h I__2221 (
            .O(N__9688),
            .I(N__9685));
    Span4Mux_v I__2220 (
            .O(N__9685),
            .I(N__9682));
    Span4Mux_v I__2219 (
            .O(N__9682),
            .I(N__9679));
    Sp12to4 I__2218 (
            .O(N__9679),
            .I(N__9676));
    Odrv12 I__2217 (
            .O(N__9676),
            .I(N_59_i));
    InMux I__2216 (
            .O(N__9673),
            .I(N__9670));
    LocalMux I__2215 (
            .O(N__9670),
            .I(\U712_BYTE_ENABLE.N_557 ));
    CascadeMux I__2214 (
            .O(N__9667),
            .I(N__9660));
    InMux I__2213 (
            .O(N__9666),
            .I(N__9655));
    CascadeMux I__2212 (
            .O(N__9665),
            .I(N__9652));
    CascadeMux I__2211 (
            .O(N__9664),
            .I(N__9649));
    CascadeMux I__2210 (
            .O(N__9663),
            .I(N__9645));
    InMux I__2209 (
            .O(N__9660),
            .I(N__9640));
    CascadeMux I__2208 (
            .O(N__9659),
            .I(N__9637));
    CascadeMux I__2207 (
            .O(N__9658),
            .I(N__9630));
    LocalMux I__2206 (
            .O(N__9655),
            .I(N__9625));
    InMux I__2205 (
            .O(N__9652),
            .I(N__9622));
    InMux I__2204 (
            .O(N__9649),
            .I(N__9617));
    InMux I__2203 (
            .O(N__9648),
            .I(N__9613));
    InMux I__2202 (
            .O(N__9645),
            .I(N__9606));
    InMux I__2201 (
            .O(N__9644),
            .I(N__9606));
    InMux I__2200 (
            .O(N__9643),
            .I(N__9606));
    LocalMux I__2199 (
            .O(N__9640),
            .I(N__9603));
    InMux I__2198 (
            .O(N__9637),
            .I(N__9600));
    InMux I__2197 (
            .O(N__9636),
            .I(N__9597));
    InMux I__2196 (
            .O(N__9635),
            .I(N__9592));
    InMux I__2195 (
            .O(N__9634),
            .I(N__9592));
    InMux I__2194 (
            .O(N__9633),
            .I(N__9589));
    InMux I__2193 (
            .O(N__9630),
            .I(N__9586));
    InMux I__2192 (
            .O(N__9629),
            .I(N__9580));
    InMux I__2191 (
            .O(N__9628),
            .I(N__9580));
    Span4Mux_v I__2190 (
            .O(N__9625),
            .I(N__9572));
    LocalMux I__2189 (
            .O(N__9622),
            .I(N__9572));
    InMux I__2188 (
            .O(N__9621),
            .I(N__9567));
    InMux I__2187 (
            .O(N__9620),
            .I(N__9567));
    LocalMux I__2186 (
            .O(N__9617),
            .I(N__9564));
    InMux I__2185 (
            .O(N__9616),
            .I(N__9561));
    LocalMux I__2184 (
            .O(N__9613),
            .I(N__9556));
    LocalMux I__2183 (
            .O(N__9606),
            .I(N__9556));
    Span4Mux_v I__2182 (
            .O(N__9603),
            .I(N__9547));
    LocalMux I__2181 (
            .O(N__9600),
            .I(N__9547));
    LocalMux I__2180 (
            .O(N__9597),
            .I(N__9547));
    LocalMux I__2179 (
            .O(N__9592),
            .I(N__9547));
    LocalMux I__2178 (
            .O(N__9589),
            .I(N__9544));
    LocalMux I__2177 (
            .O(N__9586),
            .I(N__9541));
    InMux I__2176 (
            .O(N__9585),
            .I(N__9538));
    LocalMux I__2175 (
            .O(N__9580),
            .I(N__9535));
    InMux I__2174 (
            .O(N__9579),
            .I(N__9532));
    InMux I__2173 (
            .O(N__9578),
            .I(N__9527));
    InMux I__2172 (
            .O(N__9577),
            .I(N__9527));
    Span4Mux_v I__2171 (
            .O(N__9572),
            .I(N__9520));
    LocalMux I__2170 (
            .O(N__9567),
            .I(N__9520));
    Span4Mux_v I__2169 (
            .O(N__9564),
            .I(N__9520));
    LocalMux I__2168 (
            .O(N__9561),
            .I(N__9513));
    Span4Mux_h I__2167 (
            .O(N__9556),
            .I(N__9513));
    Span4Mux_v I__2166 (
            .O(N__9547),
            .I(N__9513));
    Span4Mux_v I__2165 (
            .O(N__9544),
            .I(N__9506));
    Span4Mux_h I__2164 (
            .O(N__9541),
            .I(N__9506));
    LocalMux I__2163 (
            .O(N__9538),
            .I(N__9506));
    Span12Mux_h I__2162 (
            .O(N__9535),
            .I(N__9501));
    LocalMux I__2161 (
            .O(N__9532),
            .I(N__9501));
    LocalMux I__2160 (
            .O(N__9527),
            .I(CPU_CYCLEm));
    Odrv4 I__2159 (
            .O(N__9520),
            .I(CPU_CYCLEm));
    Odrv4 I__2158 (
            .O(N__9513),
            .I(CPU_CYCLEm));
    Odrv4 I__2157 (
            .O(N__9506),
            .I(CPU_CYCLEm));
    Odrv12 I__2156 (
            .O(N__9501),
            .I(CPU_CYCLEm));
    InMux I__2155 (
            .O(N__9490),
            .I(N__9487));
    LocalMux I__2154 (
            .O(N__9487),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2153 (
            .O(N__9484),
            .I(N__9481));
    LocalMux I__2152 (
            .O(N__9481),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2151 (
            .O(N__9478),
            .I(N__9475));
    LocalMux I__2150 (
            .O(N__9475),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2149 (
            .O(N__9472),
            .I(N__9469));
    LocalMux I__2148 (
            .O(N__9469),
            .I(N__9466));
    Span4Mux_h I__2147 (
            .O(N__9466),
            .I(N__9463));
    Odrv4 I__2146 (
            .O(N__9463),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__2145 (
            .O(N__9460),
            .I(N__9457));
    LocalMux I__2144 (
            .O(N__9457),
            .I(N__9452));
    InMux I__2143 (
            .O(N__9456),
            .I(N__9449));
    InMux I__2142 (
            .O(N__9455),
            .I(N__9445));
    Span4Mux_h I__2141 (
            .O(N__9452),
            .I(N__9440));
    LocalMux I__2140 (
            .O(N__9449),
            .I(N__9440));
    InMux I__2139 (
            .O(N__9448),
            .I(N__9437));
    LocalMux I__2138 (
            .O(N__9445),
            .I(N__9430));
    Sp12to4 I__2137 (
            .O(N__9440),
            .I(N__9430));
    LocalMux I__2136 (
            .O(N__9437),
            .I(N__9430));
    Span12Mux_v I__2135 (
            .O(N__9430),
            .I(N__9427));
    Span12Mux_h I__2134 (
            .O(N__9427),
            .I(N__9424));
    Odrv12 I__2133 (
            .O(N__9424),
            .I(DRA_c_3));
    InMux I__2132 (
            .O(N__9421),
            .I(N__9418));
    LocalMux I__2131 (
            .O(N__9418),
            .I(N__9415));
    Span4Mux_h I__2130 (
            .O(N__9415),
            .I(N__9412));
    Odrv4 I__2129 (
            .O(N__9412),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__2128 (
            .O(N__9409),
            .I(N__9402));
    InMux I__2127 (
            .O(N__9408),
            .I(N__9402));
    InMux I__2126 (
            .O(N__9407),
            .I(N__9399));
    LocalMux I__2125 (
            .O(N__9402),
            .I(N__9395));
    LocalMux I__2124 (
            .O(N__9399),
            .I(N__9392));
    InMux I__2123 (
            .O(N__9398),
            .I(N__9389));
    Span4Mux_v I__2122 (
            .O(N__9395),
            .I(N__9382));
    Span4Mux_h I__2121 (
            .O(N__9392),
            .I(N__9382));
    LocalMux I__2120 (
            .O(N__9389),
            .I(N__9382));
    Span4Mux_v I__2119 (
            .O(N__9382),
            .I(N__9379));
    Span4Mux_v I__2118 (
            .O(N__9379),
            .I(N__9376));
    Sp12to4 I__2117 (
            .O(N__9376),
            .I(N__9373));
    Span12Mux_h I__2116 (
            .O(N__9373),
            .I(N__9370));
    Odrv12 I__2115 (
            .O(N__9370),
            .I(DRA_c_4));
    InMux I__2114 (
            .O(N__9367),
            .I(N__9364));
    LocalMux I__2113 (
            .O(N__9364),
            .I(N__9361));
    Odrv4 I__2112 (
            .O(N__9361),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    IoInMux I__2111 (
            .O(N__9358),
            .I(N__9355));
    LocalMux I__2110 (
            .O(N__9355),
            .I(N__9352));
    Span4Mux_s2_v I__2109 (
            .O(N__9352),
            .I(N__9349));
    Span4Mux_v I__2108 (
            .O(N__9349),
            .I(N__9346));
    Sp12to4 I__2107 (
            .O(N__9346),
            .I(N__9343));
    Odrv12 I__2106 (
            .O(N__9343),
            .I(un1_UDSn_i_0_0));
    InMux I__2105 (
            .O(N__9340),
            .I(N__9334));
    InMux I__2104 (
            .O(N__9339),
            .I(N__9334));
    LocalMux I__2103 (
            .O(N__9334),
            .I(N__9331));
    Span4Mux_v I__2102 (
            .O(N__9331),
            .I(N__9328));
    Span4Mux_h I__2101 (
            .O(N__9328),
            .I(N__9325));
    Span4Mux_v I__2100 (
            .O(N__9325),
            .I(N__9321));
    InMux I__2099 (
            .O(N__9324),
            .I(N__9318));
    Odrv4 I__2098 (
            .O(N__9321),
            .I(DS_ENm));
    LocalMux I__2097 (
            .O(N__9318),
            .I(DS_ENm));
    IoInMux I__2096 (
            .O(N__9313),
            .I(N__9310));
    LocalMux I__2095 (
            .O(N__9310),
            .I(N__9307));
    Span12Mux_s6_v I__2094 (
            .O(N__9307),
            .I(N__9304));
    Odrv12 I__2093 (
            .O(N__9304),
            .I(un1_LDSn_i_0_0));
    CascadeMux I__2092 (
            .O(N__9301),
            .I(N__9298));
    InMux I__2091 (
            .O(N__9298),
            .I(N__9295));
    LocalMux I__2090 (
            .O(N__9295),
            .I(N__9292));
    Odrv12 I__2089 (
            .O(N__9292),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2088 (
            .O(N__9289),
            .I(N__9286));
    LocalMux I__2087 (
            .O(N__9286),
            .I(N__9282));
    InMux I__2086 (
            .O(N__9285),
            .I(N__9279));
    Odrv12 I__2085 (
            .O(N__9282),
            .I(DBRn_c_i));
    LocalMux I__2084 (
            .O(N__9279),
            .I(DBRn_c_i));
    InMux I__2083 (
            .O(N__9274),
            .I(N__9271));
    LocalMux I__2082 (
            .O(N__9271),
            .I(N__9267));
    InMux I__2081 (
            .O(N__9270),
            .I(N__9264));
    Span4Mux_h I__2080 (
            .O(N__9267),
            .I(N__9261));
    LocalMux I__2079 (
            .O(N__9264),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    Odrv4 I__2078 (
            .O(N__9261),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    IoInMux I__2077 (
            .O(N__9256),
            .I(N__9253));
    LocalMux I__2076 (
            .O(N__9253),
            .I(N__9250));
    IoSpan4Mux I__2075 (
            .O(N__9250),
            .I(N__9247));
    Span4Mux_s1_h I__2074 (
            .O(N__9247),
            .I(N__9244));
    Sp12to4 I__2073 (
            .O(N__9244),
            .I(N__9241));
    Span12Mux_h I__2072 (
            .O(N__9241),
            .I(N__9238));
    Span12Mux_v I__2071 (
            .O(N__9238),
            .I(N__9235));
    Odrv12 I__2070 (
            .O(N__9235),
            .I(N_58_i));
    CascadeMux I__2069 (
            .O(N__9232),
            .I(N__9229));
    InMux I__2068 (
            .O(N__9229),
            .I(N__9225));
    InMux I__2067 (
            .O(N__9228),
            .I(N__9222));
    LocalMux I__2066 (
            .O(N__9225),
            .I(N__9219));
    LocalMux I__2065 (
            .O(N__9222),
            .I(N__9216));
    Odrv4 I__2064 (
            .O(N__9219),
            .I(\U712_BYTE_ENABLE.N_410 ));
    Odrv4 I__2063 (
            .O(N__9216),
            .I(\U712_BYTE_ENABLE.N_410 ));
    CascadeMux I__2062 (
            .O(N__9211),
            .I(N__9208));
    InMux I__2061 (
            .O(N__9208),
            .I(N__9205));
    LocalMux I__2060 (
            .O(N__9205),
            .I(\U712_BYTE_ENABLE.N_559 ));
    IoInMux I__2059 (
            .O(N__9202),
            .I(N__9199));
    LocalMux I__2058 (
            .O(N__9199),
            .I(N__9196));
    IoSpan4Mux I__2057 (
            .O(N__9196),
            .I(N__9193));
    Span4Mux_s3_v I__2056 (
            .O(N__9193),
            .I(N__9190));
    Odrv4 I__2055 (
            .O(N__9190),
            .I(N_129_i));
    IoInMux I__2054 (
            .O(N__9187),
            .I(N__9184));
    LocalMux I__2053 (
            .O(N__9184),
            .I(N__9181));
    IoSpan4Mux I__2052 (
            .O(N__9181),
            .I(N__9178));
    Sp12to4 I__2051 (
            .O(N__9178),
            .I(N__9175));
    Span12Mux_s7_v I__2050 (
            .O(N__9175),
            .I(N__9172));
    Odrv12 I__2049 (
            .O(N__9172),
            .I(CASn_c));
    InMux I__2048 (
            .O(N__9169),
            .I(N__9165));
    InMux I__2047 (
            .O(N__9168),
            .I(N__9162));
    LocalMux I__2046 (
            .O(N__9165),
            .I(N__9155));
    LocalMux I__2045 (
            .O(N__9162),
            .I(N__9155));
    CascadeMux I__2044 (
            .O(N__9161),
            .I(N__9152));
    InMux I__2043 (
            .O(N__9160),
            .I(N__9149));
    Span4Mux_h I__2042 (
            .O(N__9155),
            .I(N__9144));
    InMux I__2041 (
            .O(N__9152),
            .I(N__9141));
    LocalMux I__2040 (
            .O(N__9149),
            .I(N__9138));
    InMux I__2039 (
            .O(N__9148),
            .I(N__9133));
    InMux I__2038 (
            .O(N__9147),
            .I(N__9133));
    Span4Mux_h I__2037 (
            .O(N__9144),
            .I(N__9130));
    LocalMux I__2036 (
            .O(N__9141),
            .I(N__9123));
    Span4Mux_v I__2035 (
            .O(N__9138),
            .I(N__9123));
    LocalMux I__2034 (
            .O(N__9133),
            .I(N__9123));
    Odrv4 I__2033 (
            .O(N__9130),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    Odrv4 I__2032 (
            .O(N__9123),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    IoInMux I__2031 (
            .O(N__9118),
            .I(N__9115));
    LocalMux I__2030 (
            .O(N__9115),
            .I(N__9112));
    IoSpan4Mux I__2029 (
            .O(N__9112),
            .I(N__9109));
    Sp12to4 I__2028 (
            .O(N__9109),
            .I(N__9106));
    Span12Mux_s9_v I__2027 (
            .O(N__9106),
            .I(N__9103));
    Odrv12 I__2026 (
            .O(N__9103),
            .I(RASn_c));
    InMux I__2025 (
            .O(N__9100),
            .I(N__9097));
    LocalMux I__2024 (
            .O(N__9097),
            .I(N__9094));
    Span12Mux_h I__2023 (
            .O(N__9094),
            .I(N__9091));
    Odrv12 I__2022 (
            .O(N__9091),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    InMux I__2021 (
            .O(N__9088),
            .I(N__9083));
    CascadeMux I__2020 (
            .O(N__9087),
            .I(N__9080));
    CascadeMux I__2019 (
            .O(N__9086),
            .I(N__9077));
    LocalMux I__2018 (
            .O(N__9083),
            .I(N__9065));
    InMux I__2017 (
            .O(N__9080),
            .I(N__9062));
    InMux I__2016 (
            .O(N__9077),
            .I(N__9059));
    InMux I__2015 (
            .O(N__9076),
            .I(N__9052));
    InMux I__2014 (
            .O(N__9075),
            .I(N__9052));
    InMux I__2013 (
            .O(N__9074),
            .I(N__9052));
    InMux I__2012 (
            .O(N__9073),
            .I(N__9047));
    InMux I__2011 (
            .O(N__9072),
            .I(N__9044));
    InMux I__2010 (
            .O(N__9071),
            .I(N__9039));
    InMux I__2009 (
            .O(N__9070),
            .I(N__9039));
    InMux I__2008 (
            .O(N__9069),
            .I(N__9036));
    InMux I__2007 (
            .O(N__9068),
            .I(N__9032));
    Span4Mux_v I__2006 (
            .O(N__9065),
            .I(N__9023));
    LocalMux I__2005 (
            .O(N__9062),
            .I(N__9023));
    LocalMux I__2004 (
            .O(N__9059),
            .I(N__9023));
    LocalMux I__2003 (
            .O(N__9052),
            .I(N__9023));
    InMux I__2002 (
            .O(N__9051),
            .I(N__9016));
    InMux I__2001 (
            .O(N__9050),
            .I(N__9016));
    LocalMux I__2000 (
            .O(N__9047),
            .I(N__9011));
    LocalMux I__1999 (
            .O(N__9044),
            .I(N__9011));
    LocalMux I__1998 (
            .O(N__9039),
            .I(N__9006));
    LocalMux I__1997 (
            .O(N__9036),
            .I(N__9006));
    InMux I__1996 (
            .O(N__9035),
            .I(N__8998));
    LocalMux I__1995 (
            .O(N__9032),
            .I(N__8991));
    Span4Mux_h I__1994 (
            .O(N__9023),
            .I(N__8991));
    InMux I__1993 (
            .O(N__9022),
            .I(N__8988));
    InMux I__1992 (
            .O(N__9021),
            .I(N__8985));
    LocalMux I__1991 (
            .O(N__9016),
            .I(N__8982));
    Span4Mux_v I__1990 (
            .O(N__9011),
            .I(N__8977));
    Span4Mux_v I__1989 (
            .O(N__9006),
            .I(N__8977));
    InMux I__1988 (
            .O(N__9005),
            .I(N__8970));
    InMux I__1987 (
            .O(N__9004),
            .I(N__8970));
    InMux I__1986 (
            .O(N__9003),
            .I(N__8970));
    InMux I__1985 (
            .O(N__9002),
            .I(N__8967));
    InMux I__1984 (
            .O(N__9001),
            .I(N__8964));
    LocalMux I__1983 (
            .O(N__8998),
            .I(N__8961));
    InMux I__1982 (
            .O(N__8997),
            .I(N__8956));
    InMux I__1981 (
            .O(N__8996),
            .I(N__8956));
    Span4Mux_h I__1980 (
            .O(N__8991),
            .I(N__8951));
    LocalMux I__1979 (
            .O(N__8988),
            .I(N__8951));
    LocalMux I__1978 (
            .O(N__8985),
            .I(N__8942));
    Span12Mux_s11_v I__1977 (
            .O(N__8982),
            .I(N__8942));
    Sp12to4 I__1976 (
            .O(N__8977),
            .I(N__8942));
    LocalMux I__1975 (
            .O(N__8970),
            .I(N__8942));
    LocalMux I__1974 (
            .O(N__8967),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1973 (
            .O(N__8964),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1972 (
            .O(N__8961),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1971 (
            .O(N__8956),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1970 (
            .O(N__8951),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__1969 (
            .O(N__8942),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    InMux I__1968 (
            .O(N__8929),
            .I(N__8923));
    InMux I__1967 (
            .O(N__8928),
            .I(N__8916));
    InMux I__1966 (
            .O(N__8927),
            .I(N__8916));
    InMux I__1965 (
            .O(N__8926),
            .I(N__8913));
    LocalMux I__1964 (
            .O(N__8923),
            .I(N__8910));
    InMux I__1963 (
            .O(N__8922),
            .I(N__8905));
    InMux I__1962 (
            .O(N__8921),
            .I(N__8905));
    LocalMux I__1961 (
            .O(N__8916),
            .I(N__8902));
    LocalMux I__1960 (
            .O(N__8913),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    Odrv4 I__1959 (
            .O(N__8910),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    LocalMux I__1958 (
            .O(N__8905),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    Odrv4 I__1957 (
            .O(N__8902),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    CascadeMux I__1956 (
            .O(N__8893),
            .I(N__8885));
    CascadeMux I__1955 (
            .O(N__8892),
            .I(N__8882));
    CascadeMux I__1954 (
            .O(N__8891),
            .I(N__8879));
    CascadeMux I__1953 (
            .O(N__8890),
            .I(N__8876));
    InMux I__1952 (
            .O(N__8889),
            .I(N__8871));
    InMux I__1951 (
            .O(N__8888),
            .I(N__8868));
    InMux I__1950 (
            .O(N__8885),
            .I(N__8864));
    InMux I__1949 (
            .O(N__8882),
            .I(N__8861));
    InMux I__1948 (
            .O(N__8879),
            .I(N__8856));
    InMux I__1947 (
            .O(N__8876),
            .I(N__8856));
    InMux I__1946 (
            .O(N__8875),
            .I(N__8851));
    InMux I__1945 (
            .O(N__8874),
            .I(N__8851));
    LocalMux I__1944 (
            .O(N__8871),
            .I(N__8848));
    LocalMux I__1943 (
            .O(N__8868),
            .I(N__8845));
    InMux I__1942 (
            .O(N__8867),
            .I(N__8842));
    LocalMux I__1941 (
            .O(N__8864),
            .I(\U712_CHIP_RAM.N_412 ));
    LocalMux I__1940 (
            .O(N__8861),
            .I(\U712_CHIP_RAM.N_412 ));
    LocalMux I__1939 (
            .O(N__8856),
            .I(\U712_CHIP_RAM.N_412 ));
    LocalMux I__1938 (
            .O(N__8851),
            .I(\U712_CHIP_RAM.N_412 ));
    Odrv4 I__1937 (
            .O(N__8848),
            .I(\U712_CHIP_RAM.N_412 ));
    Odrv4 I__1936 (
            .O(N__8845),
            .I(\U712_CHIP_RAM.N_412 ));
    LocalMux I__1935 (
            .O(N__8842),
            .I(\U712_CHIP_RAM.N_412 ));
    CascadeMux I__1934 (
            .O(N__8827),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_ ));
    IoInMux I__1933 (
            .O(N__8824),
            .I(N__8821));
    LocalMux I__1932 (
            .O(N__8821),
            .I(N__8818));
    IoSpan4Mux I__1931 (
            .O(N__8818),
            .I(N__8815));
    Span4Mux_s3_h I__1930 (
            .O(N__8815),
            .I(N__8812));
    Sp12to4 I__1929 (
            .O(N__8812),
            .I(N__8809));
    Span12Mux_h I__1928 (
            .O(N__8809),
            .I(N__8806));
    Odrv12 I__1927 (
            .O(N__8806),
            .I(CMA_c_4));
    InMux I__1926 (
            .O(N__8803),
            .I(N__8800));
    LocalMux I__1925 (
            .O(N__8800),
            .I(N__8770));
    ClkMux I__1924 (
            .O(N__8799),
            .I(N__8680));
    ClkMux I__1923 (
            .O(N__8798),
            .I(N__8680));
    ClkMux I__1922 (
            .O(N__8797),
            .I(N__8680));
    ClkMux I__1921 (
            .O(N__8796),
            .I(N__8680));
    ClkMux I__1920 (
            .O(N__8795),
            .I(N__8680));
    ClkMux I__1919 (
            .O(N__8794),
            .I(N__8680));
    ClkMux I__1918 (
            .O(N__8793),
            .I(N__8680));
    ClkMux I__1917 (
            .O(N__8792),
            .I(N__8680));
    ClkMux I__1916 (
            .O(N__8791),
            .I(N__8680));
    ClkMux I__1915 (
            .O(N__8790),
            .I(N__8680));
    ClkMux I__1914 (
            .O(N__8789),
            .I(N__8680));
    ClkMux I__1913 (
            .O(N__8788),
            .I(N__8680));
    ClkMux I__1912 (
            .O(N__8787),
            .I(N__8680));
    ClkMux I__1911 (
            .O(N__8786),
            .I(N__8680));
    ClkMux I__1910 (
            .O(N__8785),
            .I(N__8680));
    ClkMux I__1909 (
            .O(N__8784),
            .I(N__8680));
    ClkMux I__1908 (
            .O(N__8783),
            .I(N__8680));
    ClkMux I__1907 (
            .O(N__8782),
            .I(N__8680));
    ClkMux I__1906 (
            .O(N__8781),
            .I(N__8680));
    ClkMux I__1905 (
            .O(N__8780),
            .I(N__8680));
    ClkMux I__1904 (
            .O(N__8779),
            .I(N__8680));
    ClkMux I__1903 (
            .O(N__8778),
            .I(N__8680));
    ClkMux I__1902 (
            .O(N__8777),
            .I(N__8680));
    ClkMux I__1901 (
            .O(N__8776),
            .I(N__8680));
    ClkMux I__1900 (
            .O(N__8775),
            .I(N__8680));
    ClkMux I__1899 (
            .O(N__8774),
            .I(N__8680));
    ClkMux I__1898 (
            .O(N__8773),
            .I(N__8680));
    Glb2LocalMux I__1897 (
            .O(N__8770),
            .I(N__8680));
    ClkMux I__1896 (
            .O(N__8769),
            .I(N__8680));
    ClkMux I__1895 (
            .O(N__8768),
            .I(N__8680));
    ClkMux I__1894 (
            .O(N__8767),
            .I(N__8680));
    ClkMux I__1893 (
            .O(N__8766),
            .I(N__8680));
    ClkMux I__1892 (
            .O(N__8765),
            .I(N__8680));
    ClkMux I__1891 (
            .O(N__8764),
            .I(N__8680));
    ClkMux I__1890 (
            .O(N__8763),
            .I(N__8680));
    ClkMux I__1889 (
            .O(N__8762),
            .I(N__8680));
    ClkMux I__1888 (
            .O(N__8761),
            .I(N__8680));
    ClkMux I__1887 (
            .O(N__8760),
            .I(N__8680));
    ClkMux I__1886 (
            .O(N__8759),
            .I(N__8680));
    GlobalMux I__1885 (
            .O(N__8680),
            .I(CLK80_PLL));
    CEMux I__1884 (
            .O(N__8677),
            .I(N__8671));
    CEMux I__1883 (
            .O(N__8676),
            .I(N__8668));
    CEMux I__1882 (
            .O(N__8675),
            .I(N__8664));
    CEMux I__1881 (
            .O(N__8674),
            .I(N__8660));
    LocalMux I__1880 (
            .O(N__8671),
            .I(N__8655));
    LocalMux I__1879 (
            .O(N__8668),
            .I(N__8655));
    CEMux I__1878 (
            .O(N__8667),
            .I(N__8652));
    LocalMux I__1877 (
            .O(N__8664),
            .I(N__8649));
    CEMux I__1876 (
            .O(N__8663),
            .I(N__8646));
    LocalMux I__1875 (
            .O(N__8660),
            .I(N__8643));
    Span4Mux_v I__1874 (
            .O(N__8655),
            .I(N__8638));
    LocalMux I__1873 (
            .O(N__8652),
            .I(N__8638));
    Span4Mux_h I__1872 (
            .O(N__8649),
            .I(N__8633));
    LocalMux I__1871 (
            .O(N__8646),
            .I(N__8633));
    Span4Mux_h I__1870 (
            .O(N__8643),
            .I(N__8630));
    Span4Mux_v I__1869 (
            .O(N__8638),
            .I(N__8627));
    Span4Mux_h I__1868 (
            .O(N__8633),
            .I(N__8624));
    Odrv4 I__1867 (
            .O(N__8630),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__1866 (
            .O(N__8627),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    Odrv4 I__1865 (
            .O(N__8624),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__1864 (
            .O(N__8617),
            .I(N__8614));
    LocalMux I__1863 (
            .O(N__8614),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__1862 (
            .O(N__8611),
            .I(N__8608));
    LocalMux I__1861 (
            .O(N__8608),
            .I(N__8605));
    IoSpan4Mux I__1860 (
            .O(N__8605),
            .I(N__8602));
    Span4Mux_s2_h I__1859 (
            .O(N__8602),
            .I(N__8599));
    Sp12to4 I__1858 (
            .O(N__8599),
            .I(N__8596));
    Span12Mux_h I__1857 (
            .O(N__8596),
            .I(N__8593));
    Odrv12 I__1856 (
            .O(N__8593),
            .I(CMA_c_6));
    InMux I__1855 (
            .O(N__8590),
            .I(N__8587));
    LocalMux I__1854 (
            .O(N__8587),
            .I(N__8584));
    Span4Mux_v I__1853 (
            .O(N__8584),
            .I(N__8581));
    Span4Mux_v I__1852 (
            .O(N__8581),
            .I(N__8578));
    Sp12to4 I__1851 (
            .O(N__8578),
            .I(N__8575));
    Span12Mux_h I__1850 (
            .O(N__8575),
            .I(N__8572));
    Odrv12 I__1849 (
            .O(N__8572),
            .I(A_c_17));
    IoInMux I__1848 (
            .O(N__8569),
            .I(N__8566));
    LocalMux I__1847 (
            .O(N__8566),
            .I(N__8563));
    Span4Mux_s3_h I__1846 (
            .O(N__8563),
            .I(N__8560));
    Sp12to4 I__1845 (
            .O(N__8560),
            .I(N__8557));
    Span12Mux_s9_v I__1844 (
            .O(N__8557),
            .I(N__8554));
    Span12Mux_h I__1843 (
            .O(N__8554),
            .I(N__8551));
    Odrv12 I__1842 (
            .O(N__8551),
            .I(CMA_c_8));
    InMux I__1841 (
            .O(N__8548),
            .I(N__8545));
    LocalMux I__1840 (
            .O(N__8545),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1839 (
            .O(N__8542),
            .I(N__8539));
    LocalMux I__1838 (
            .O(N__8539),
            .I(N__8536));
    Span12Mux_s3_h I__1837 (
            .O(N__8536),
            .I(N__8533));
    Span12Mux_h I__1836 (
            .O(N__8533),
            .I(N__8530));
    Odrv12 I__1835 (
            .O(N__8530),
            .I(CMA_c_7));
    InMux I__1834 (
            .O(N__8527),
            .I(N__8524));
    LocalMux I__1833 (
            .O(N__8524),
            .I(N__8520));
    InMux I__1832 (
            .O(N__8523),
            .I(N__8517));
    Odrv4 I__1831 (
            .O(N__8520),
            .I(\U712_CHIP_RAM.CMA_5_i_0_8 ));
    LocalMux I__1830 (
            .O(N__8517),
            .I(\U712_CHIP_RAM.CMA_5_i_0_8 ));
    InMux I__1829 (
            .O(N__8512),
            .I(N__8509));
    LocalMux I__1828 (
            .O(N__8509),
            .I(N__8506));
    Span4Mux_v I__1827 (
            .O(N__8506),
            .I(N__8503));
    Span4Mux_v I__1826 (
            .O(N__8503),
            .I(N__8500));
    Sp12to4 I__1825 (
            .O(N__8500),
            .I(N__8497));
    Span12Mux_h I__1824 (
            .O(N__8497),
            .I(N__8494));
    Odrv12 I__1823 (
            .O(N__8494),
            .I(A_c_19));
    IoInMux I__1822 (
            .O(N__8491),
            .I(N__8488));
    LocalMux I__1821 (
            .O(N__8488),
            .I(N__8485));
    Span4Mux_s3_h I__1820 (
            .O(N__8485),
            .I(N__8482));
    Sp12to4 I__1819 (
            .O(N__8482),
            .I(N__8479));
    Span12Mux_s11_v I__1818 (
            .O(N__8479),
            .I(N__8476));
    Odrv12 I__1817 (
            .O(N__8476),
            .I(CMA_c_9));
    InMux I__1816 (
            .O(N__8473),
            .I(N__8470));
    LocalMux I__1815 (
            .O(N__8470),
            .I(N__8467));
    Odrv4 I__1814 (
            .O(N__8467),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__1813 (
            .O(N__8464),
            .I(N__8461));
    LocalMux I__1812 (
            .O(N__8461),
            .I(N__8458));
    Span4Mux_s2_h I__1811 (
            .O(N__8458),
            .I(N__8455));
    Span4Mux_v I__1810 (
            .O(N__8455),
            .I(N__8452));
    Sp12to4 I__1809 (
            .O(N__8452),
            .I(N__8449));
    Span12Mux_h I__1808 (
            .O(N__8449),
            .I(N__8446));
    Odrv12 I__1807 (
            .O(N__8446),
            .I(CMA_c_3));
    InMux I__1806 (
            .O(N__8443),
            .I(N__8440));
    LocalMux I__1805 (
            .O(N__8440),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__1804 (
            .O(N__8437),
            .I(N__8434));
    LocalMux I__1803 (
            .O(N__8434),
            .I(N__8431));
    Odrv4 I__1802 (
            .O(N__8431),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__1801 (
            .O(N__8428),
            .I(N__8425));
    LocalMux I__1800 (
            .O(N__8425),
            .I(N__8422));
    Odrv4 I__1799 (
            .O(N__8422),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    CascadeMux I__1798 (
            .O(N__8419),
            .I(N__8416));
    InMux I__1797 (
            .O(N__8416),
            .I(N__8413));
    LocalMux I__1796 (
            .O(N__8413),
            .I(N__8410));
    Odrv4 I__1795 (
            .O(N__8410),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    CascadeMux I__1794 (
            .O(N__8407),
            .I(\U712_BYTE_ENABLE.N_563_cascade_ ));
    IoInMux I__1793 (
            .O(N__8404),
            .I(N__8401));
    LocalMux I__1792 (
            .O(N__8401),
            .I(N__8398));
    Span4Mux_s2_v I__1791 (
            .O(N__8398),
            .I(N__8395));
    Span4Mux_h I__1790 (
            .O(N__8395),
            .I(N__8392));
    Sp12to4 I__1789 (
            .O(N__8392),
            .I(N__8389));
    Span12Mux_s10_v I__1788 (
            .O(N__8389),
            .I(N__8386));
    Odrv12 I__1787 (
            .O(N__8386),
            .I(N_56_i));
    IoInMux I__1786 (
            .O(N__8383),
            .I(N__8380));
    LocalMux I__1785 (
            .O(N__8380),
            .I(N__8377));
    IoSpan4Mux I__1784 (
            .O(N__8377),
            .I(N__8374));
    Sp12to4 I__1783 (
            .O(N__8374),
            .I(N__8371));
    Span12Mux_s7_v I__1782 (
            .O(N__8371),
            .I(N__8368));
    Odrv12 I__1781 (
            .O(N__8368),
            .I(WEn_c));
    InMux I__1780 (
            .O(N__8365),
            .I(N__8361));
    InMux I__1779 (
            .O(N__8364),
            .I(N__8358));
    LocalMux I__1778 (
            .O(N__8361),
            .I(N__8355));
    LocalMux I__1777 (
            .O(N__8358),
            .I(N__8347));
    Span4Mux_h I__1776 (
            .O(N__8355),
            .I(N__8347));
    InMux I__1775 (
            .O(N__8354),
            .I(N__8344));
    InMux I__1774 (
            .O(N__8353),
            .I(N__8341));
    CascadeMux I__1773 (
            .O(N__8352),
            .I(N__8338));
    Span4Mux_v I__1772 (
            .O(N__8347),
            .I(N__8331));
    LocalMux I__1771 (
            .O(N__8344),
            .I(N__8331));
    LocalMux I__1770 (
            .O(N__8341),
            .I(N__8331));
    InMux I__1769 (
            .O(N__8338),
            .I(N__8328));
    Span4Mux_h I__1768 (
            .O(N__8331),
            .I(N__8325));
    LocalMux I__1767 (
            .O(N__8328),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__1766 (
            .O(N__8325),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1765 (
            .O(N__8320),
            .I(N__8317));
    LocalMux I__1764 (
            .O(N__8317),
            .I(N__8314));
    Span4Mux_s3_v I__1763 (
            .O(N__8314),
            .I(N__8311));
    Span4Mux_v I__1762 (
            .O(N__8311),
            .I(N__8308));
    Span4Mux_h I__1761 (
            .O(N__8308),
            .I(N__8305));
    Odrv4 I__1760 (
            .O(N__8305),
            .I(CRCSn_c));
    InMux I__1759 (
            .O(N__8302),
            .I(N__8299));
    LocalMux I__1758 (
            .O(N__8299),
            .I(N__8292));
    InMux I__1757 (
            .O(N__8298),
            .I(N__8289));
    InMux I__1756 (
            .O(N__8297),
            .I(N__8286));
    CascadeMux I__1755 (
            .O(N__8296),
            .I(N__8283));
    CascadeMux I__1754 (
            .O(N__8295),
            .I(N__8280));
    Span4Mux_h I__1753 (
            .O(N__8292),
            .I(N__8277));
    LocalMux I__1752 (
            .O(N__8289),
            .I(N__8274));
    LocalMux I__1751 (
            .O(N__8286),
            .I(N__8271));
    InMux I__1750 (
            .O(N__8283),
            .I(N__8268));
    InMux I__1749 (
            .O(N__8280),
            .I(N__8265));
    Span4Mux_v I__1748 (
            .O(N__8277),
            .I(N__8262));
    Span4Mux_v I__1747 (
            .O(N__8274),
            .I(N__8259));
    Span4Mux_h I__1746 (
            .O(N__8271),
            .I(N__8254));
    LocalMux I__1745 (
            .O(N__8268),
            .I(N__8254));
    LocalMux I__1744 (
            .O(N__8265),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1743 (
            .O(N__8262),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1742 (
            .O(N__8259),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1741 (
            .O(N__8254),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    InMux I__1740 (
            .O(N__8245),
            .I(N__8242));
    LocalMux I__1739 (
            .O(N__8242),
            .I(N__8239));
    Odrv12 I__1738 (
            .O(N__8239),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__1737 (
            .O(N__8236),
            .I(N__8233));
    LocalMux I__1736 (
            .O(N__8233),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ));
    InMux I__1735 (
            .O(N__8230),
            .I(N__8227));
    LocalMux I__1734 (
            .O(N__8227),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__1733 (
            .O(N__8224),
            .I(N__8221));
    LocalMux I__1732 (
            .O(N__8221),
            .I(N__8218));
    Odrv12 I__1731 (
            .O(N__8218),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    IoInMux I__1730 (
            .O(N__8215),
            .I(N__8212));
    LocalMux I__1729 (
            .O(N__8212),
            .I(N__8209));
    IoSpan4Mux I__1728 (
            .O(N__8209),
            .I(N__8206));
    Span4Mux_s2_h I__1727 (
            .O(N__8206),
            .I(N__8203));
    Sp12to4 I__1726 (
            .O(N__8203),
            .I(N__8200));
    Span12Mux_h I__1725 (
            .O(N__8200),
            .I(N__8197));
    Odrv12 I__1724 (
            .O(N__8197),
            .I(CMA_c_5));
    CascadeMux I__1723 (
            .O(N__8194),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ));
    InMux I__1722 (
            .O(N__8191),
            .I(N__8188));
    LocalMux I__1721 (
            .O(N__8188),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    InMux I__1720 (
            .O(N__8185),
            .I(N__8179));
    InMux I__1719 (
            .O(N__8184),
            .I(N__8176));
    InMux I__1718 (
            .O(N__8183),
            .I(N__8173));
    InMux I__1717 (
            .O(N__8182),
            .I(N__8170));
    LocalMux I__1716 (
            .O(N__8179),
            .I(N__8163));
    LocalMux I__1715 (
            .O(N__8176),
            .I(N__8163));
    LocalMux I__1714 (
            .O(N__8173),
            .I(N__8163));
    LocalMux I__1713 (
            .O(N__8170),
            .I(N__8158));
    Span4Mux_h I__1712 (
            .O(N__8163),
            .I(N__8158));
    Sp12to4 I__1711 (
            .O(N__8158),
            .I(N__8155));
    Span12Mux_v I__1710 (
            .O(N__8155),
            .I(N__8152));
    Odrv12 I__1709 (
            .O(N__8152),
            .I(CLK40_PLL_i));
    IoInMux I__1708 (
            .O(N__8149),
            .I(N__8145));
    IoInMux I__1707 (
            .O(N__8148),
            .I(N__8142));
    LocalMux I__1706 (
            .O(N__8145),
            .I(N__8138));
    LocalMux I__1705 (
            .O(N__8142),
            .I(N__8135));
    IoInMux I__1704 (
            .O(N__8141),
            .I(N__8132));
    Span4Mux_s2_v I__1703 (
            .O(N__8138),
            .I(N__8129));
    Span4Mux_s2_v I__1702 (
            .O(N__8135),
            .I(N__8126));
    LocalMux I__1701 (
            .O(N__8132),
            .I(N__8123));
    Span4Mux_v I__1700 (
            .O(N__8129),
            .I(N__8120));
    Span4Mux_v I__1699 (
            .O(N__8126),
            .I(N__8117));
    Span4Mux_s3_h I__1698 (
            .O(N__8123),
            .I(N__8114));
    Sp12to4 I__1697 (
            .O(N__8120),
            .I(N__8109));
    Sp12to4 I__1696 (
            .O(N__8117),
            .I(N__8109));
    Span4Mux_h I__1695 (
            .O(N__8114),
            .I(N__8106));
    Span12Mux_s8_h I__1694 (
            .O(N__8109),
            .I(N__8103));
    Span4Mux_h I__1693 (
            .O(N__8106),
            .I(N__8100));
    Span12Mux_v I__1692 (
            .O(N__8103),
            .I(N__8097));
    Span4Mux_h I__1691 (
            .O(N__8100),
            .I(N__8094));
    Odrv12 I__1690 (
            .O(N__8097),
            .I(CLK40_PLL_i_i));
    Odrv4 I__1689 (
            .O(N__8094),
            .I(CLK40_PLL_i_i));
    InMux I__1688 (
            .O(N__8089),
            .I(N__8085));
    InMux I__1687 (
            .O(N__8088),
            .I(N__8082));
    LocalMux I__1686 (
            .O(N__8085),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__1685 (
            .O(N__8082),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__1684 (
            .O(N__8077),
            .I(N__8074));
    LocalMux I__1683 (
            .O(N__8074),
            .I(\U712_CYCLE_TERM.N_598 ));
    CascadeMux I__1682 (
            .O(N__8071),
            .I(N__8066));
    InMux I__1681 (
            .O(N__8070),
            .I(N__8063));
    InMux I__1680 (
            .O(N__8069),
            .I(N__8060));
    InMux I__1679 (
            .O(N__8066),
            .I(N__8057));
    LocalMux I__1678 (
            .O(N__8063),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    LocalMux I__1677 (
            .O(N__8060),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    LocalMux I__1676 (
            .O(N__8057),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    InMux I__1675 (
            .O(N__8050),
            .I(N__8046));
    InMux I__1674 (
            .O(N__8049),
            .I(N__8043));
    LocalMux I__1673 (
            .O(N__8046),
            .I(\U712_CYCLE_TERM.N_440 ));
    LocalMux I__1672 (
            .O(N__8043),
            .I(\U712_CYCLE_TERM.N_440 ));
    InMux I__1671 (
            .O(N__8038),
            .I(N__8035));
    LocalMux I__1670 (
            .O(N__8035),
            .I(\U712_CYCLE_TERM.un13_0 ));
    InMux I__1669 (
            .O(N__8032),
            .I(N__8015));
    InMux I__1668 (
            .O(N__8031),
            .I(N__8015));
    InMux I__1667 (
            .O(N__8030),
            .I(N__8015));
    InMux I__1666 (
            .O(N__8029),
            .I(N__8008));
    InMux I__1665 (
            .O(N__8028),
            .I(N__8008));
    InMux I__1664 (
            .O(N__8027),
            .I(N__8008));
    InMux I__1663 (
            .O(N__8026),
            .I(N__8004));
    InMux I__1662 (
            .O(N__8025),
            .I(N__8001));
    InMux I__1661 (
            .O(N__8024),
            .I(N__7996));
    InMux I__1660 (
            .O(N__8023),
            .I(N__7991));
    InMux I__1659 (
            .O(N__8022),
            .I(N__7991));
    LocalMux I__1658 (
            .O(N__8015),
            .I(N__7979));
    LocalMux I__1657 (
            .O(N__8008),
            .I(N__7979));
    InMux I__1656 (
            .O(N__8007),
            .I(N__7976));
    LocalMux I__1655 (
            .O(N__8004),
            .I(N__7972));
    LocalMux I__1654 (
            .O(N__8001),
            .I(N__7969));
    InMux I__1653 (
            .O(N__8000),
            .I(N__7964));
    InMux I__1652 (
            .O(N__7999),
            .I(N__7964));
    LocalMux I__1651 (
            .O(N__7996),
            .I(N__7954));
    LocalMux I__1650 (
            .O(N__7991),
            .I(N__7954));
    InMux I__1649 (
            .O(N__7990),
            .I(N__7951));
    InMux I__1648 (
            .O(N__7989),
            .I(N__7944));
    InMux I__1647 (
            .O(N__7988),
            .I(N__7944));
    InMux I__1646 (
            .O(N__7987),
            .I(N__7941));
    InMux I__1645 (
            .O(N__7986),
            .I(N__7938));
    InMux I__1644 (
            .O(N__7985),
            .I(N__7933));
    InMux I__1643 (
            .O(N__7984),
            .I(N__7933));
    Span4Mux_v I__1642 (
            .O(N__7979),
            .I(N__7928));
    LocalMux I__1641 (
            .O(N__7976),
            .I(N__7928));
    InMux I__1640 (
            .O(N__7975),
            .I(N__7925));
    Span4Mux_v I__1639 (
            .O(N__7972),
            .I(N__7917));
    Span4Mux_v I__1638 (
            .O(N__7969),
            .I(N__7917));
    LocalMux I__1637 (
            .O(N__7964),
            .I(N__7917));
    InMux I__1636 (
            .O(N__7963),
            .I(N__7908));
    InMux I__1635 (
            .O(N__7962),
            .I(N__7908));
    InMux I__1634 (
            .O(N__7961),
            .I(N__7908));
    InMux I__1633 (
            .O(N__7960),
            .I(N__7908));
    InMux I__1632 (
            .O(N__7959),
            .I(N__7905));
    Span4Mux_v I__1631 (
            .O(N__7954),
            .I(N__7900));
    LocalMux I__1630 (
            .O(N__7951),
            .I(N__7900));
    InMux I__1629 (
            .O(N__7950),
            .I(N__7897));
    InMux I__1628 (
            .O(N__7949),
            .I(N__7894));
    LocalMux I__1627 (
            .O(N__7944),
            .I(N__7885));
    LocalMux I__1626 (
            .O(N__7941),
            .I(N__7885));
    LocalMux I__1625 (
            .O(N__7938),
            .I(N__7885));
    LocalMux I__1624 (
            .O(N__7933),
            .I(N__7885));
    Span4Mux_v I__1623 (
            .O(N__7928),
            .I(N__7880));
    LocalMux I__1622 (
            .O(N__7925),
            .I(N__7880));
    InMux I__1621 (
            .O(N__7924),
            .I(N__7877));
    Span4Mux_h I__1620 (
            .O(N__7917),
            .I(N__7872));
    LocalMux I__1619 (
            .O(N__7908),
            .I(N__7872));
    LocalMux I__1618 (
            .O(N__7905),
            .I(N__7865));
    Span4Mux_v I__1617 (
            .O(N__7900),
            .I(N__7865));
    LocalMux I__1616 (
            .O(N__7897),
            .I(N__7865));
    LocalMux I__1615 (
            .O(N__7894),
            .I(N__7862));
    Span4Mux_v I__1614 (
            .O(N__7885),
            .I(N__7857));
    Span4Mux_v I__1613 (
            .O(N__7880),
            .I(N__7857));
    LocalMux I__1612 (
            .O(N__7877),
            .I(N__7854));
    Span4Mux_v I__1611 (
            .O(N__7872),
            .I(N__7847));
    Span4Mux_v I__1610 (
            .O(N__7865),
            .I(N__7847));
    Span4Mux_v I__1609 (
            .O(N__7862),
            .I(N__7847));
    Sp12to4 I__1608 (
            .O(N__7857),
            .I(N__7844));
    Span12Mux_v I__1607 (
            .O(N__7854),
            .I(N__7839));
    Sp12to4 I__1606 (
            .O(N__7847),
            .I(N__7839));
    Span12Mux_h I__1605 (
            .O(N__7844),
            .I(N__7836));
    Span12Mux_h I__1604 (
            .O(N__7839),
            .I(N__7833));
    Odrv12 I__1603 (
            .O(N__7836),
            .I(RESETn_c));
    Odrv12 I__1602 (
            .O(N__7833),
            .I(RESETn_c));
    InMux I__1601 (
            .O(N__7828),
            .I(N__7825));
    LocalMux I__1600 (
            .O(N__7825),
            .I(\U712_CYCLE_TERM.N_566 ));
    CascadeMux I__1599 (
            .O(N__7822),
            .I(\U712_CYCLE_TERM.un13_0_cascade_ ));
    CascadeMux I__1598 (
            .O(N__7819),
            .I(N__7816));
    InMux I__1597 (
            .O(N__7816),
            .I(N__7813));
    LocalMux I__1596 (
            .O(N__7813),
            .I(N__7810));
    Odrv12 I__1595 (
            .O(N__7810),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    InMux I__1594 (
            .O(N__7807),
            .I(N__7804));
    LocalMux I__1593 (
            .O(N__7804),
            .I(N__7797));
    CascadeMux I__1592 (
            .O(N__7803),
            .I(N__7787));
    CascadeMux I__1591 (
            .O(N__7802),
            .I(N__7784));
    InMux I__1590 (
            .O(N__7801),
            .I(N__7779));
    InMux I__1589 (
            .O(N__7800),
            .I(N__7776));
    Span4Mux_h I__1588 (
            .O(N__7797),
            .I(N__7773));
    InMux I__1587 (
            .O(N__7796),
            .I(N__7768));
    InMux I__1586 (
            .O(N__7795),
            .I(N__7768));
    InMux I__1585 (
            .O(N__7794),
            .I(N__7765));
    InMux I__1584 (
            .O(N__7793),
            .I(N__7760));
    InMux I__1583 (
            .O(N__7792),
            .I(N__7760));
    InMux I__1582 (
            .O(N__7791),
            .I(N__7753));
    InMux I__1581 (
            .O(N__7790),
            .I(N__7753));
    InMux I__1580 (
            .O(N__7787),
            .I(N__7753));
    InMux I__1579 (
            .O(N__7784),
            .I(N__7746));
    InMux I__1578 (
            .O(N__7783),
            .I(N__7746));
    InMux I__1577 (
            .O(N__7782),
            .I(N__7746));
    LocalMux I__1576 (
            .O(N__7779),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1575 (
            .O(N__7776),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1574 (
            .O(N__7773),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1573 (
            .O(N__7768),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1572 (
            .O(N__7765),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1571 (
            .O(N__7760),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1570 (
            .O(N__7753),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1569 (
            .O(N__7746),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1568 (
            .O(N__7729),
            .I(N__7726));
    LocalMux I__1567 (
            .O(N__7726),
            .I(N__7723));
    Span4Mux_h I__1566 (
            .O(N__7723),
            .I(N__7720));
    Odrv4 I__1565 (
            .O(N__7720),
            .I(\U712_CHIP_RAM.N_93 ));
    IoInMux I__1564 (
            .O(N__7717),
            .I(N__7714));
    LocalMux I__1563 (
            .O(N__7714),
            .I(N__7711));
    IoSpan4Mux I__1562 (
            .O(N__7711),
            .I(N__7707));
    InMux I__1561 (
            .O(N__7710),
            .I(N__7704));
    Span4Mux_s2_v I__1560 (
            .O(N__7707),
            .I(N__7701));
    LocalMux I__1559 (
            .O(N__7704),
            .I(N__7698));
    Sp12to4 I__1558 (
            .O(N__7701),
            .I(N__7695));
    Span4Mux_v I__1557 (
            .O(N__7698),
            .I(N__7692));
    Span12Mux_s8_v I__1556 (
            .O(N__7695),
            .I(N__7689));
    Sp12to4 I__1555 (
            .O(N__7692),
            .I(N__7686));
    Span12Mux_v I__1554 (
            .O(N__7689),
            .I(N__7681));
    Span12Mux_h I__1553 (
            .O(N__7686),
            .I(N__7681));
    Span12Mux_h I__1552 (
            .O(N__7681),
            .I(N__7678));
    Odrv12 I__1551 (
            .O(N__7678),
            .I(A_c_10));
    InMux I__1550 (
            .O(N__7675),
            .I(N__7672));
    LocalMux I__1549 (
            .O(N__7672),
            .I(N__7669));
    Odrv12 I__1548 (
            .O(N__7669),
            .I(\U712_CHIP_RAM.N_455 ));
    IoInMux I__1547 (
            .O(N__7666),
            .I(N__7662));
    InMux I__1546 (
            .O(N__7665),
            .I(N__7659));
    LocalMux I__1545 (
            .O(N__7662),
            .I(N__7656));
    LocalMux I__1544 (
            .O(N__7659),
            .I(N__7653));
    Span12Mux_s9_h I__1543 (
            .O(N__7656),
            .I(N__7649));
    Span4Mux_v I__1542 (
            .O(N__7653),
            .I(N__7646));
    InMux I__1541 (
            .O(N__7652),
            .I(N__7643));
    Span12Mux_v I__1540 (
            .O(N__7649),
            .I(N__7639));
    Span4Mux_h I__1539 (
            .O(N__7646),
            .I(N__7636));
    LocalMux I__1538 (
            .O(N__7643),
            .I(N__7633));
    InMux I__1537 (
            .O(N__7642),
            .I(N__7630));
    Odrv12 I__1536 (
            .O(N__7639),
            .I(TACK_OUTn));
    Odrv4 I__1535 (
            .O(N__7636),
            .I(TACK_OUTn));
    Odrv4 I__1534 (
            .O(N__7633),
            .I(TACK_OUTn));
    LocalMux I__1533 (
            .O(N__7630),
            .I(TACK_OUTn));
    InMux I__1532 (
            .O(N__7621),
            .I(N__7617));
    InMux I__1531 (
            .O(N__7620),
            .I(N__7614));
    LocalMux I__1530 (
            .O(N__7617),
            .I(\U712_CYCLE_TERM.RAM_CYCLEZ0 ));
    LocalMux I__1529 (
            .O(N__7614),
            .I(\U712_CYCLE_TERM.RAM_CYCLEZ0 ));
    IoInMux I__1528 (
            .O(N__7609),
            .I(N__7606));
    LocalMux I__1527 (
            .O(N__7606),
            .I(N__7603));
    Span4Mux_s3_h I__1526 (
            .O(N__7603),
            .I(N__7600));
    Span4Mux_h I__1525 (
            .O(N__7600),
            .I(N__7596));
    InMux I__1524 (
            .O(N__7599),
            .I(N__7593));
    Sp12to4 I__1523 (
            .O(N__7596),
            .I(N__7590));
    LocalMux I__1522 (
            .O(N__7593),
            .I(N__7587));
    Span12Mux_v I__1521 (
            .O(N__7590),
            .I(N__7580));
    Span12Mux_s7_h I__1520 (
            .O(N__7587),
            .I(N__7580));
    InMux I__1519 (
            .O(N__7586),
            .I(N__7577));
    InMux I__1518 (
            .O(N__7585),
            .I(N__7574));
    Odrv12 I__1517 (
            .O(N__7580),
            .I(TACK_EN));
    LocalMux I__1516 (
            .O(N__7577),
            .I(TACK_EN));
    LocalMux I__1515 (
            .O(N__7574),
            .I(TACK_EN));
    IoInMux I__1514 (
            .O(N__7567),
            .I(N__7564));
    LocalMux I__1513 (
            .O(N__7564),
            .I(N__7561));
    Span4Mux_s2_v I__1512 (
            .O(N__7561),
            .I(N__7558));
    Sp12to4 I__1511 (
            .O(N__7558),
            .I(N__7555));
    Span12Mux_s11_h I__1510 (
            .O(N__7555),
            .I(N__7552));
    Span12Mux_v I__1509 (
            .O(N__7552),
            .I(N__7549));
    Odrv12 I__1508 (
            .O(N__7549),
            .I(U712_CYCLE_TERM_TCIn_0_i));
    IoInMux I__1507 (
            .O(N__7546),
            .I(N__7543));
    LocalMux I__1506 (
            .O(N__7543),
            .I(N__7540));
    Span4Mux_s2_v I__1505 (
            .O(N__7540),
            .I(N__7537));
    Span4Mux_h I__1504 (
            .O(N__7537),
            .I(N__7534));
    Sp12to4 I__1503 (
            .O(N__7534),
            .I(N__7530));
    InMux I__1502 (
            .O(N__7533),
            .I(N__7527));
    Span12Mux_s9_v I__1501 (
            .O(N__7530),
            .I(N__7524));
    LocalMux I__1500 (
            .O(N__7527),
            .I(N__7521));
    Odrv12 I__1499 (
            .O(N__7524),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__1498 (
            .O(N__7521),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1497 (
            .O(N__7516),
            .I(\U712_CHIP_RAM.N_412_cascade_ ));
    InMux I__1496 (
            .O(N__7513),
            .I(N__7510));
    LocalMux I__1495 (
            .O(N__7510),
            .I(N__7507));
    Span4Mux_v I__1494 (
            .O(N__7507),
            .I(N__7504));
    Sp12to4 I__1493 (
            .O(N__7504),
            .I(N__7501));
    Span12Mux_h I__1492 (
            .O(N__7501),
            .I(N__7498));
    Span12Mux_v I__1491 (
            .O(N__7498),
            .I(N__7495));
    Odrv12 I__1490 (
            .O(N__7495),
            .I(A_c_3));
    InMux I__1489 (
            .O(N__7492),
            .I(N__7489));
    LocalMux I__1488 (
            .O(N__7489),
            .I(\U712_CHIP_RAM.N_478 ));
    InMux I__1487 (
            .O(N__7486),
            .I(N__7483));
    LocalMux I__1486 (
            .O(N__7483),
            .I(N__7480));
    Span4Mux_h I__1485 (
            .O(N__7480),
            .I(N__7477));
    Odrv4 I__1484 (
            .O(N__7477),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ));
    InMux I__1483 (
            .O(N__7474),
            .I(N__7471));
    LocalMux I__1482 (
            .O(N__7471),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ));
    CascadeMux I__1481 (
            .O(N__7468),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_ ));
    IoInMux I__1480 (
            .O(N__7465),
            .I(N__7462));
    LocalMux I__1479 (
            .O(N__7462),
            .I(N__7459));
    Span12Mux_s11_v I__1478 (
            .O(N__7459),
            .I(N__7456));
    Odrv12 I__1477 (
            .O(N__7456),
            .I(CMA_c_0));
    IoInMux I__1476 (
            .O(N__7453),
            .I(N__7450));
    LocalMux I__1475 (
            .O(N__7450),
            .I(N__7447));
    Span4Mux_s3_v I__1474 (
            .O(N__7447),
            .I(N__7444));
    Span4Mux_v I__1473 (
            .O(N__7444),
            .I(N__7441));
    Span4Mux_v I__1472 (
            .O(N__7441),
            .I(N__7438));
    Odrv4 I__1471 (
            .O(N__7438),
            .I(CMA_c_2));
    InMux I__1470 (
            .O(N__7435),
            .I(N__7432));
    LocalMux I__1469 (
            .O(N__7432),
            .I(N__7429));
    Span4Mux_v I__1468 (
            .O(N__7429),
            .I(N__7426));
    Span4Mux_v I__1467 (
            .O(N__7426),
            .I(N__7423));
    Sp12to4 I__1466 (
            .O(N__7423),
            .I(N__7420));
    Span12Mux_h I__1465 (
            .O(N__7420),
            .I(N__7417));
    Odrv12 I__1464 (
            .O(N__7417),
            .I(A_c_4));
    IoInMux I__1463 (
            .O(N__7414),
            .I(N__7411));
    LocalMux I__1462 (
            .O(N__7411),
            .I(N__7408));
    IoSpan4Mux I__1461 (
            .O(N__7408),
            .I(N__7405));
    Span4Mux_s2_v I__1460 (
            .O(N__7405),
            .I(N__7402));
    Sp12to4 I__1459 (
            .O(N__7402),
            .I(N__7398));
    InMux I__1458 (
            .O(N__7401),
            .I(N__7395));
    Span12Mux_s8_v I__1457 (
            .O(N__7398),
            .I(N__7392));
    LocalMux I__1456 (
            .O(N__7395),
            .I(N__7389));
    Span12Mux_v I__1455 (
            .O(N__7392),
            .I(N__7386));
    Span12Mux_v I__1454 (
            .O(N__7389),
            .I(N__7383));
    Span12Mux_h I__1453 (
            .O(N__7386),
            .I(N__7380));
    Span12Mux_h I__1452 (
            .O(N__7383),
            .I(N__7377));
    Odrv12 I__1451 (
            .O(N__7380),
            .I(A_c_11));
    Odrv12 I__1450 (
            .O(N__7377),
            .I(A_c_11));
    InMux I__1449 (
            .O(N__7372),
            .I(N__7367));
    InMux I__1448 (
            .O(N__7371),
            .I(N__7362));
    InMux I__1447 (
            .O(N__7370),
            .I(N__7362));
    LocalMux I__1446 (
            .O(N__7367),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__1445 (
            .O(N__7362),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    CascadeMux I__1444 (
            .O(N__7357),
            .I(N__7354));
    InMux I__1443 (
            .O(N__7354),
            .I(N__7351));
    LocalMux I__1442 (
            .O(N__7351),
            .I(N__7345));
    InMux I__1441 (
            .O(N__7350),
            .I(N__7338));
    InMux I__1440 (
            .O(N__7349),
            .I(N__7338));
    InMux I__1439 (
            .O(N__7348),
            .I(N__7338));
    Odrv4 I__1438 (
            .O(N__7345),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1437 (
            .O(N__7338),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__1436 (
            .O(N__7333),
            .I(N__7329));
    InMux I__1435 (
            .O(N__7332),
            .I(N__7326));
    LocalMux I__1434 (
            .O(N__7329),
            .I(\U712_REG_SM.N_407 ));
    LocalMux I__1433 (
            .O(N__7326),
            .I(\U712_REG_SM.N_407 ));
    CascadeMux I__1432 (
            .O(N__7321),
            .I(N__7317));
    InMux I__1431 (
            .O(N__7320),
            .I(N__7311));
    InMux I__1430 (
            .O(N__7317),
            .I(N__7308));
    InMux I__1429 (
            .O(N__7316),
            .I(N__7305));
    InMux I__1428 (
            .O(N__7315),
            .I(N__7302));
    InMux I__1427 (
            .O(N__7314),
            .I(N__7298));
    LocalMux I__1426 (
            .O(N__7311),
            .I(N__7295));
    LocalMux I__1425 (
            .O(N__7308),
            .I(N__7290));
    LocalMux I__1424 (
            .O(N__7305),
            .I(N__7290));
    LocalMux I__1423 (
            .O(N__7302),
            .I(N__7287));
    InMux I__1422 (
            .O(N__7301),
            .I(N__7284));
    LocalMux I__1421 (
            .O(N__7298),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv12 I__1420 (
            .O(N__7295),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv4 I__1419 (
            .O(N__7290),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv4 I__1418 (
            .O(N__7287),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1417 (
            .O(N__7284),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    CascadeMux I__1416 (
            .O(N__7273),
            .I(N__7269));
    InMux I__1415 (
            .O(N__7272),
            .I(N__7261));
    InMux I__1414 (
            .O(N__7269),
            .I(N__7256));
    InMux I__1413 (
            .O(N__7268),
            .I(N__7256));
    InMux I__1412 (
            .O(N__7267),
            .I(N__7247));
    InMux I__1411 (
            .O(N__7266),
            .I(N__7247));
    InMux I__1410 (
            .O(N__7265),
            .I(N__7247));
    InMux I__1409 (
            .O(N__7264),
            .I(N__7247));
    LocalMux I__1408 (
            .O(N__7261),
            .I(N__7240));
    LocalMux I__1407 (
            .O(N__7256),
            .I(N__7240));
    LocalMux I__1406 (
            .O(N__7247),
            .I(N__7240));
    Odrv4 I__1405 (
            .O(N__7240),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    InMux I__1404 (
            .O(N__7237),
            .I(N__7232));
    InMux I__1403 (
            .O(N__7236),
            .I(N__7229));
    CascadeMux I__1402 (
            .O(N__7235),
            .I(N__7225));
    LocalMux I__1401 (
            .O(N__7232),
            .I(N__7222));
    LocalMux I__1400 (
            .O(N__7229),
            .I(N__7219));
    InMux I__1399 (
            .O(N__7228),
            .I(N__7216));
    InMux I__1398 (
            .O(N__7225),
            .I(N__7213));
    Sp12to4 I__1397 (
            .O(N__7222),
            .I(N__7210));
    Sp12to4 I__1396 (
            .O(N__7219),
            .I(N__7205));
    LocalMux I__1395 (
            .O(N__7216),
            .I(N__7205));
    LocalMux I__1394 (
            .O(N__7213),
            .I(N__7202));
    Span12Mux_v I__1393 (
            .O(N__7210),
            .I(N__7199));
    Span12Mux_h I__1392 (
            .O(N__7205),
            .I(N__7196));
    Span12Mux_v I__1391 (
            .O(N__7202),
            .I(N__7193));
    Span12Mux_h I__1390 (
            .O(N__7199),
            .I(N__7188));
    Span12Mux_v I__1389 (
            .O(N__7196),
            .I(N__7188));
    Span12Mux_h I__1388 (
            .O(N__7193),
            .I(N__7185));
    Odrv12 I__1387 (
            .O(N__7188),
            .I(RnW_c));
    Odrv12 I__1386 (
            .O(N__7185),
            .I(RnW_c));
    InMux I__1385 (
            .O(N__7180),
            .I(N__7175));
    InMux I__1384 (
            .O(N__7179),
            .I(N__7172));
    InMux I__1383 (
            .O(N__7178),
            .I(N__7169));
    LocalMux I__1382 (
            .O(N__7175),
            .I(N__7162));
    LocalMux I__1381 (
            .O(N__7172),
            .I(N__7162));
    LocalMux I__1380 (
            .O(N__7169),
            .I(N__7157));
    InMux I__1379 (
            .O(N__7168),
            .I(N__7154));
    InMux I__1378 (
            .O(N__7167),
            .I(N__7151));
    Span4Mux_h I__1377 (
            .O(N__7162),
            .I(N__7148));
    InMux I__1376 (
            .O(N__7161),
            .I(N__7145));
    InMux I__1375 (
            .O(N__7160),
            .I(N__7140));
    Span4Mux_h I__1374 (
            .O(N__7157),
            .I(N__7133));
    LocalMux I__1373 (
            .O(N__7154),
            .I(N__7133));
    LocalMux I__1372 (
            .O(N__7151),
            .I(N__7133));
    Sp12to4 I__1371 (
            .O(N__7148),
            .I(N__7129));
    LocalMux I__1370 (
            .O(N__7145),
            .I(N__7126));
    InMux I__1369 (
            .O(N__7144),
            .I(N__7121));
    InMux I__1368 (
            .O(N__7143),
            .I(N__7121));
    LocalMux I__1367 (
            .O(N__7140),
            .I(N__7118));
    Span4Mux_v I__1366 (
            .O(N__7133),
            .I(N__7115));
    InMux I__1365 (
            .O(N__7132),
            .I(N__7112));
    Odrv12 I__1364 (
            .O(N__7129),
            .I(WRITE_CYCLEm));
    Odrv4 I__1363 (
            .O(N__7126),
            .I(WRITE_CYCLEm));
    LocalMux I__1362 (
            .O(N__7121),
            .I(WRITE_CYCLEm));
    Odrv4 I__1361 (
            .O(N__7118),
            .I(WRITE_CYCLEm));
    Odrv4 I__1360 (
            .O(N__7115),
            .I(WRITE_CYCLEm));
    LocalMux I__1359 (
            .O(N__7112),
            .I(WRITE_CYCLEm));
    IoInMux I__1358 (
            .O(N__7099),
            .I(N__7096));
    LocalMux I__1357 (
            .O(N__7096),
            .I(N__7093));
    Span4Mux_s1_h I__1356 (
            .O(N__7093),
            .I(N__7090));
    Span4Mux_h I__1355 (
            .O(N__7090),
            .I(N__7087));
    Sp12to4 I__1354 (
            .O(N__7087),
            .I(N__7084));
    Span12Mux_s10_v I__1353 (
            .O(N__7084),
            .I(N__7081));
    Span12Mux_h I__1352 (
            .O(N__7081),
            .I(N__7078));
    Odrv12 I__1351 (
            .O(N__7078),
            .I(N_483));
    IoInMux I__1350 (
            .O(N__7075),
            .I(N__7072));
    LocalMux I__1349 (
            .O(N__7072),
            .I(N__7069));
    Span12Mux_s8_v I__1348 (
            .O(N__7069),
            .I(N__7066));
    Odrv12 I__1347 (
            .O(N__7066),
            .I(CMA_c_10));
    IoInMux I__1346 (
            .O(N__7063),
            .I(N__7060));
    LocalMux I__1345 (
            .O(N__7060),
            .I(N__7057));
    Odrv12 I__1344 (
            .O(N__7057),
            .I(CMA_c_1));
    InMux I__1343 (
            .O(N__7054),
            .I(N__7051));
    LocalMux I__1342 (
            .O(N__7051),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i ));
    CascadeMux I__1341 (
            .O(N__7048),
            .I(\U712_CYCLE_TERM.TACK_EN_RNOZ0Z_0_cascade_ ));
    CascadeMux I__1340 (
            .O(N__7045),
            .I(\U712_CYCLE_TERM.N_598_cascade_ ));
    CascadeMux I__1339 (
            .O(N__7042),
            .I(N__7038));
    InMux I__1338 (
            .O(N__7041),
            .I(N__7034));
    InMux I__1337 (
            .O(N__7038),
            .I(N__7031));
    InMux I__1336 (
            .O(N__7037),
            .I(N__7028));
    LocalMux I__1335 (
            .O(N__7034),
            .I(N__7025));
    LocalMux I__1334 (
            .O(N__7031),
            .I(N__7022));
    LocalMux I__1333 (
            .O(N__7028),
            .I(\U712_REG_SM.N_422 ));
    Odrv4 I__1332 (
            .O(N__7025),
            .I(\U712_REG_SM.N_422 ));
    Odrv12 I__1331 (
            .O(N__7022),
            .I(\U712_REG_SM.N_422 ));
    InMux I__1330 (
            .O(N__7015),
            .I(N__7012));
    LocalMux I__1329 (
            .O(N__7012),
            .I(N__7009));
    Span4Mux_h I__1328 (
            .O(N__7009),
            .I(N__7006));
    Odrv4 I__1327 (
            .O(N__7006),
            .I(\U712_REG_SM.N_514 ));
    CascadeMux I__1326 (
            .O(N__7003),
            .I(N__6999));
    InMux I__1325 (
            .O(N__7002),
            .I(N__6994));
    InMux I__1324 (
            .O(N__6999),
            .I(N__6987));
    InMux I__1323 (
            .O(N__6998),
            .I(N__6987));
    InMux I__1322 (
            .O(N__6997),
            .I(N__6987));
    LocalMux I__1321 (
            .O(N__6994),
            .I(REG_TACK));
    LocalMux I__1320 (
            .O(N__6987),
            .I(REG_TACK));
    CascadeMux I__1319 (
            .O(N__6982),
            .I(N__6979));
    InMux I__1318 (
            .O(N__6979),
            .I(N__6973));
    InMux I__1317 (
            .O(N__6978),
            .I(N__6966));
    InMux I__1316 (
            .O(N__6977),
            .I(N__6966));
    InMux I__1315 (
            .O(N__6976),
            .I(N__6966));
    LocalMux I__1314 (
            .O(N__6973),
            .I(N__6963));
    LocalMux I__1313 (
            .O(N__6966),
            .I(N__6960));
    Span4Mux_h I__1312 (
            .O(N__6963),
            .I(N__6957));
    Span4Mux_h I__1311 (
            .O(N__6960),
            .I(N__6954));
    Odrv4 I__1310 (
            .O(N__6957),
            .I(CPU_TACKm));
    Odrv4 I__1309 (
            .O(N__6954),
            .I(CPU_TACKm));
    InMux I__1308 (
            .O(N__6949),
            .I(N__6941));
    InMux I__1307 (
            .O(N__6948),
            .I(N__6941));
    InMux I__1306 (
            .O(N__6947),
            .I(N__6936));
    InMux I__1305 (
            .O(N__6946),
            .I(N__6936));
    LocalMux I__1304 (
            .O(N__6941),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__1303 (
            .O(N__6936),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__1302 (
            .O(N__6931),
            .I(\U712_CYCLE_TERM.N_571_cascade_ ));
    InMux I__1301 (
            .O(N__6928),
            .I(N__6924));
    InMux I__1300 (
            .O(N__6927),
            .I(N__6921));
    LocalMux I__1299 (
            .O(N__6924),
            .I(\U712_REG_SM.N_480 ));
    LocalMux I__1298 (
            .O(N__6921),
            .I(\U712_REG_SM.N_480 ));
    InMux I__1297 (
            .O(N__6916),
            .I(N__6913));
    LocalMux I__1296 (
            .O(N__6913),
            .I(\U712_REG_SM.REG_TACK_RNOZ0Z_0 ));
    InMux I__1295 (
            .O(N__6910),
            .I(N__6906));
    InMux I__1294 (
            .O(N__6909),
            .I(N__6903));
    LocalMux I__1293 (
            .O(N__6906),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__1292 (
            .O(N__6903),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__1291 (
            .O(N__6898),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__1290 (
            .O(N__6895),
            .I(N__6891));
    InMux I__1289 (
            .O(N__6894),
            .I(N__6888));
    LocalMux I__1288 (
            .O(N__6891),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__1287 (
            .O(N__6888),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__1286 (
            .O(N__6883),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__1285 (
            .O(N__6880),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    InMux I__1284 (
            .O(N__6877),
            .I(N__6873));
    InMux I__1283 (
            .O(N__6876),
            .I(N__6870));
    LocalMux I__1282 (
            .O(N__6873),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__1281 (
            .O(N__6870),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    ClkMux I__1280 (
            .O(N__6865),
            .I(N__6841));
    ClkMux I__1279 (
            .O(N__6864),
            .I(N__6841));
    ClkMux I__1278 (
            .O(N__6863),
            .I(N__6841));
    ClkMux I__1277 (
            .O(N__6862),
            .I(N__6841));
    ClkMux I__1276 (
            .O(N__6861),
            .I(N__6841));
    ClkMux I__1275 (
            .O(N__6860),
            .I(N__6841));
    ClkMux I__1274 (
            .O(N__6859),
            .I(N__6841));
    ClkMux I__1273 (
            .O(N__6858),
            .I(N__6841));
    GlobalMux I__1272 (
            .O(N__6841),
            .I(N__6838));
    gio2CtrlBuf I__1271 (
            .O(N__6838),
            .I(C1_c_g));
    InMux I__1270 (
            .O(N__6835),
            .I(N__6832));
    LocalMux I__1269 (
            .O(N__6832),
            .I(N__6829));
    Span4Mux_v I__1268 (
            .O(N__6829),
            .I(N__6826));
    Sp12to4 I__1267 (
            .O(N__6826),
            .I(N__6823));
    Span12Mux_h I__1266 (
            .O(N__6823),
            .I(N__6820));
    Span12Mux_v I__1265 (
            .O(N__6820),
            .I(N__6817));
    Odrv12 I__1264 (
            .O(N__6817),
            .I(A_c_2));
    IoInMux I__1263 (
            .O(N__6814),
            .I(N__6810));
    InMux I__1262 (
            .O(N__6813),
            .I(N__6807));
    LocalMux I__1261 (
            .O(N__6810),
            .I(N__6804));
    LocalMux I__1260 (
            .O(N__6807),
            .I(N__6801));
    Span12Mux_s4_v I__1259 (
            .O(N__6804),
            .I(N__6798));
    Span4Mux_h I__1258 (
            .O(N__6801),
            .I(N__6795));
    Span12Mux_v I__1257 (
            .O(N__6798),
            .I(N__6792));
    Span4Mux_v I__1256 (
            .O(N__6795),
            .I(N__6789));
    Span12Mux_h I__1255 (
            .O(N__6792),
            .I(N__6786));
    Sp12to4 I__1254 (
            .O(N__6789),
            .I(N__6783));
    Odrv12 I__1253 (
            .O(N__6786),
            .I(A_c_9));
    Odrv12 I__1252 (
            .O(N__6783),
            .I(A_c_9));
    SRMux I__1251 (
            .O(N__6778),
            .I(N__6775));
    LocalMux I__1250 (
            .O(N__6775),
            .I(N__6772));
    Span4Mux_h I__1249 (
            .O(N__6772),
            .I(N__6769));
    Odrv4 I__1248 (
            .O(N__6769),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    CascadeMux I__1247 (
            .O(N__6766),
            .I(\U712_CHIP_RAM.REFRESH_RST_cascade_ ));
    InMux I__1246 (
            .O(N__6763),
            .I(N__6756));
    InMux I__1245 (
            .O(N__6762),
            .I(N__6753));
    CascadeMux I__1244 (
            .O(N__6761),
            .I(N__6748));
    InMux I__1243 (
            .O(N__6760),
            .I(N__6744));
    InMux I__1242 (
            .O(N__6759),
            .I(N__6741));
    LocalMux I__1241 (
            .O(N__6756),
            .I(N__6731));
    LocalMux I__1240 (
            .O(N__6753),
            .I(N__6731));
    InMux I__1239 (
            .O(N__6752),
            .I(N__6728));
    InMux I__1238 (
            .O(N__6751),
            .I(N__6721));
    InMux I__1237 (
            .O(N__6748),
            .I(N__6721));
    InMux I__1236 (
            .O(N__6747),
            .I(N__6721));
    LocalMux I__1235 (
            .O(N__6744),
            .I(N__6718));
    LocalMux I__1234 (
            .O(N__6741),
            .I(N__6715));
    InMux I__1233 (
            .O(N__6740),
            .I(N__6710));
    InMux I__1232 (
            .O(N__6739),
            .I(N__6710));
    InMux I__1231 (
            .O(N__6738),
            .I(N__6707));
    InMux I__1230 (
            .O(N__6737),
            .I(N__6704));
    InMux I__1229 (
            .O(N__6736),
            .I(N__6701));
    Span4Mux_h I__1228 (
            .O(N__6731),
            .I(N__6694));
    LocalMux I__1227 (
            .O(N__6728),
            .I(N__6694));
    LocalMux I__1226 (
            .O(N__6721),
            .I(N__6694));
    Span4Mux_v I__1225 (
            .O(N__6718),
            .I(N__6689));
    Span4Mux_v I__1224 (
            .O(N__6715),
            .I(N__6689));
    LocalMux I__1223 (
            .O(N__6710),
            .I(N__6686));
    LocalMux I__1222 (
            .O(N__6707),
            .I(N__6681));
    LocalMux I__1221 (
            .O(N__6704),
            .I(N__6681));
    LocalMux I__1220 (
            .O(N__6701),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1219 (
            .O(N__6694),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1218 (
            .O(N__6689),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1217 (
            .O(N__6686),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv12 I__1216 (
            .O(N__6681),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CascadeMux I__1215 (
            .O(N__6670),
            .I(N__6666));
    InMux I__1214 (
            .O(N__6669),
            .I(N__6662));
    InMux I__1213 (
            .O(N__6666),
            .I(N__6658));
    InMux I__1212 (
            .O(N__6665),
            .I(N__6655));
    LocalMux I__1211 (
            .O(N__6662),
            .I(N__6648));
    InMux I__1210 (
            .O(N__6661),
            .I(N__6645));
    LocalMux I__1209 (
            .O(N__6658),
            .I(N__6642));
    LocalMux I__1208 (
            .O(N__6655),
            .I(N__6639));
    InMux I__1207 (
            .O(N__6654),
            .I(N__6636));
    InMux I__1206 (
            .O(N__6653),
            .I(N__6633));
    InMux I__1205 (
            .O(N__6652),
            .I(N__6628));
    InMux I__1204 (
            .O(N__6651),
            .I(N__6628));
    Odrv4 I__1203 (
            .O(N__6648),
            .I(\U712_CHIP_RAM.N_595 ));
    LocalMux I__1202 (
            .O(N__6645),
            .I(\U712_CHIP_RAM.N_595 ));
    Odrv4 I__1201 (
            .O(N__6642),
            .I(\U712_CHIP_RAM.N_595 ));
    Odrv4 I__1200 (
            .O(N__6639),
            .I(\U712_CHIP_RAM.N_595 ));
    LocalMux I__1199 (
            .O(N__6636),
            .I(\U712_CHIP_RAM.N_595 ));
    LocalMux I__1198 (
            .O(N__6633),
            .I(\U712_CHIP_RAM.N_595 ));
    LocalMux I__1197 (
            .O(N__6628),
            .I(\U712_CHIP_RAM.N_595 ));
    CEMux I__1196 (
            .O(N__6613),
            .I(N__6610));
    LocalMux I__1195 (
            .O(N__6610),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0 ));
    InMux I__1194 (
            .O(N__6607),
            .I(N__6604));
    LocalMux I__1193 (
            .O(N__6604),
            .I(\U712_REG_SM.N_443 ));
    CascadeMux I__1192 (
            .O(N__6601),
            .I(N__6597));
    InMux I__1191 (
            .O(N__6600),
            .I(N__6588));
    InMux I__1190 (
            .O(N__6597),
            .I(N__6588));
    InMux I__1189 (
            .O(N__6596),
            .I(N__6581));
    InMux I__1188 (
            .O(N__6595),
            .I(N__6581));
    InMux I__1187 (
            .O(N__6594),
            .I(N__6581));
    CascadeMux I__1186 (
            .O(N__6593),
            .I(N__6574));
    LocalMux I__1185 (
            .O(N__6588),
            .I(N__6568));
    LocalMux I__1184 (
            .O(N__6581),
            .I(N__6568));
    InMux I__1183 (
            .O(N__6580),
            .I(N__6565));
    InMux I__1182 (
            .O(N__6579),
            .I(N__6562));
    InMux I__1181 (
            .O(N__6578),
            .I(N__6559));
    InMux I__1180 (
            .O(N__6577),
            .I(N__6552));
    InMux I__1179 (
            .O(N__6574),
            .I(N__6552));
    InMux I__1178 (
            .O(N__6573),
            .I(N__6552));
    Span4Mux_v I__1177 (
            .O(N__6568),
            .I(N__6549));
    LocalMux I__1176 (
            .O(N__6565),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1175 (
            .O(N__6562),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1174 (
            .O(N__6559),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1173 (
            .O(N__6552),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1172 (
            .O(N__6549),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__1171 (
            .O(N__6538),
            .I(N__6531));
    InMux I__1170 (
            .O(N__6537),
            .I(N__6522));
    InMux I__1169 (
            .O(N__6536),
            .I(N__6522));
    InMux I__1168 (
            .O(N__6535),
            .I(N__6522));
    CascadeMux I__1167 (
            .O(N__6534),
            .I(N__6519));
    LocalMux I__1166 (
            .O(N__6531),
            .I(N__6516));
    CascadeMux I__1165 (
            .O(N__6530),
            .I(N__6513));
    CascadeMux I__1164 (
            .O(N__6529),
            .I(N__6509));
    LocalMux I__1163 (
            .O(N__6522),
            .I(N__6502));
    InMux I__1162 (
            .O(N__6519),
            .I(N__6499));
    Span4Mux_v I__1161 (
            .O(N__6516),
            .I(N__6496));
    InMux I__1160 (
            .O(N__6513),
            .I(N__6493));
    InMux I__1159 (
            .O(N__6512),
            .I(N__6490));
    InMux I__1158 (
            .O(N__6509),
            .I(N__6479));
    InMux I__1157 (
            .O(N__6508),
            .I(N__6479));
    InMux I__1156 (
            .O(N__6507),
            .I(N__6479));
    InMux I__1155 (
            .O(N__6506),
            .I(N__6479));
    InMux I__1154 (
            .O(N__6505),
            .I(N__6479));
    Span4Mux_v I__1153 (
            .O(N__6502),
            .I(N__6476));
    LocalMux I__1152 (
            .O(N__6499),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1151 (
            .O(N__6496),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1150 (
            .O(N__6493),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1149 (
            .O(N__6490),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1148 (
            .O(N__6479),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1147 (
            .O(N__6476),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    IoInMux I__1146 (
            .O(N__6463),
            .I(N__6459));
    IoInMux I__1145 (
            .O(N__6462),
            .I(N__6456));
    LocalMux I__1144 (
            .O(N__6459),
            .I(N__6453));
    LocalMux I__1143 (
            .O(N__6456),
            .I(N__6450));
    Span4Mux_s3_v I__1142 (
            .O(N__6453),
            .I(N__6447));
    Span4Mux_s3_v I__1141 (
            .O(N__6450),
            .I(N__6444));
    Sp12to4 I__1140 (
            .O(N__6447),
            .I(N__6441));
    Sp12to4 I__1139 (
            .O(N__6444),
            .I(N__6438));
    Span12Mux_s9_h I__1138 (
            .O(N__6441),
            .I(N__6435));
    Span12Mux_s10_h I__1137 (
            .O(N__6438),
            .I(N__6432));
    Span12Mux_v I__1136 (
            .O(N__6435),
            .I(N__6426));
    Span12Mux_v I__1135 (
            .O(N__6432),
            .I(N__6426));
    InMux I__1134 (
            .O(N__6431),
            .I(N__6423));
    Odrv12 I__1133 (
            .O(N__6426),
            .I(ASn_c));
    LocalMux I__1132 (
            .O(N__6423),
            .I(ASn_c));
    InMux I__1131 (
            .O(N__6418),
            .I(N__6412));
    InMux I__1130 (
            .O(N__6417),
            .I(N__6412));
    LocalMux I__1129 (
            .O(N__6412),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    IoInMux I__1128 (
            .O(N__6409),
            .I(N__6406));
    LocalMux I__1127 (
            .O(N__6406),
            .I(N__6403));
    Span4Mux_s3_v I__1126 (
            .O(N__6403),
            .I(N__6400));
    Span4Mux_v I__1125 (
            .O(N__6400),
            .I(N__6397));
    Span4Mux_v I__1124 (
            .O(N__6397),
            .I(N__6394));
    Odrv4 I__1123 (
            .O(N__6394),
            .I(RESETn_c_i));
    IoInMux I__1122 (
            .O(N__6391),
            .I(N__6388));
    LocalMux I__1121 (
            .O(N__6388),
            .I(N__6385));
    Span4Mux_s3_v I__1120 (
            .O(N__6385),
            .I(N__6382));
    Span4Mux_h I__1119 (
            .O(N__6382),
            .I(N__6379));
    Span4Mux_v I__1118 (
            .O(N__6379),
            .I(N__6376));
    Odrv4 I__1117 (
            .O(N__6376),
            .I(N_549));
    InMux I__1116 (
            .O(N__6373),
            .I(N__6369));
    InMux I__1115 (
            .O(N__6372),
            .I(N__6366));
    LocalMux I__1114 (
            .O(N__6369),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    LocalMux I__1113 (
            .O(N__6366),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__1112 (
            .O(N__6361),
            .I(bfn_11_5_0_));
    InMux I__1111 (
            .O(N__6358),
            .I(N__6354));
    InMux I__1110 (
            .O(N__6357),
            .I(N__6351));
    LocalMux I__1109 (
            .O(N__6354),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    LocalMux I__1108 (
            .O(N__6351),
            .I(\U712_CHIP_RAM.REFRESH5lto1 ));
    InMux I__1107 (
            .O(N__6346),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__1106 (
            .O(N__6343),
            .I(N__6339));
    InMux I__1105 (
            .O(N__6342),
            .I(N__6336));
    LocalMux I__1104 (
            .O(N__6339),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    LocalMux I__1103 (
            .O(N__6336),
            .I(\U712_CHIP_RAM.REFRESH5lto2 ));
    InMux I__1102 (
            .O(N__6331),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__1101 (
            .O(N__6328),
            .I(N__6324));
    InMux I__1100 (
            .O(N__6327),
            .I(N__6321));
    LocalMux I__1099 (
            .O(N__6324),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__1098 (
            .O(N__6321),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__1097 (
            .O(N__6316),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    CascadeMux I__1096 (
            .O(N__6313),
            .I(N__6309));
    InMux I__1095 (
            .O(N__6312),
            .I(N__6306));
    InMux I__1094 (
            .O(N__6309),
            .I(N__6303));
    LocalMux I__1093 (
            .O(N__6306),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__1092 (
            .O(N__6303),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__1091 (
            .O(N__6298),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__1090 (
            .O(N__6295),
            .I(N__6292));
    LocalMux I__1089 (
            .O(N__6292),
            .I(\U712_REG_SM.STATE_COUNT_srsts_i_i_i_a2_0_0_0 ));
    InMux I__1088 (
            .O(N__6289),
            .I(N__6283));
    InMux I__1087 (
            .O(N__6288),
            .I(N__6276));
    InMux I__1086 (
            .O(N__6287),
            .I(N__6276));
    InMux I__1085 (
            .O(N__6286),
            .I(N__6276));
    LocalMux I__1084 (
            .O(N__6283),
            .I(N__6269));
    LocalMux I__1083 (
            .O(N__6276),
            .I(N__6269));
    InMux I__1082 (
            .O(N__6275),
            .I(N__6264));
    InMux I__1081 (
            .O(N__6274),
            .I(N__6264));
    Odrv12 I__1080 (
            .O(N__6269),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1079 (
            .O(N__6264),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    InMux I__1078 (
            .O(N__6259),
            .I(N__6256));
    LocalMux I__1077 (
            .O(N__6256),
            .I(N__6249));
    InMux I__1076 (
            .O(N__6255),
            .I(N__6242));
    InMux I__1075 (
            .O(N__6254),
            .I(N__6242));
    InMux I__1074 (
            .O(N__6253),
            .I(N__6242));
    InMux I__1073 (
            .O(N__6252),
            .I(N__6237));
    Sp12to4 I__1072 (
            .O(N__6249),
            .I(N__6232));
    LocalMux I__1071 (
            .O(N__6242),
            .I(N__6232));
    InMux I__1070 (
            .O(N__6241),
            .I(N__6227));
    InMux I__1069 (
            .O(N__6240),
            .I(N__6227));
    LocalMux I__1068 (
            .O(N__6237),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    Odrv12 I__1067 (
            .O(N__6232),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    LocalMux I__1066 (
            .O(N__6227),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    InMux I__1065 (
            .O(N__6220),
            .I(N__6213));
    InMux I__1064 (
            .O(N__6219),
            .I(N__6213));
    InMux I__1063 (
            .O(N__6218),
            .I(N__6210));
    LocalMux I__1062 (
            .O(N__6213),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__1061 (
            .O(N__6210),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__1060 (
            .O(N__6205),
            .I(N__6202));
    LocalMux I__1059 (
            .O(N__6202),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    InMux I__1058 (
            .O(N__6199),
            .I(N__6196));
    LocalMux I__1057 (
            .O(N__6196),
            .I(N__6192));
    InMux I__1056 (
            .O(N__6195),
            .I(N__6189));
    Odrv12 I__1055 (
            .O(N__6192),
            .I(\U712_REG_SM.START_RST_0_sqmuxa ));
    LocalMux I__1054 (
            .O(N__6189),
            .I(\U712_REG_SM.START_RST_0_sqmuxa ));
    InMux I__1053 (
            .O(N__6184),
            .I(N__6181));
    LocalMux I__1052 (
            .O(N__6181),
            .I(\U712_REG_SM.un1_STATE_COUNT_4_i_i_0_0 ));
    InMux I__1051 (
            .O(N__6178),
            .I(N__6175));
    LocalMux I__1050 (
            .O(N__6175),
            .I(\U712_REG_SM.DS_EN_RNOZ0Z_0 ));
    CascadeMux I__1049 (
            .O(N__6172),
            .I(N__6169));
    InMux I__1048 (
            .O(N__6169),
            .I(N__6166));
    LocalMux I__1047 (
            .O(N__6166),
            .I(N__6163));
    Odrv4 I__1046 (
            .O(N__6163),
            .I(\U712_REG_SM.N_515 ));
    InMux I__1045 (
            .O(N__6160),
            .I(N__6157));
    LocalMux I__1044 (
            .O(N__6157),
            .I(N__6154));
    Odrv4 I__1043 (
            .O(N__6154),
            .I(\U712_CHIP_RAM.N_537 ));
    InMux I__1042 (
            .O(N__6151),
            .I(N__6147));
    InMux I__1041 (
            .O(N__6150),
            .I(N__6142));
    LocalMux I__1040 (
            .O(N__6147),
            .I(N__6139));
    InMux I__1039 (
            .O(N__6146),
            .I(N__6136));
    InMux I__1038 (
            .O(N__6145),
            .I(N__6133));
    LocalMux I__1037 (
            .O(N__6142),
            .I(N__6130));
    Span4Mux_v I__1036 (
            .O(N__6139),
            .I(N__6125));
    LocalMux I__1035 (
            .O(N__6136),
            .I(N__6125));
    LocalMux I__1034 (
            .O(N__6133),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    Odrv4 I__1033 (
            .O(N__6130),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    Odrv4 I__1032 (
            .O(N__6125),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    InMux I__1031 (
            .O(N__6118),
            .I(N__6115));
    LocalMux I__1030 (
            .O(N__6115),
            .I(N__6112));
    Odrv4 I__1029 (
            .O(N__6112),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0_0 ));
    InMux I__1028 (
            .O(N__6109),
            .I(N__6098));
    InMux I__1027 (
            .O(N__6108),
            .I(N__6098));
    CascadeMux I__1026 (
            .O(N__6107),
            .I(N__6094));
    CascadeMux I__1025 (
            .O(N__6106),
            .I(N__6090));
    InMux I__1024 (
            .O(N__6105),
            .I(N__6083));
    InMux I__1023 (
            .O(N__6104),
            .I(N__6077));
    InMux I__1022 (
            .O(N__6103),
            .I(N__6077));
    LocalMux I__1021 (
            .O(N__6098),
            .I(N__6074));
    InMux I__1020 (
            .O(N__6097),
            .I(N__6071));
    InMux I__1019 (
            .O(N__6094),
            .I(N__6068));
    InMux I__1018 (
            .O(N__6093),
            .I(N__6063));
    InMux I__1017 (
            .O(N__6090),
            .I(N__6063));
    InMux I__1016 (
            .O(N__6089),
            .I(N__6056));
    InMux I__1015 (
            .O(N__6088),
            .I(N__6056));
    CascadeMux I__1014 (
            .O(N__6087),
            .I(N__6053));
    CascadeMux I__1013 (
            .O(N__6086),
            .I(N__6049));
    LocalMux I__1012 (
            .O(N__6083),
            .I(N__6045));
    InMux I__1011 (
            .O(N__6082),
            .I(N__6042));
    LocalMux I__1010 (
            .O(N__6077),
            .I(N__6039));
    Span4Mux_v I__1009 (
            .O(N__6074),
            .I(N__6032));
    LocalMux I__1008 (
            .O(N__6071),
            .I(N__6032));
    LocalMux I__1007 (
            .O(N__6068),
            .I(N__6032));
    LocalMux I__1006 (
            .O(N__6063),
            .I(N__6029));
    InMux I__1005 (
            .O(N__6062),
            .I(N__6026));
    InMux I__1004 (
            .O(N__6061),
            .I(N__6023));
    LocalMux I__1003 (
            .O(N__6056),
            .I(N__6020));
    InMux I__1002 (
            .O(N__6053),
            .I(N__6017));
    InMux I__1001 (
            .O(N__6052),
            .I(N__6014));
    InMux I__1000 (
            .O(N__6049),
            .I(N__6009));
    InMux I__999 (
            .O(N__6048),
            .I(N__6009));
    Span4Mux_v I__998 (
            .O(N__6045),
            .I(N__5998));
    LocalMux I__997 (
            .O(N__6042),
            .I(N__5998));
    Span4Mux_v I__996 (
            .O(N__6039),
            .I(N__5998));
    Span4Mux_h I__995 (
            .O(N__6032),
            .I(N__5998));
    Span4Mux_v I__994 (
            .O(N__6029),
            .I(N__5998));
    LocalMux I__993 (
            .O(N__6026),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__992 (
            .O(N__6023),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__991 (
            .O(N__6020),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__990 (
            .O(N__6017),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__989 (
            .O(N__6014),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__988 (
            .O(N__6009),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__987 (
            .O(N__5998),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    CascadeMux I__986 (
            .O(N__5983),
            .I(N__5979));
    InMux I__985 (
            .O(N__5982),
            .I(N__5972));
    InMux I__984 (
            .O(N__5979),
            .I(N__5969));
    InMux I__983 (
            .O(N__5978),
            .I(N__5965));
    CascadeMux I__982 (
            .O(N__5977),
            .I(N__5959));
    CascadeMux I__981 (
            .O(N__5976),
            .I(N__5955));
    CascadeMux I__980 (
            .O(N__5975),
            .I(N__5949));
    LocalMux I__979 (
            .O(N__5972),
            .I(N__5943));
    LocalMux I__978 (
            .O(N__5969),
            .I(N__5943));
    InMux I__977 (
            .O(N__5968),
            .I(N__5938));
    LocalMux I__976 (
            .O(N__5965),
            .I(N__5935));
    InMux I__975 (
            .O(N__5964),
            .I(N__5928));
    InMux I__974 (
            .O(N__5963),
            .I(N__5928));
    InMux I__973 (
            .O(N__5962),
            .I(N__5928));
    InMux I__972 (
            .O(N__5959),
            .I(N__5922));
    InMux I__971 (
            .O(N__5958),
            .I(N__5915));
    InMux I__970 (
            .O(N__5955),
            .I(N__5915));
    InMux I__969 (
            .O(N__5954),
            .I(N__5915));
    InMux I__968 (
            .O(N__5953),
            .I(N__5912));
    InMux I__967 (
            .O(N__5952),
            .I(N__5909));
    InMux I__966 (
            .O(N__5949),
            .I(N__5906));
    InMux I__965 (
            .O(N__5948),
            .I(N__5903));
    Span12Mux_h I__964 (
            .O(N__5943),
            .I(N__5900));
    InMux I__963 (
            .O(N__5942),
            .I(N__5895));
    InMux I__962 (
            .O(N__5941),
            .I(N__5895));
    LocalMux I__961 (
            .O(N__5938),
            .I(N__5890));
    Span4Mux_h I__960 (
            .O(N__5935),
            .I(N__5890));
    LocalMux I__959 (
            .O(N__5928),
            .I(N__5887));
    InMux I__958 (
            .O(N__5927),
            .I(N__5884));
    InMux I__957 (
            .O(N__5926),
            .I(N__5879));
    InMux I__956 (
            .O(N__5925),
            .I(N__5879));
    LocalMux I__955 (
            .O(N__5922),
            .I(N__5874));
    LocalMux I__954 (
            .O(N__5915),
            .I(N__5874));
    LocalMux I__953 (
            .O(N__5912),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__952 (
            .O(N__5909),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__951 (
            .O(N__5906),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__950 (
            .O(N__5903),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv12 I__949 (
            .O(N__5900),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__948 (
            .O(N__5895),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__947 (
            .O(N__5890),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__946 (
            .O(N__5887),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__945 (
            .O(N__5884),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__944 (
            .O(N__5879),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv12 I__943 (
            .O(N__5874),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__942 (
            .O(N__5851),
            .I(N__5847));
    InMux I__941 (
            .O(N__5850),
            .I(N__5844));
    LocalMux I__940 (
            .O(N__5847),
            .I(\U712_CHIP_RAM.N_703 ));
    LocalMux I__939 (
            .O(N__5844),
            .I(\U712_CHIP_RAM.N_703 ));
    CascadeMux I__938 (
            .O(N__5839),
            .I(\U712_CHIP_RAM.N_530_cascade_ ));
    InMux I__937 (
            .O(N__5836),
            .I(N__5831));
    InMux I__936 (
            .O(N__5835),
            .I(N__5826));
    InMux I__935 (
            .O(N__5834),
            .I(N__5823));
    LocalMux I__934 (
            .O(N__5831),
            .I(N__5820));
    InMux I__933 (
            .O(N__5830),
            .I(N__5817));
    InMux I__932 (
            .O(N__5829),
            .I(N__5814));
    LocalMux I__931 (
            .O(N__5826),
            .I(N__5809));
    LocalMux I__930 (
            .O(N__5823),
            .I(N__5809));
    Odrv4 I__929 (
            .O(N__5820),
            .I(\U712_CHIP_RAM.N_600 ));
    LocalMux I__928 (
            .O(N__5817),
            .I(\U712_CHIP_RAM.N_600 ));
    LocalMux I__927 (
            .O(N__5814),
            .I(\U712_CHIP_RAM.N_600 ));
    Odrv4 I__926 (
            .O(N__5809),
            .I(\U712_CHIP_RAM.N_600 ));
    CascadeMux I__925 (
            .O(N__5800),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_ ));
    CEMux I__924 (
            .O(N__5797),
            .I(N__5794));
    LocalMux I__923 (
            .O(N__5794),
            .I(N__5791));
    Span4Mux_h I__922 (
            .O(N__5791),
            .I(N__5788));
    Odrv4 I__921 (
            .O(N__5788),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0 ));
    InMux I__920 (
            .O(N__5785),
            .I(N__5781));
    InMux I__919 (
            .O(N__5784),
            .I(N__5778));
    LocalMux I__918 (
            .O(N__5781),
            .I(N__5775));
    LocalMux I__917 (
            .O(N__5778),
            .I(N__5772));
    Span4Mux_v I__916 (
            .O(N__5775),
            .I(N__5769));
    Span4Mux_v I__915 (
            .O(N__5772),
            .I(N__5766));
    Sp12to4 I__914 (
            .O(N__5769),
            .I(N__5763));
    Span4Mux_h I__913 (
            .O(N__5766),
            .I(N__5760));
    Span12Mux_h I__912 (
            .O(N__5763),
            .I(N__5755));
    Sp12to4 I__911 (
            .O(N__5760),
            .I(N__5755));
    Span12Mux_v I__910 (
            .O(N__5755),
            .I(N__5752));
    Odrv12 I__909 (
            .O(N__5752),
            .I(AWEn_c));
    InMux I__908 (
            .O(N__5749),
            .I(N__5746));
    LocalMux I__907 (
            .O(N__5746),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ));
    IoInMux I__906 (
            .O(N__5743),
            .I(N__5740));
    LocalMux I__905 (
            .O(N__5740),
            .I(N__5737));
    IoSpan4Mux I__904 (
            .O(N__5737),
            .I(N__5734));
    Span4Mux_s2_v I__903 (
            .O(N__5734),
            .I(N__5731));
    Sp12to4 I__902 (
            .O(N__5731),
            .I(N__5727));
    InMux I__901 (
            .O(N__5730),
            .I(N__5724));
    Odrv12 I__900 (
            .O(N__5727),
            .I(DBDIR_c));
    LocalMux I__899 (
            .O(N__5724),
            .I(DBDIR_c));
    InMux I__898 (
            .O(N__5719),
            .I(N__5716));
    LocalMux I__897 (
            .O(N__5716),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ));
    InMux I__896 (
            .O(N__5713),
            .I(N__5710));
    LocalMux I__895 (
            .O(N__5710),
            .I(\U712_CHIP_RAM.DBENn_8_0 ));
    InMux I__894 (
            .O(N__5707),
            .I(N__5703));
    InMux I__893 (
            .O(N__5706),
            .I(N__5700));
    LocalMux I__892 (
            .O(N__5703),
            .I(\U712_REG_SM.START_RSTZ0 ));
    LocalMux I__891 (
            .O(N__5700),
            .I(\U712_REG_SM.START_RSTZ0 ));
    CascadeMux I__890 (
            .O(N__5695),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_ ));
    IoInMux I__889 (
            .O(N__5692),
            .I(N__5689));
    LocalMux I__888 (
            .O(N__5689),
            .I(N__5686));
    Span4Mux_s3_v I__887 (
            .O(N__5686),
            .I(N__5683));
    Sp12to4 I__886 (
            .O(N__5683),
            .I(N__5680));
    Span12Mux_h I__885 (
            .O(N__5680),
            .I(N__5677));
    Span12Mux_v I__884 (
            .O(N__5677),
            .I(N__5673));
    InMux I__883 (
            .O(N__5676),
            .I(N__5670));
    Odrv12 I__882 (
            .O(N__5673),
            .I(LATCH_CLK_c));
    LocalMux I__881 (
            .O(N__5670),
            .I(LATCH_CLK_c));
    CascadeMux I__880 (
            .O(N__5665),
            .I(N__5661));
    InMux I__879 (
            .O(N__5664),
            .I(N__5658));
    InMux I__878 (
            .O(N__5661),
            .I(N__5655));
    LocalMux I__877 (
            .O(N__5658),
            .I(\U712_CHIP_RAM.N_528 ));
    LocalMux I__876 (
            .O(N__5655),
            .I(\U712_CHIP_RAM.N_528 ));
    InMux I__875 (
            .O(N__5650),
            .I(N__5647));
    LocalMux I__874 (
            .O(N__5647),
            .I(N__5641));
    InMux I__873 (
            .O(N__5646),
            .I(N__5638));
    InMux I__872 (
            .O(N__5645),
            .I(N__5633));
    InMux I__871 (
            .O(N__5644),
            .I(N__5633));
    Span4Mux_h I__870 (
            .O(N__5641),
            .I(N__5630));
    LocalMux I__869 (
            .O(N__5638),
            .I(N__5625));
    LocalMux I__868 (
            .O(N__5633),
            .I(N__5625));
    Odrv4 I__867 (
            .O(N__5630),
            .I(DBR_SYNCZ0Z_1));
    Odrv12 I__866 (
            .O(N__5625),
            .I(DBR_SYNCZ0Z_1));
    CascadeMux I__865 (
            .O(N__5620),
            .I(\U712_REG_SM.N_482_cascade_ ));
    InMux I__864 (
            .O(N__5617),
            .I(N__5614));
    LocalMux I__863 (
            .O(N__5614),
            .I(N__5611));
    Span4Mux_v I__862 (
            .O(N__5611),
            .I(N__5608));
    Span4Mux_h I__861 (
            .O(N__5608),
            .I(N__5604));
    IoInMux I__860 (
            .O(N__5607),
            .I(N__5601));
    Sp12to4 I__859 (
            .O(N__5604),
            .I(N__5598));
    LocalMux I__858 (
            .O(N__5601),
            .I(N__5595));
    Span12Mux_v I__857 (
            .O(N__5598),
            .I(N__5592));
    IoSpan4Mux I__856 (
            .O(N__5595),
            .I(N__5589));
    Odrv12 I__855 (
            .O(N__5592),
            .I(RAMENn_c));
    Odrv4 I__854 (
            .O(N__5589),
            .I(RAMENn_c));
    CascadeMux I__853 (
            .O(N__5584),
            .I(N__5581));
    InMux I__852 (
            .O(N__5581),
            .I(N__5578));
    LocalMux I__851 (
            .O(N__5578),
            .I(N__5575));
    Odrv4 I__850 (
            .O(N__5575),
            .I(\U712_CHIP_RAM.N_527 ));
    InMux I__849 (
            .O(N__5572),
            .I(N__5569));
    LocalMux I__848 (
            .O(N__5569),
            .I(N__5566));
    Span4Mux_v I__847 (
            .O(N__5566),
            .I(N__5562));
    InMux I__846 (
            .O(N__5565),
            .I(N__5559));
    Sp12to4 I__845 (
            .O(N__5562),
            .I(N__5554));
    LocalMux I__844 (
            .O(N__5559),
            .I(N__5554));
    Span12Mux_h I__843 (
            .O(N__5554),
            .I(N__5551));
    Span12Mux_v I__842 (
            .O(N__5551),
            .I(N__5548));
    Odrv12 I__841 (
            .O(N__5548),
            .I(TSn_c));
    InMux I__840 (
            .O(N__5545),
            .I(N__5542));
    LocalMux I__839 (
            .O(N__5542),
            .I(N__5537));
    InMux I__838 (
            .O(N__5541),
            .I(N__5534));
    InMux I__837 (
            .O(N__5540),
            .I(N__5531));
    Odrv4 I__836 (
            .O(N__5537),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__835 (
            .O(N__5534),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__834 (
            .O(N__5531),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__833 (
            .O(N__5524),
            .I(N__5520));
    InMux I__832 (
            .O(N__5523),
            .I(N__5517));
    LocalMux I__831 (
            .O(N__5520),
            .I(N__5514));
    LocalMux I__830 (
            .O(N__5517),
            .I(\U712_CHIP_RAM.N_553 ));
    Odrv12 I__829 (
            .O(N__5514),
            .I(\U712_CHIP_RAM.N_553 ));
    CascadeMux I__828 (
            .O(N__5509),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_ ));
    InMux I__827 (
            .O(N__5506),
            .I(N__5503));
    LocalMux I__826 (
            .O(N__5503),
            .I(\U712_CHIP_RAM.N_597 ));
    CascadeMux I__825 (
            .O(N__5500),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_ ));
    CascadeMux I__824 (
            .O(N__5497),
            .I(\U712_REG_SM.N_429_cascade_ ));
    CascadeMux I__823 (
            .O(N__5494),
            .I(\U712_REG_SM.N_511_cascade_ ));
    InMux I__822 (
            .O(N__5491),
            .I(N__5488));
    LocalMux I__821 (
            .O(N__5488),
            .I(N__5485));
    Span4Mux_h I__820 (
            .O(N__5485),
            .I(N__5482));
    Odrv4 I__819 (
            .O(N__5482),
            .I(\U712_REG_SM.N_694 ));
    InMux I__818 (
            .O(N__5479),
            .I(N__5476));
    LocalMux I__817 (
            .O(N__5476),
            .I(N__5473));
    Span4Mux_h I__816 (
            .O(N__5473),
            .I(N__5470));
    Odrv4 I__815 (
            .O(N__5470),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ));
    InMux I__814 (
            .O(N__5467),
            .I(N__5463));
    InMux I__813 (
            .O(N__5466),
            .I(N__5460));
    LocalMux I__812 (
            .O(N__5463),
            .I(\U712_CHIP_RAM.N_700 ));
    LocalMux I__811 (
            .O(N__5460),
            .I(\U712_CHIP_RAM.N_700 ));
    InMux I__810 (
            .O(N__5455),
            .I(N__5452));
    LocalMux I__809 (
            .O(N__5452),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0_a2_0_1 ));
    InMux I__808 (
            .O(N__5449),
            .I(N__5442));
    CascadeMux I__807 (
            .O(N__5448),
            .I(N__5439));
    CascadeMux I__806 (
            .O(N__5447),
            .I(N__5436));
    InMux I__805 (
            .O(N__5446),
            .I(N__5433));
    CascadeMux I__804 (
            .O(N__5445),
            .I(N__5427));
    LocalMux I__803 (
            .O(N__5442),
            .I(N__5423));
    InMux I__802 (
            .O(N__5439),
            .I(N__5420));
    InMux I__801 (
            .O(N__5436),
            .I(N__5417));
    LocalMux I__800 (
            .O(N__5433),
            .I(N__5414));
    InMux I__799 (
            .O(N__5432),
            .I(N__5411));
    InMux I__798 (
            .O(N__5431),
            .I(N__5408));
    InMux I__797 (
            .O(N__5430),
            .I(N__5405));
    InMux I__796 (
            .O(N__5427),
            .I(N__5399));
    InMux I__795 (
            .O(N__5426),
            .I(N__5396));
    Span4Mux_v I__794 (
            .O(N__5423),
            .I(N__5393));
    LocalMux I__793 (
            .O(N__5420),
            .I(N__5386));
    LocalMux I__792 (
            .O(N__5417),
            .I(N__5386));
    Span4Mux_v I__791 (
            .O(N__5414),
            .I(N__5386));
    LocalMux I__790 (
            .O(N__5411),
            .I(N__5379));
    LocalMux I__789 (
            .O(N__5408),
            .I(N__5379));
    LocalMux I__788 (
            .O(N__5405),
            .I(N__5379));
    InMux I__787 (
            .O(N__5404),
            .I(N__5376));
    InMux I__786 (
            .O(N__5403),
            .I(N__5373));
    InMux I__785 (
            .O(N__5402),
            .I(N__5370));
    LocalMux I__784 (
            .O(N__5399),
            .I(\U712_CHIP_RAM.N_578 ));
    LocalMux I__783 (
            .O(N__5396),
            .I(\U712_CHIP_RAM.N_578 ));
    Odrv4 I__782 (
            .O(N__5393),
            .I(\U712_CHIP_RAM.N_578 ));
    Odrv4 I__781 (
            .O(N__5386),
            .I(\U712_CHIP_RAM.N_578 ));
    Odrv12 I__780 (
            .O(N__5379),
            .I(\U712_CHIP_RAM.N_578 ));
    LocalMux I__779 (
            .O(N__5376),
            .I(\U712_CHIP_RAM.N_578 ));
    LocalMux I__778 (
            .O(N__5373),
            .I(\U712_CHIP_RAM.N_578 ));
    LocalMux I__777 (
            .O(N__5370),
            .I(\U712_CHIP_RAM.N_578 ));
    InMux I__776 (
            .O(N__5353),
            .I(N__5350));
    LocalMux I__775 (
            .O(N__5350),
            .I(N__5343));
    InMux I__774 (
            .O(N__5349),
            .I(N__5337));
    InMux I__773 (
            .O(N__5348),
            .I(N__5332));
    InMux I__772 (
            .O(N__5347),
            .I(N__5332));
    InMux I__771 (
            .O(N__5346),
            .I(N__5329));
    Span4Mux_h I__770 (
            .O(N__5343),
            .I(N__5326));
    InMux I__769 (
            .O(N__5342),
            .I(N__5323));
    InMux I__768 (
            .O(N__5341),
            .I(N__5320));
    InMux I__767 (
            .O(N__5340),
            .I(N__5317));
    LocalMux I__766 (
            .O(N__5337),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__765 (
            .O(N__5332),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__764 (
            .O(N__5329),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    Odrv4 I__763 (
            .O(N__5326),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__762 (
            .O(N__5323),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__761 (
            .O(N__5320),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__760 (
            .O(N__5317),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__759 (
            .O(N__5302),
            .I(N__5299));
    LocalMux I__758 (
            .O(N__5299),
            .I(\U712_CHIP_RAM.N_405 ));
    InMux I__757 (
            .O(N__5296),
            .I(N__5291));
    InMux I__756 (
            .O(N__5295),
            .I(N__5288));
    InMux I__755 (
            .O(N__5294),
            .I(N__5285));
    LocalMux I__754 (
            .O(N__5291),
            .I(\U712_CHIP_RAM.N_699 ));
    LocalMux I__753 (
            .O(N__5288),
            .I(\U712_CHIP_RAM.N_699 ));
    LocalMux I__752 (
            .O(N__5285),
            .I(\U712_CHIP_RAM.N_699 ));
    CascadeMux I__751 (
            .O(N__5278),
            .I(\U712_CHIP_RAM.N_597_cascade_ ));
    CascadeMux I__750 (
            .O(N__5275),
            .I(N__5272));
    InMux I__749 (
            .O(N__5272),
            .I(N__5269));
    LocalMux I__748 (
            .O(N__5269),
            .I(N__5266));
    Odrv4 I__747 (
            .O(N__5266),
            .I(\U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0 ));
    InMux I__746 (
            .O(N__5263),
            .I(N__5260));
    LocalMux I__745 (
            .O(N__5260),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    IoInMux I__744 (
            .O(N__5257),
            .I(N__5253));
    InMux I__743 (
            .O(N__5256),
            .I(N__5250));
    LocalMux I__742 (
            .O(N__5253),
            .I(N__5247));
    LocalMux I__741 (
            .O(N__5250),
            .I(N__5244));
    IoSpan4Mux I__740 (
            .O(N__5247),
            .I(N__5241));
    Span12Mux_h I__739 (
            .O(N__5244),
            .I(N__5238));
    IoSpan4Mux I__738 (
            .O(N__5241),
            .I(N__5235));
    Span12Mux_v I__737 (
            .O(N__5238),
            .I(N__5232));
    IoSpan4Mux I__736 (
            .O(N__5235),
            .I(N__5229));
    Odrv12 I__735 (
            .O(N__5232),
            .I(C1_c));
    Odrv4 I__734 (
            .O(N__5229),
            .I(C1_c));
    InMux I__733 (
            .O(N__5224),
            .I(N__5221));
    LocalMux I__732 (
            .O(N__5221),
            .I(N__5218));
    Odrv4 I__731 (
            .O(N__5218),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    CascadeMux I__730 (
            .O(N__5215),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_ ));
    InMux I__729 (
            .O(N__5212),
            .I(N__5209));
    LocalMux I__728 (
            .O(N__5209),
            .I(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ));
    InMux I__727 (
            .O(N__5206),
            .I(N__5202));
    CascadeMux I__726 (
            .O(N__5205),
            .I(N__5199));
    LocalMux I__725 (
            .O(N__5202),
            .I(N__5195));
    InMux I__724 (
            .O(N__5199),
            .I(N__5192));
    InMux I__723 (
            .O(N__5198),
            .I(N__5189));
    Span4Mux_h I__722 (
            .O(N__5195),
            .I(N__5186));
    LocalMux I__721 (
            .O(N__5192),
            .I(N__5181));
    LocalMux I__720 (
            .O(N__5189),
            .I(N__5181));
    Odrv4 I__719 (
            .O(N__5186),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__718 (
            .O(N__5181),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__717 (
            .O(N__5176),
            .I(N__5173));
    LocalMux I__716 (
            .O(N__5173),
            .I(N__5170));
    Odrv12 I__715 (
            .O(N__5170),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ));
    CascadeMux I__714 (
            .O(N__5167),
            .I(N__5164));
    InMux I__713 (
            .O(N__5164),
            .I(N__5159));
    InMux I__712 (
            .O(N__5163),
            .I(N__5154));
    InMux I__711 (
            .O(N__5162),
            .I(N__5151));
    LocalMux I__710 (
            .O(N__5159),
            .I(N__5146));
    InMux I__709 (
            .O(N__5158),
            .I(N__5141));
    InMux I__708 (
            .O(N__5157),
            .I(N__5141));
    LocalMux I__707 (
            .O(N__5154),
            .I(N__5134));
    LocalMux I__706 (
            .O(N__5151),
            .I(N__5134));
    InMux I__705 (
            .O(N__5150),
            .I(N__5129));
    InMux I__704 (
            .O(N__5149),
            .I(N__5129));
    Span4Mux_h I__703 (
            .O(N__5146),
            .I(N__5126));
    LocalMux I__702 (
            .O(N__5141),
            .I(N__5123));
    InMux I__701 (
            .O(N__5140),
            .I(N__5120));
    InMux I__700 (
            .O(N__5139),
            .I(N__5117));
    Odrv12 I__699 (
            .O(N__5134),
            .I(\U712_CHIP_RAM.N_589 ));
    LocalMux I__698 (
            .O(N__5129),
            .I(\U712_CHIP_RAM.N_589 ));
    Odrv4 I__697 (
            .O(N__5126),
            .I(\U712_CHIP_RAM.N_589 ));
    Odrv4 I__696 (
            .O(N__5123),
            .I(\U712_CHIP_RAM.N_589 ));
    LocalMux I__695 (
            .O(N__5120),
            .I(\U712_CHIP_RAM.N_589 ));
    LocalMux I__694 (
            .O(N__5117),
            .I(\U712_CHIP_RAM.N_589 ));
    CascadeMux I__693 (
            .O(N__5104),
            .I(N__5100));
    InMux I__692 (
            .O(N__5103),
            .I(N__5097));
    InMux I__691 (
            .O(N__5100),
            .I(N__5094));
    LocalMux I__690 (
            .O(N__5097),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    LocalMux I__689 (
            .O(N__5094),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    CascadeMux I__688 (
            .O(N__5089),
            .I(\U712_REG_SM.N_694_cascade_ ));
    CascadeMux I__687 (
            .O(N__5086),
            .I(\U712_REG_SM.N_522_cascade_ ));
    IoInMux I__686 (
            .O(N__5083),
            .I(N__5080));
    LocalMux I__685 (
            .O(N__5080),
            .I(N__5077));
    IoSpan4Mux I__684 (
            .O(N__5077),
            .I(N__5074));
    Span4Mux_s3_h I__683 (
            .O(N__5074),
            .I(N__5071));
    Span4Mux_h I__682 (
            .O(N__5071),
            .I(N__5068));
    Span4Mux_h I__681 (
            .O(N__5068),
            .I(N__5065));
    Span4Mux_h I__680 (
            .O(N__5065),
            .I(N__5061));
    InMux I__679 (
            .O(N__5064),
            .I(N__5058));
    Sp12to4 I__678 (
            .O(N__5061),
            .I(N__5053));
    LocalMux I__677 (
            .O(N__5058),
            .I(N__5053));
    Span12Mux_h I__676 (
            .O(N__5053),
            .I(N__5050));
    Span12Mux_v I__675 (
            .O(N__5050),
            .I(N__5047));
    Odrv12 I__674 (
            .O(N__5047),
            .I(C3_c));
    InMux I__673 (
            .O(N__5044),
            .I(N__5041));
    LocalMux I__672 (
            .O(N__5041),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__671 (
            .O(N__5038),
            .I(N__5034));
    InMux I__670 (
            .O(N__5037),
            .I(N__5031));
    LocalMux I__669 (
            .O(N__5034),
            .I(\U712_CHIP_RAM.N_697 ));
    LocalMux I__668 (
            .O(N__5031),
            .I(\U712_CHIP_RAM.N_697 ));
    InMux I__667 (
            .O(N__5026),
            .I(N__5023));
    LocalMux I__666 (
            .O(N__5023),
            .I(N__5019));
    InMux I__665 (
            .O(N__5022),
            .I(N__5016));
    Span4Mux_h I__664 (
            .O(N__5019),
            .I(N__5013));
    LocalMux I__663 (
            .O(N__5016),
            .I(N__5010));
    Odrv4 I__662 (
            .O(N__5013),
            .I(\U712_CHIP_RAM.N_551 ));
    Odrv4 I__661 (
            .O(N__5010),
            .I(\U712_CHIP_RAM.N_551 ));
    CascadeMux I__660 (
            .O(N__5005),
            .I(N__4998));
    CascadeMux I__659 (
            .O(N__5004),
            .I(N__4995));
    CascadeMux I__658 (
            .O(N__5003),
            .I(N__4992));
    CascadeMux I__657 (
            .O(N__5002),
            .I(N__4989));
    InMux I__656 (
            .O(N__5001),
            .I(N__4986));
    InMux I__655 (
            .O(N__4998),
            .I(N__4981));
    InMux I__654 (
            .O(N__4995),
            .I(N__4981));
    InMux I__653 (
            .O(N__4992),
            .I(N__4975));
    InMux I__652 (
            .O(N__4989),
            .I(N__4975));
    LocalMux I__651 (
            .O(N__4986),
            .I(N__4967));
    LocalMux I__650 (
            .O(N__4981),
            .I(N__4967));
    InMux I__649 (
            .O(N__4980),
            .I(N__4964));
    LocalMux I__648 (
            .O(N__4975),
            .I(N__4961));
    InMux I__647 (
            .O(N__4974),
            .I(N__4956));
    InMux I__646 (
            .O(N__4973),
            .I(N__4956));
    InMux I__645 (
            .O(N__4972),
            .I(N__4953));
    Odrv4 I__644 (
            .O(N__4967),
            .I(\U712_CHIP_RAM.N_580 ));
    LocalMux I__643 (
            .O(N__4964),
            .I(\U712_CHIP_RAM.N_580 ));
    Odrv12 I__642 (
            .O(N__4961),
            .I(\U712_CHIP_RAM.N_580 ));
    LocalMux I__641 (
            .O(N__4956),
            .I(\U712_CHIP_RAM.N_580 ));
    LocalMux I__640 (
            .O(N__4953),
            .I(\U712_CHIP_RAM.N_580 ));
    InMux I__639 (
            .O(N__4942),
            .I(N__4939));
    LocalMux I__638 (
            .O(N__4939),
            .I(N__4936));
    Span4Mux_h I__637 (
            .O(N__4936),
            .I(N__4933));
    Odrv4 I__636 (
            .O(N__4933),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    InMux I__635 (
            .O(N__4930),
            .I(N__4927));
    LocalMux I__634 (
            .O(N__4927),
            .I(N__4924));
    Odrv4 I__633 (
            .O(N__4924),
            .I(\U712_CHIP_RAM.N_505 ));
    CascadeMux I__632 (
            .O(N__4921),
            .I(N__4918));
    InMux I__631 (
            .O(N__4918),
            .I(N__4915));
    LocalMux I__630 (
            .O(N__4915),
            .I(\U712_CHIP_RAM.N_437 ));
    InMux I__629 (
            .O(N__4912),
            .I(N__4909));
    LocalMux I__628 (
            .O(N__4909),
            .I(\U712_CHIP_RAM.N_587 ));
    InMux I__627 (
            .O(N__4906),
            .I(N__4903));
    LocalMux I__626 (
            .O(N__4903),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__625 (
            .O(N__4900),
            .I(N__4884));
    InMux I__624 (
            .O(N__4899),
            .I(N__4884));
    InMux I__623 (
            .O(N__4898),
            .I(N__4884));
    InMux I__622 (
            .O(N__4897),
            .I(N__4884));
    InMux I__621 (
            .O(N__4896),
            .I(N__4879));
    InMux I__620 (
            .O(N__4895),
            .I(N__4879));
    InMux I__619 (
            .O(N__4894),
            .I(N__4874));
    InMux I__618 (
            .O(N__4893),
            .I(N__4874));
    LocalMux I__617 (
            .O(N__4884),
            .I(\U712_CHIP_RAM.N_70 ));
    LocalMux I__616 (
            .O(N__4879),
            .I(\U712_CHIP_RAM.N_70 ));
    LocalMux I__615 (
            .O(N__4874),
            .I(\U712_CHIP_RAM.N_70 ));
    CEMux I__614 (
            .O(N__4867),
            .I(N__4863));
    CEMux I__613 (
            .O(N__4866),
            .I(N__4860));
    LocalMux I__612 (
            .O(N__4863),
            .I(N__4857));
    LocalMux I__611 (
            .O(N__4860),
            .I(N__4854));
    Span4Mux_h I__610 (
            .O(N__4857),
            .I(N__4851));
    Odrv4 I__609 (
            .O(N__4854),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv4 I__608 (
            .O(N__4851),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__607 (
            .O(N__4846),
            .I(N__4843));
    LocalMux I__606 (
            .O(N__4843),
            .I(N__4840));
    Span4Mux_v I__605 (
            .O(N__4840),
            .I(N__4837));
    Sp12to4 I__604 (
            .O(N__4837),
            .I(N__4834));
    Span12Mux_h I__603 (
            .O(N__4834),
            .I(N__4831));
    Odrv12 I__602 (
            .O(N__4831),
            .I(REGSPACEn_c));
    CascadeMux I__601 (
            .O(N__4828),
            .I(\U712_REG_SM.N_513_cascade_ ));
    InMux I__600 (
            .O(N__4825),
            .I(N__4816));
    InMux I__599 (
            .O(N__4824),
            .I(N__4805));
    InMux I__598 (
            .O(N__4823),
            .I(N__4802));
    InMux I__597 (
            .O(N__4822),
            .I(N__4797));
    InMux I__596 (
            .O(N__4821),
            .I(N__4797));
    InMux I__595 (
            .O(N__4820),
            .I(N__4792));
    InMux I__594 (
            .O(N__4819),
            .I(N__4792));
    LocalMux I__593 (
            .O(N__4816),
            .I(N__4789));
    InMux I__592 (
            .O(N__4815),
            .I(N__4786));
    InMux I__591 (
            .O(N__4814),
            .I(N__4783));
    InMux I__590 (
            .O(N__4813),
            .I(N__4778));
    InMux I__589 (
            .O(N__4812),
            .I(N__4778));
    InMux I__588 (
            .O(N__4811),
            .I(N__4775));
    InMux I__587 (
            .O(N__4810),
            .I(N__4768));
    InMux I__586 (
            .O(N__4809),
            .I(N__4768));
    InMux I__585 (
            .O(N__4808),
            .I(N__4768));
    LocalMux I__584 (
            .O(N__4805),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__583 (
            .O(N__4802),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__582 (
            .O(N__4797),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__581 (
            .O(N__4792),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__580 (
            .O(N__4789),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__579 (
            .O(N__4786),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__578 (
            .O(N__4783),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__577 (
            .O(N__4778),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__576 (
            .O(N__4775),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__575 (
            .O(N__4768),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__574 (
            .O(N__4747),
            .I(N__4744));
    LocalMux I__573 (
            .O(N__4744),
            .I(\U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1 ));
    CascadeMux I__572 (
            .O(N__4741),
            .I(\U712_CHIP_RAM.N_697_cascade_ ));
    InMux I__571 (
            .O(N__4738),
            .I(N__4735));
    LocalMux I__570 (
            .O(N__4735),
            .I(N__4732));
    Odrv4 I__569 (
            .O(N__4732),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2 ));
    CascadeMux I__568 (
            .O(N__4729),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2_cascade_ ));
    InMux I__567 (
            .O(N__4726),
            .I(N__4723));
    LocalMux I__566 (
            .O(N__4723),
            .I(\U712_CHIP_RAM.N_539 ));
    CascadeMux I__565 (
            .O(N__4720),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_ ));
    CEMux I__564 (
            .O(N__4717),
            .I(N__4714));
    LocalMux I__563 (
            .O(N__4714),
            .I(N__4711));
    Odrv4 I__562 (
            .O(N__4711),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0 ));
    InMux I__561 (
            .O(N__4708),
            .I(N__4705));
    LocalMux I__560 (
            .O(N__4705),
            .I(N__4698));
    InMux I__559 (
            .O(N__4704),
            .I(N__4695));
    InMux I__558 (
            .O(N__4703),
            .I(N__4692));
    InMux I__557 (
            .O(N__4702),
            .I(N__4687));
    InMux I__556 (
            .O(N__4701),
            .I(N__4687));
    Odrv4 I__555 (
            .O(N__4698),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__554 (
            .O(N__4695),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__553 (
            .O(N__4692),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__552 (
            .O(N__4687),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__551 (
            .O(N__4678),
            .I(\U712_CHIP_RAM.N_442_cascade_ ));
    InMux I__550 (
            .O(N__4675),
            .I(N__4672));
    LocalMux I__549 (
            .O(N__4672),
            .I(\U712_CHIP_RAM.BANK0_RNOZ0Z_3 ));
    CascadeMux I__548 (
            .O(N__4669),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ));
    InMux I__547 (
            .O(N__4666),
            .I(N__4663));
    LocalMux I__546 (
            .O(N__4663),
            .I(\U712_CHIP_RAM.BANK0_RNOZ0Z_1 ));
    InMux I__545 (
            .O(N__4660),
            .I(N__4657));
    LocalMux I__544 (
            .O(N__4657),
            .I(N__4654));
    Span4Mux_h I__543 (
            .O(N__4654),
            .I(N__4651));
    Span4Mux_v I__542 (
            .O(N__4651),
            .I(N__4648));
    Sp12to4 I__541 (
            .O(N__4648),
            .I(N__4645));
    Odrv12 I__540 (
            .O(N__4645),
            .I(A_c_20));
    InMux I__539 (
            .O(N__4642),
            .I(N__4639));
    LocalMux I__538 (
            .O(N__4639),
            .I(N__4636));
    Odrv12 I__537 (
            .O(N__4636),
            .I(\U712_CHIP_RAM.BANK0_RNOZ0Z_2 ));
    CascadeMux I__536 (
            .O(N__4633),
            .I(\U712_CHIP_RAM.N_605_cascade_ ));
    InMux I__535 (
            .O(N__4630),
            .I(N__4626));
    InMux I__534 (
            .O(N__4629),
            .I(N__4623));
    LocalMux I__533 (
            .O(N__4626),
            .I(N__4620));
    LocalMux I__532 (
            .O(N__4623),
            .I(\U712_CHIP_RAM.N_605 ));
    Odrv4 I__531 (
            .O(N__4620),
            .I(\U712_CHIP_RAM.N_605 ));
    CascadeMux I__530 (
            .O(N__4615),
            .I(\U712_CHIP_RAM.N_554_cascade_ ));
    IoInMux I__529 (
            .O(N__4612),
            .I(N__4609));
    LocalMux I__528 (
            .O(N__4609),
            .I(N__4606));
    Span4Mux_s1_v I__527 (
            .O(N__4606),
            .I(N__4603));
    Sp12to4 I__526 (
            .O(N__4603),
            .I(N__4600));
    Span12Mux_h I__525 (
            .O(N__4600),
            .I(N__4597));
    Span12Mux_v I__524 (
            .O(N__4597),
            .I(N__4593));
    InMux I__523 (
            .O(N__4596),
            .I(N__4590));
    Odrv12 I__522 (
            .O(N__4593),
            .I(BANK0_c));
    LocalMux I__521 (
            .O(N__4590),
            .I(BANK0_c));
    InMux I__520 (
            .O(N__4585),
            .I(N__4582));
    LocalMux I__519 (
            .O(N__4582),
            .I(\U712_CHIP_RAM.N_588 ));
    CascadeMux I__518 (
            .O(N__4579),
            .I(\U712_CHIP_RAM.N_553_cascade_ ));
    CascadeMux I__517 (
            .O(N__4576),
            .I(\U712_CHIP_RAM.N_437_cascade_ ));
    InMux I__516 (
            .O(N__4573),
            .I(N__4569));
    InMux I__515 (
            .O(N__4572),
            .I(N__4566));
    LocalMux I__514 (
            .O(N__4569),
            .I(\U712_CHIP_RAM.N_414 ));
    LocalMux I__513 (
            .O(N__4566),
            .I(\U712_CHIP_RAM.N_414 ));
    InMux I__512 (
            .O(N__4561),
            .I(N__4558));
    LocalMux I__511 (
            .O(N__4558),
            .I(\U712_CHIP_RAM.N_507 ));
    CascadeMux I__510 (
            .O(N__4555),
            .I(\U712_CHIP_RAM.N_507_cascade_ ));
    InMux I__509 (
            .O(N__4552),
            .I(N__4549));
    LocalMux I__508 (
            .O(N__4549),
            .I(N__4546));
    Odrv4 I__507 (
            .O(N__4546),
            .I(\U712_CHIP_RAM.N_506 ));
    CascadeMux I__506 (
            .O(N__4543),
            .I(N__4539));
    InMux I__505 (
            .O(N__4542),
            .I(N__4536));
    InMux I__504 (
            .O(N__4539),
            .I(N__4532));
    LocalMux I__503 (
            .O(N__4536),
            .I(N__4529));
    InMux I__502 (
            .O(N__4535),
            .I(N__4526));
    LocalMux I__501 (
            .O(N__4532),
            .I(\U712_CHIP_RAM.N_696 ));
    Odrv4 I__500 (
            .O(N__4529),
            .I(\U712_CHIP_RAM.N_696 ));
    LocalMux I__499 (
            .O(N__4526),
            .I(\U712_CHIP_RAM.N_696 ));
    InMux I__498 (
            .O(N__4519),
            .I(N__4516));
    LocalMux I__497 (
            .O(N__4516),
            .I(N__4513));
    Odrv4 I__496 (
            .O(N__4513),
            .I(\U712_CHIP_RAM.N_534 ));
    InMux I__495 (
            .O(N__4510),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__494 (
            .O(N__4507),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__493 (
            .O(N__4504),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__492 (
            .O(N__4501),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__491 (
            .O(N__4498),
            .I(N__4494));
    InMux I__490 (
            .O(N__4497),
            .I(N__4491));
    LocalMux I__489 (
            .O(N__4494),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__488 (
            .O(N__4491),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__487 (
            .O(N__4486),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__486 (
            .O(N__4483),
            .I(N__4479));
    InMux I__485 (
            .O(N__4482),
            .I(N__4476));
    LocalMux I__484 (
            .O(N__4479),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__483 (
            .O(N__4476),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__482 (
            .O(N__4471),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__481 (
            .O(N__4468),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    InMux I__480 (
            .O(N__4465),
            .I(N__4461));
    InMux I__479 (
            .O(N__4464),
            .I(N__4458));
    LocalMux I__478 (
            .O(N__4461),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__477 (
            .O(N__4458),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__476 (
            .O(N__4453),
            .I(N__4450));
    LocalMux I__475 (
            .O(N__4450),
            .I(N__4447));
    Span4Mux_h I__474 (
            .O(N__4447),
            .I(N__4444));
    Sp12to4 I__473 (
            .O(N__4444),
            .I(N__4441));
    Span12Mux_v I__472 (
            .O(N__4441),
            .I(N__4438));
    Odrv12 I__471 (
            .O(N__4438),
            .I(A_c_8));
    InMux I__470 (
            .O(N__4435),
            .I(N__4432));
    LocalMux I__469 (
            .O(N__4432),
            .I(N__4429));
    Span12Mux_v I__468 (
            .O(N__4429),
            .I(N__4426));
    Odrv12 I__467 (
            .O(N__4426),
            .I(A_c_15));
    CascadeMux I__466 (
            .O(N__4423),
            .I(\U712_CHIP_RAM.N_578_cascade_ ));
    InMux I__465 (
            .O(N__4420),
            .I(N__4417));
    LocalMux I__464 (
            .O(N__4417),
            .I(\U712_CHIP_RAM.N_545 ));
    CascadeMux I__463 (
            .O(N__4414),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER18_cascade_ ));
    CascadeMux I__462 (
            .O(N__4411),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_cascade_ ));
    InMux I__461 (
            .O(N__4408),
            .I(N__4405));
    LocalMux I__460 (
            .O(N__4405),
            .I(\U712_CHIP_RAM.N_552 ));
    CascadeMux I__459 (
            .O(N__4402),
            .I(\U712_CHIP_RAM.N_504_cascade_ ));
    InMux I__458 (
            .O(N__4399),
            .I(N__4396));
    LocalMux I__457 (
            .O(N__4396),
            .I(N__4393));
    Odrv4 I__456 (
            .O(N__4393),
            .I(\U712_CHIP_RAM.N_404 ));
    CascadeMux I__455 (
            .O(N__4390),
            .I(\U712_CHIP_RAM.N_404_cascade_ ));
    InMux I__454 (
            .O(N__4387),
            .I(N__4384));
    LocalMux I__453 (
            .O(N__4384),
            .I(N__4381));
    Span4Mux_v I__452 (
            .O(N__4381),
            .I(N__4378));
    Span4Mux_v I__451 (
            .O(N__4378),
            .I(N__4375));
    Sp12to4 I__450 (
            .O(N__4375),
            .I(N__4372));
    Odrv12 I__449 (
            .O(N__4372),
            .I(A_c_5));
    InMux I__448 (
            .O(N__4369),
            .I(N__4366));
    LocalMux I__447 (
            .O(N__4366),
            .I(N__4363));
    Span4Mux_v I__446 (
            .O(N__4363),
            .I(N__4360));
    Sp12to4 I__445 (
            .O(N__4360),
            .I(N__4357));
    Odrv12 I__444 (
            .O(N__4357),
            .I(A_c_12));
    InMux I__443 (
            .O(N__4354),
            .I(N__4351));
    LocalMux I__442 (
            .O(N__4351),
            .I(\U712_CHIP_RAM.N_591 ));
    IoInMux I__441 (
            .O(N__4348),
            .I(N__4345));
    LocalMux I__440 (
            .O(N__4345),
            .I(N__4342));
    Span12Mux_s9_v I__439 (
            .O(N__4342),
            .I(N__4339));
    Odrv12 I__438 (
            .O(N__4339),
            .I(VBENn_c));
    InMux I__437 (
            .O(N__4336),
            .I(N__4333));
    LocalMux I__436 (
            .O(N__4333),
            .I(N__4330));
    Span4Mux_v I__435 (
            .O(N__4330),
            .I(N__4327));
    Span4Mux_v I__434 (
            .O(N__4327),
            .I(N__4324));
    Sp12to4 I__433 (
            .O(N__4324),
            .I(N__4321));
    Odrv12 I__432 (
            .O(N__4321),
            .I(A_c_14));
    InMux I__431 (
            .O(N__4318),
            .I(N__4315));
    LocalMux I__430 (
            .O(N__4315),
            .I(N__4312));
    Span4Mux_v I__429 (
            .O(N__4312),
            .I(N__4309));
    Span4Mux_v I__428 (
            .O(N__4309),
            .I(N__4306));
    Sp12to4 I__427 (
            .O(N__4306),
            .I(N__4303));
    Odrv12 I__426 (
            .O(N__4303),
            .I(A_c_7));
    CascadeMux I__425 (
            .O(N__4300),
            .I(\U712_CHIP_RAM.N_543_cascade_ ));
    CascadeMux I__424 (
            .O(N__4297),
            .I(\U712_CHIP_RAM.N_322_cascade_ ));
    InMux I__423 (
            .O(N__4294),
            .I(N__4291));
    LocalMux I__422 (
            .O(N__4291),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0_0 ));
    InMux I__421 (
            .O(N__4288),
            .I(N__4285));
    LocalMux I__420 (
            .O(N__4285),
            .I(\U712_CHIP_RAM.CLK_EN_6_0_a3_0_a2_1 ));
    CascadeMux I__419 (
            .O(N__4282),
            .I(\U712_CHIP_RAM.N_599_cascade_ ));
    InMux I__418 (
            .O(N__4279),
            .I(N__4276));
    LocalMux I__417 (
            .O(N__4276),
            .I(\U712_CHIP_RAM.CLK_EN_6_0 ));
    IoInMux I__416 (
            .O(N__4273),
            .I(N__4270));
    LocalMux I__415 (
            .O(N__4270),
            .I(N__4267));
    Span4Mux_s1_v I__414 (
            .O(N__4267),
            .I(N__4264));
    Span4Mux_v I__413 (
            .O(N__4264),
            .I(N__4261));
    Span4Mux_v I__412 (
            .O(N__4261),
            .I(N__4258));
    Span4Mux_v I__411 (
            .O(N__4258),
            .I(N__4255));
    Odrv4 I__410 (
            .O(N__4255),
            .I(U712_CYCLE_TERM_TBIn_0_i));
    IoInMux I__409 (
            .O(N__4252),
            .I(N__4249));
    LocalMux I__408 (
            .O(N__4249),
            .I(N__4246));
    Span4Mux_s2_v I__407 (
            .O(N__4246),
            .I(N__4243));
    Span4Mux_v I__406 (
            .O(N__4243),
            .I(N__4240));
    Span4Mux_h I__405 (
            .O(N__4240),
            .I(N__4237));
    Odrv4 I__404 (
            .O(N__4237),
            .I(CLK80_PLL_i_i));
    IoInMux I__403 (
            .O(N__4234),
            .I(N__4231));
    LocalMux I__402 (
            .O(N__4231),
            .I(N__4228));
    IoSpan4Mux I__401 (
            .O(N__4228),
            .I(N__4225));
    Span4Mux_s3_h I__400 (
            .O(N__4225),
            .I(N__4222));
    Span4Mux_h I__399 (
            .O(N__4222),
            .I(N__4219));
    Odrv4 I__398 (
            .O(N__4219),
            .I(DBRn_c_i_0));
    IoInMux I__397 (
            .O(N__4216),
            .I(N__4213));
    LocalMux I__396 (
            .O(N__4213),
            .I(N__4210));
    Span12Mux_s10_h I__395 (
            .O(N__4210),
            .I(N__4207));
    Span12Mux_h I__394 (
            .O(N__4207),
            .I(N__4203));
    InMux I__393 (
            .O(N__4206),
            .I(N__4200));
    Odrv12 I__392 (
            .O(N__4203),
            .I(CLK_EN_c));
    LocalMux I__391 (
            .O(N__4200),
            .I(CLK_EN_c));
    InMux I__390 (
            .O(N__4195),
            .I(N__4191));
    InMux I__389 (
            .O(N__4194),
            .I(N__4188));
    LocalMux I__388 (
            .O(N__4191),
            .I(N__4183));
    LocalMux I__387 (
            .O(N__4188),
            .I(N__4183));
    Span12Mux_h I__386 (
            .O(N__4183),
            .I(N__4180));
    Span12Mux_v I__385 (
            .O(N__4180),
            .I(N__4177));
    Odrv12 I__384 (
            .O(N__4177),
            .I(DBRn_c));
    InMux I__383 (
            .O(N__4174),
            .I(N__4171));
    LocalMux I__382 (
            .O(N__4171),
            .I(N__4168));
    Odrv4 I__381 (
            .O(N__4168),
            .I(DBR_SYNCZ0Z_0));
    InMux I__380 (
            .O(N__4165),
            .I(N__4162));
    LocalMux I__379 (
            .O(N__4162),
            .I(N__4159));
    Span4Mux_v I__378 (
            .O(N__4159),
            .I(N__4156));
    Span4Mux_v I__377 (
            .O(N__4156),
            .I(N__4153));
    Sp12to4 I__376 (
            .O(N__4153),
            .I(N__4150));
    Odrv12 I__375 (
            .O(N__4150),
            .I(A_c_18));
    InMux I__374 (
            .O(N__4147),
            .I(N__4144));
    LocalMux I__373 (
            .O(N__4144),
            .I(N__4141));
    Span4Mux_v I__372 (
            .O(N__4141),
            .I(N__4138));
    Span4Mux_v I__371 (
            .O(N__4138),
            .I(N__4135));
    Sp12to4 I__370 (
            .O(N__4135),
            .I(N__4132));
    Odrv12 I__369 (
            .O(N__4132),
            .I(A_c_16));
    InMux I__368 (
            .O(N__4129),
            .I(N__4126));
    LocalMux I__367 (
            .O(N__4126),
            .I(N__4123));
    Span4Mux_v I__366 (
            .O(N__4123),
            .I(N__4120));
    Span4Mux_v I__365 (
            .O(N__4120),
            .I(N__4117));
    Sp12to4 I__364 (
            .O(N__4117),
            .I(N__4114));
    Odrv12 I__363 (
            .O(N__4114),
            .I(A_c_6));
    InMux I__362 (
            .O(N__4111),
            .I(N__4108));
    LocalMux I__361 (
            .O(N__4108),
            .I(N__4105));
    Odrv12 I__360 (
            .O(N__4105),
            .I(A_c_13));
    IoInMux I__359 (
            .O(N__4102),
            .I(N__4099));
    LocalMux I__358 (
            .O(N__4099),
            .I(N__4096));
    IoSpan4Mux I__357 (
            .O(N__4096),
            .I(N__4093));
    Span4Mux_s2_v I__356 (
            .O(N__4093),
            .I(N__4090));
    Sp12to4 I__355 (
            .O(N__4090),
            .I(N__4087));
    Span12Mux_v I__354 (
            .O(N__4087),
            .I(N__4084));
    Odrv12 I__353 (
            .O(N__4084),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__6861));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__6863));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__6865));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .I(N__6860));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__6862));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__6858));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__6859));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__5257),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__6409),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4234),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__5083),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUTn_RNI3QLB_LC_3_8_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_RNI3QLB_LC_3_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_OUTn_RNI3QLB_LC_3_8_7 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_RNI3QLB_LC_3_8_7  (
            .in0(N__7665),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7599),
            .lcout(U712_CYCLE_TERM_TBIn_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_5_1_2.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_5_1_2.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_5_1_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_5_1_2 (
            .in0(N__8803),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_5_9_4.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_5_9_4.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_5_9_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_5_9_4 (
            .in0(N__4194),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_10_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_5_10_7  (
            .in0(N__9285),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10279),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_6_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_6_6_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_6_6_6 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_6_6_6  (
            .in0(N__4206),
            .in1(N__4279),
            .in2(_gnd_net_),
            .in3(N__5479),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8787),
            .ce(),
            .sr(N__10259));
    defparam DBR_SYNC_1_LC_6_7_7.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_6_7_7.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_6_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_6_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4174),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8791),
            .ce(),
            .sr(N__10256));
    defparam DBR_SYNC_0_LC_6_9_5.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_6_9_5.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_6_9_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 DBR_SYNC_0_LC_6_9_5 (
            .in0(N__4195),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8797),
            .ce(),
            .sr(N__10244));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_7_4_0  (
            .in0(N__4165),
            .in1(N__4147),
            .in2(_gnd_net_),
            .in3(N__9035),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_7_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_7_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_7_5_3  (
            .in0(N__4129),
            .in1(N__4111),
            .in2(_gnd_net_),
            .in3(N__8997),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_3_LC_7_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_3_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_3_LC_7_5_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_3_LC_7_5_6  (
            .in0(N__9585),
            .in1(N__7178),
            .in2(_gnd_net_),
            .in3(N__5978),
            .lcout(\U712_CHIP_RAM.CLK_EN_6_0_a3_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_7_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_7_5_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_7_5_7  (
            .in0(N__4336),
            .in1(N__4318),
            .in2(_gnd_net_),
            .in3(N__8996),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_6_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_6_0  (
            .in0(N__4399),
            .in1(N__4630),
            .in2(N__5448),
            .in3(N__5348),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_543_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_7_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_7_6_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_7_6_1  (
            .in0(N__4294),
            .in1(N__4420),
            .in2(N__4300),
            .in3(N__5001),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_322_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_7_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_7_6_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__6151),
            .in2(N__4297),
            .in3(N__9002),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8782),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_7_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_7_6_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_1_LC_7_6_3  (
            .in0(N__4821),
            .in1(N__8026),
            .in2(N__5983),
            .in3(N__6109),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_7_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_2_LC_7_6_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_2_LC_7_6_5  (
            .in0(N__4822),
            .in1(N__7801),
            .in2(_gnd_net_),
            .in3(N__6108),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_599_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_6_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_7_6_6  (
            .in0(N__4288),
            .in1(N__5347),
            .in2(N__4282),
            .in3(N__5426),
            .lcout(\U712_CHIP_RAM.CLK_EN_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_7_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_LC_7_7_0 .LUT_INIT=16'b1010101010101110;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_LC_7_7_0  (
            .in0(N__4519),
            .in1(N__9633),
            .in2(N__7802),
            .in3(N__7161),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8788),
            .ce(N__4717),
            .sr(N__10250));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_1_LC_7_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_1_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_1_LC_7_7_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_1_LC_7_7_2  (
            .in0(N__7783),
            .in1(N__4972),
            .in2(N__6106),
            .in3(N__4812),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_504_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5PDS6_3_LC_7_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5PDS6_3_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5PDS6_3_LC_7_7_3 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5PDS6_3_LC_7_7_3  (
            .in0(N__4813),
            .in1(N__6093),
            .in2(N__4402),
            .in3(N__4535),
            .lcout(\U712_CHIP_RAM.N_414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI85LA2_4_LC_7_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI85LA2_4_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI85LA2_4_LC_7_7_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI85LA2_4_LC_7_7_4  (
            .in0(N__7782),
            .in1(N__5341),
            .in2(_gnd_net_),
            .in3(N__5402),
            .lcout(\U712_CHIP_RAM.N_696 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_7_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_7_8_1 .LUT_INIT=16'b0000001101000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_7_8_1  (
            .in0(N__4814),
            .in1(N__6097),
            .in2(N__5976),
            .in3(N__7793),
            .lcout(\U712_CHIP_RAM.N_404 ),
            .ltout(\U712_CHIP_RAM.N_404_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIM81M2_LC_7_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIM81M2_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIM81M2_LC_7_8_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIM81M2_LC_7_8_2  (
            .in0(N__5342),
            .in1(_gnd_net_),
            .in2(N__4390),
            .in3(N__4708),
            .lcout(\U712_CHIP_RAM.N_591 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_8_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_8_3  (
            .in0(N__5958),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4573),
            .lcout(\U712_CHIP_RAM.N_505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_7_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_7_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_7_8_4  (
            .in0(N__4387),
            .in1(N__4369),
            .in2(_gnd_net_),
            .in3(N__9022),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_7_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_7_8_5 .LUT_INIT=16'b1000110010001000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_7_8_5  (
            .in0(N__5954),
            .in1(N__7792),
            .in2(N__6107),
            .in3(N__7132),
            .lcout(\U712_CHIP_RAM.N_588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIF4EE6_LC_7_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIF4EE6_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIF4EE6_LC_7_9_1 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIF4EE6_LC_7_9_1  (
            .in0(N__4354),
            .in1(N__8025),
            .in2(N__5167),
            .in3(N__5446),
            .lcout(\U712_CHIP_RAM.N_551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a3_0_a2_LC_8_5_3 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a3_0_a2_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a3_0_a2_LC_8_5_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a3_0_a2_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(N__9616),
            .in2(_gnd_net_),
            .in3(N__10119),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_8_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_8_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_8_5_4  (
            .in0(N__4453),
            .in1(N__4435),
            .in2(_gnd_net_),
            .in3(N__9001),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_8_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_8_6_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_8_6_0  (
            .in0(N__4464),
            .in1(N__4482),
            .in2(_gnd_net_),
            .in3(N__4497),
            .lcout(\U712_CHIP_RAM.N_578 ),
            .ltout(\U712_CHIP_RAM.N_578_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_6_1 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_8_6_1  (
            .in0(N__5340),
            .in1(_gnd_net_),
            .in2(N__4423),
            .in3(N__4701),
            .lcout(\U712_CHIP_RAM.N_580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_6_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_6_2  (
            .in0(N__5206),
            .in1(N__8030),
            .in2(N__6670),
            .in3(N__6759),
            .lcout(\U712_CHIP_RAM.N_545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_6_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_6_3  (
            .in0(N__5982),
            .in1(N__6104),
            .in2(N__4543),
            .in3(N__4824),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_6_4 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_6_4  (
            .in0(N__4702),
            .in1(_gnd_net_),
            .in2(N__4414),
            .in3(N__8031),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8778),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_6_5 .LUT_INIT=16'b1100000011010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_6_5  (
            .in0(N__4408),
            .in1(N__6150),
            .in2(N__9161),
            .in3(N__5022),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8778),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIM2QU_3_LC_8_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIM2QU_3_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIM2QU_3_LC_8_6_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIM2QU_3_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(N__8032),
            .in2(_gnd_net_),
            .in3(N__4811),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMEP34_1_LC_8_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMEP34_1_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMEP34_1_LC_8_6_7 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIMEP34_1_LC_8_6_7  (
            .in0(N__7794),
            .in1(N__6103),
            .in2(N__4411),
            .in3(N__4980),
            .lcout(\U712_CHIP_RAM.N_506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_7_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__6062),
            .in2(_gnd_net_),
            .in3(N__5037),
            .lcout(\U712_CHIP_RAM.N_552 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_7_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_7_1  (
            .in0(N__4897),
            .in1(N__7800),
            .in2(_gnd_net_),
            .in3(N__4510),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__8783),
            .ce(N__4866),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_7_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__5953),
            .in2(_gnd_net_),
            .in3(N__4507),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_7_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_7_3  (
            .in0(N__4898),
            .in1(N__4823),
            .in2(_gnd_net_),
            .in3(N__4504),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__8783),
            .ce(N__4866),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_7_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_7_4  (
            .in0(N__4893),
            .in1(N__5349),
            .in2(_gnd_net_),
            .in3(N__4501),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__8783),
            .ce(N__4866),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_7_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_7_5  (
            .in0(N__4899),
            .in1(N__4498),
            .in2(_gnd_net_),
            .in3(N__4486),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__8783),
            .ce(N__4866),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_7_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_7_6  (
            .in0(N__4894),
            .in1(N__4483),
            .in2(_gnd_net_),
            .in3(N__4471),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__8783),
            .ce(N__4866),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_7_7  (
            .in0(N__4900),
            .in1(N__4465),
            .in2(_gnd_net_),
            .in3(N__4468),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8783),
            .ce(N__4866),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_0_LC_8_8_0 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_0_LC_8_8_0  (
            .in0(N__5830),
            .in1(N__6760),
            .in2(N__5003),
            .in3(N__5150),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_554_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_LC_8_8_1 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \U712_CHIP_RAM.BANK0_LC_8_8_1  (
            .in0(N__4596),
            .in1(N__5523),
            .in2(N__4615),
            .in3(N__4666),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8789),
            .ce(),
            .sr(N__10236));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_3_LC_8_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_3_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_3_LC_8_8_2 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_3_LC_8_8_2  (
            .in0(N__4912),
            .in1(N__4815),
            .in2(N__5002),
            .in3(N__4585),
            .lcout(\U712_CHIP_RAM.N_553 ),
            .ltout(\U712_CHIP_RAM.N_553_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_3_LC_8_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_3_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_3_LC_8_8_3 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_3_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4579),
            .in3(N__7988),
            .lcout(\U712_CHIP_RAM.N_437 ),
            .ltout(\U712_CHIP_RAM.N_437_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG9KPG_2_LC_8_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG9KPG_2_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIG9KPG_2_LC_8_8_4 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIG9KPG_2_LC_8_8_4  (
            .in0(N__4561),
            .in1(N__5432),
            .in2(N__4576),
            .in3(N__5149),
            .lcout(\U712_CHIP_RAM.N_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_2_LC_8_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_2_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_2_LC_8_8_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_2_LC_8_8_5  (
            .in0(N__5948),
            .in1(N__7989),
            .in2(_gnd_net_),
            .in3(N__4572),
            .lcout(\U712_CHIP_RAM.N_507 ),
            .ltout(\U712_CHIP_RAM.N_507_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_8_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_8_8_6 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_8_8_6  (
            .in0(N__6653),
            .in1(N__4738),
            .in2(N__4555),
            .in3(N__4552),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_8_9_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_8_9_0  (
            .in0(N__7143),
            .in1(N__4542),
            .in2(N__5975),
            .in3(N__4747),
            .lcout(\U712_CHIP_RAM.N_534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_3_LC_8_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_3_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_3_LC_8_9_1 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_3_LC_8_9_1  (
            .in0(N__5157),
            .in1(N__6747),
            .in2(_gnd_net_),
            .in3(N__5430),
            .lcout(\U712_CHIP_RAM.BANK0_RNOZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_9_2 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_8_9_2  (
            .in0(N__6751),
            .in1(N__7228),
            .in2(_gnd_net_),
            .in3(N__5784),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_442_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_8_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_8_9_3 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_8_9_3  (
            .in0(N__8007),
            .in1(N__5103),
            .in2(N__4678),
            .in3(N__7144),
            .lcout(WRITE_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8792),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_8_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_8_9_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_8_9_6  (
            .in0(N__5834),
            .in1(N__5431),
            .in2(N__6761),
            .in3(N__5158),
            .lcout(),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_8_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_1_LC_8_9_7 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_1_LC_8_9_7  (
            .in0(N__4642),
            .in1(N__4675),
            .in2(N__4669),
            .in3(N__9274),
            .lcout(\U712_CHIP_RAM.BANK0_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__7533),
            .in2(_gnd_net_),
            .in3(N__6105),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_8_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_RNO_2_LC_8_12_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_CHIP_RAM.BANK0_RNO_2_LC_8_12_5  (
            .in0(N__4660),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10613),
            .lcout(\U712_CHIP_RAM.BANK0_RNOZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_5_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_5_0  (
            .in0(N__5836),
            .in1(N__5163),
            .in2(N__5445),
            .in3(N__6738),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8773),
            .ce(N__5797),
            .sr(N__10251));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_9_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_9_6_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIHQ8R_LC_9_6_0  (
            .in0(N__8028),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4704),
            .lcout(\U712_CHIP_RAM.N_605 ),
            .ltout(\U712_CHIP_RAM.N_605_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_9_6_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_9_6_1  (
            .in0(N__5963),
            .in1(N__4820),
            .in2(N__4633),
            .in3(N__6088),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKCP34_LC_9_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKCP34_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKCP34_LC_9_6_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKCP34_LC_9_6_2  (
            .in0(N__4629),
            .in1(N__5140),
            .in2(_gnd_net_),
            .in3(N__5404),
            .lcout(\U712_CHIP_RAM.N_700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_9_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_9_6_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_9_6_3  (
            .in0(N__5964),
            .in1(N__8029),
            .in2(N__5005),
            .in3(N__7796),
            .lcout(\U712_CHIP_RAM.N_697 ),
            .ltout(\U712_CHIP_RAM.N_697_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_6_4 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_6_4  (
            .in0(N__6089),
            .in1(_gnd_net_),
            .in2(N__4741),
            .in3(N__7160),
            .lcout(\U712_CHIP_RAM.N_537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNIHJRU1_LC_9_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNIHJRU1_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNIHJRU1_LC_9_6_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNIHJRU1_LC_9_6_5  (
            .in0(N__5302),
            .in1(N__8027),
            .in2(N__5205),
            .in3(N__6737),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_9_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_9_6_6 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_9_6_6  (
            .in0(N__5467),
            .in1(N__6654),
            .in2(N__4729),
            .in3(N__5346),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_9_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_9_6_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_9_6_7  (
            .in0(N__5962),
            .in1(N__4819),
            .in2(N__5004),
            .in3(N__7795),
            .lcout(\U712_CHIP_RAM.N_539 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_9_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_9_7_0 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_9_7_0  (
            .in0(N__4726),
            .in1(N__5926),
            .in2(N__5665),
            .in3(N__5295),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_9_7_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4720),
            .in3(N__10278),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_9_7_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_9_7_2  (
            .in0(N__5139),
            .in1(N__4703),
            .in2(_gnd_net_),
            .in3(N__5403),
            .lcout(\U712_CHIP_RAM.N_595 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_9_7_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_9_7_3  (
            .in0(N__5646),
            .in1(N__5198),
            .in2(_gnd_net_),
            .in3(N__5541),
            .lcout(\U712_CHIP_RAM.N_600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_1_LC_9_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_1_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_1_LC_9_7_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_1_LC_9_7_4  (
            .in0(N__4809),
            .in1(N__7790),
            .in2(_gnd_net_),
            .in3(N__4973),
            .lcout(\U712_CHIP_RAM.N_703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_7_5 .LUT_INIT=16'b1100000011010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_7_5  (
            .in0(N__5038),
            .in1(N__6145),
            .in2(N__8352),
            .in3(N__5026),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8779),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_1_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_1_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_1_LC_9_7_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_1_LC_9_7_6  (
            .in0(N__4810),
            .in1(N__7791),
            .in2(N__6086),
            .in3(N__4974),
            .lcout(\U712_CHIP_RAM.N_699 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_9_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_9_7_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_9_7_7  (
            .in0(N__5925),
            .in1(N__6048),
            .in2(N__7803),
            .in3(N__4808),
            .lcout(\U712_CHIP_RAM.N_589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_0 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_0  (
            .in0(N__4942),
            .in1(N__4930),
            .in2(N__4921),
            .in3(N__4895),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8784),
            .ce(N__4867),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_9_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_9_8_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_9_8_1  (
            .in0(N__9770),
            .in1(N__5927),
            .in2(_gnd_net_),
            .in3(N__6052),
            .lcout(\U712_CHIP_RAM.N_587 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_2  (
            .in0(N__7987),
            .in1(N__4906),
            .in2(N__5104),
            .in3(N__4896),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8784),
            .ce(N__4867),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_9_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__5706),
            .in2(_gnd_net_),
            .in3(N__6218),
            .lcout(),
            .ltout(\U712_REG_SM.N_513_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_9_2 .LUT_INIT=16'b1100000011000100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_9_9_2  (
            .in0(N__4846),
            .in1(N__7986),
            .in2(N__4828),
            .in3(N__5565),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8790),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_9_9_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_9_9_4  (
            .in0(N__9579),
            .in1(N__4825),
            .in2(_gnd_net_),
            .in3(N__6061),
            .lcout(\U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_5  (
            .in0(N__5162),
            .in1(N__5449),
            .in2(_gnd_net_),
            .in3(N__9967),
            .lcout(\U712_CHIP_RAM.DBENn_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIPCS25_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIPCS25_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIPCS25_LC_9_9_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIPCS25_LC_9_9_7  (
            .in0(N__6752),
            .in1(N__5835),
            .in2(_gnd_net_),
            .in3(N__6665),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI347S_1_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI347S_1_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI347S_1_LC_9_10_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI347S_1_LC_9_10_2  (
            .in0(N__6578),
            .in1(N__6512),
            .in2(_gnd_net_),
            .in3(N__5650),
            .lcout(\U712_REG_SM.N_694 ),
            .ltout(\U712_REG_SM.N_694_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_10_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5089),
            .in3(N__6259),
            .lcout(),
            .ltout(\U712_REG_SM.N_522_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_10_4 .LUT_INIT=16'b1110110011100100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_9_10_4  (
            .in0(N__7985),
            .in1(N__10106),
            .in2(N__5086),
            .in3(N__6928),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8793),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_10_6 .LUT_INIT=16'b1110010011101100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_10_6  (
            .in0(N__7984),
            .in1(N__6736),
            .in2(N__5275),
            .in3(N__9774),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8793),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_11_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_11_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_9_11_2  (
            .in0(N__5064),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8795),
            .ce(),
            .sr(N__10215));
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_11_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5044),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8795),
            .ce(),
            .sr(N__10215));
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_11_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5224),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8795),
            .ce(),
            .sr(N__10215));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_12_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__5263),
            .in2(_gnd_net_),
            .in3(N__6417),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_4  (
            .in0(N__6418),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7975),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8798),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_13_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_13_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_9_13_6  (
            .in0(N__5256),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8799),
            .ce(),
            .sr(N__10213));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_5_0 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_5_0  (
            .in0(N__6342),
            .in1(N__6357),
            .in2(N__6313),
            .in3(N__6372),
            .lcout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_5_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_5_1  (
            .in0(N__6876),
            .in1(N__6894),
            .in2(_gnd_net_),
            .in3(N__6909),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_10_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_10_5_2 .LUT_INIT=16'b0000110010001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_10_5_2  (
            .in0(N__6327),
            .in1(N__8024),
            .in2(N__5215),
            .in3(N__5212),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8766),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_10_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_10_5_5 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_10_5_5  (
            .in0(N__5545),
            .in1(N__9578),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.N_527 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_6 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_5_6  (
            .in0(N__9577),
            .in1(N__5176),
            .in2(N__9301),
            .in3(N__9068),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_6_0 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_10_6_0  (
            .in0(N__7301),
            .in1(N__6594),
            .in2(_gnd_net_),
            .in3(N__6535),
            .lcout(\U712_REG_SM.N_514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_10_6_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_10_6_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_10_6_1  (
            .in0(_gnd_net_),
            .in1(N__6240),
            .in2(_gnd_net_),
            .in3(N__6274),
            .lcout(\U712_REG_SM.N_422 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_10_6_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_10_6_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(N__6595),
            .in2(_gnd_net_),
            .in3(N__6536),
            .lcout(),
            .ltout(\U712_REG_SM.N_429_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_10_6_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_10_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_10_6_3 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_10_6_3  (
            .in0(N__8022),
            .in1(N__6199),
            .in2(N__5497),
            .in3(N__6275),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8774),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_6_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_6_4 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_6_4  (
            .in0(N__6241),
            .in1(N__6596),
            .in2(_gnd_net_),
            .in3(N__6537),
            .lcout(),
            .ltout(\U712_REG_SM.N_511_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_6_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_6_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_10_6_5  (
            .in0(N__8023),
            .in1(N__7037),
            .in2(N__5494),
            .in3(N__5491),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8774),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_6 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_1_LC_10_6_6  (
            .in0(N__9739),
            .in1(N__5968),
            .in2(_gnd_net_),
            .in3(N__5296),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_7 .LUT_INIT=16'b1010101011101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_7  (
            .in0(N__5466),
            .in1(N__5455),
            .in2(N__5447),
            .in3(N__5353),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_10_7_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_10_7_1  (
            .in0(N__5540),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5644),
            .lcout(\U712_CHIP_RAM.N_405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_10_7_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_10_7_2  (
            .in0(N__9757),
            .in1(N__5942),
            .in2(_gnd_net_),
            .in3(N__5294),
            .lcout(\U712_CHIP_RAM.N_597 ),
            .ltout(\U712_CHIP_RAM.N_597_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_7_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_7_3  (
            .in0(N__6762),
            .in1(N__6661),
            .in2(N__5278),
            .in3(N__5664),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_10_7_4 .LUT_INIT=16'b0000100010101000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_10_7_4  (
            .in0(N__7999),
            .in1(N__5676),
            .in2(N__5695),
            .in3(N__7729),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8776),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_10_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_10_7_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIOBA64_LC_10_7_5  (
            .in0(N__5941),
            .in1(N__7167),
            .in2(N__6087),
            .in3(N__5850),
            .lcout(\U712_CHIP_RAM.N_528 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_10_7_6 .LUT_INIT=16'b0100110001111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_10_7_6  (
            .in0(N__5645),
            .in1(N__6252),
            .in2(N__6601),
            .in3(N__7314),
            .lcout(),
            .ltout(\U712_REG_SM.N_482_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_10_7_7 .LUT_INIT=16'b0000101100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_10_7_7  (
            .in0(N__6538),
            .in1(N__6600),
            .in2(N__5620),
            .in3(N__8000),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8776),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_8_0 .LUT_INIT=16'b1100000011000100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_8_0  (
            .in0(N__5617),
            .in1(N__7990),
            .in2(N__5584),
            .in3(N__5572),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8780),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_8_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_8_1  (
            .in0(N__6740),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6652),
            .lcout(\U712_CHIP_RAM.BANK0_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.BANK0_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFS4TD_2_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFS4TD_2_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIFS4TD_2_LC_10_8_2 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIFS4TD_2_LC_10_8_2  (
            .in0(N__5952),
            .in1(N__5524),
            .in2(N__5509),
            .in3(N__5506),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_8_3 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_8_3  (
            .in0(N__10276),
            .in1(_gnd_net_),
            .in2(N__5500),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_4 .LUT_INIT=16'b1100000011010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_8_4  (
            .in0(N__6160),
            .in1(N__6146),
            .in2(N__8295),
            .in3(N__6118),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8780),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_8_5 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_8_5  (
            .in0(N__7168),
            .in1(N__6082),
            .in2(N__5977),
            .in3(N__5851),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_530_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_8_6 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_8_6  (
            .in0(N__6651),
            .in1(N__6739),
            .in2(N__5839),
            .in3(N__5829),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_8_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_10_8_7  (
            .in0(N__10275),
            .in1(_gnd_net_),
            .in2(N__5800),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_9_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_10_9_0 .LUT_INIT=16'b1111111110001010;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_10_9_0  (
            .in0(N__7642),
            .in1(N__8184),
            .in2(N__7357),
            .in3(N__7372),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8785),
            .ce(),
            .sr(N__10217));
    defparam \U712_CHIP_RAM.DBDIR_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_10_9_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_10_9_1 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_10_9_1  (
            .in0(N__5730),
            .in1(N__5785),
            .in2(_gnd_net_),
            .in3(N__5749),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8785),
            .ce(),
            .sr(N__10217));
    defparam \U712_CHIP_RAM.DBENn_LC_10_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_10_9_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_10_9_2 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_10_9_2  (
            .in0(N__9808),
            .in1(N__5719),
            .in2(_gnd_net_),
            .in3(N__5713),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8785),
            .ce(),
            .sr(N__10217));
    defparam \U712_REG_SM.START_RST_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_10_9_3 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.START_RST_LC_10_9_3  (
            .in0(N__5707),
            .in1(N__6195),
            .in2(_gnd_net_),
            .in3(N__6289),
            .lcout(\U712_REG_SM.START_RSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8785),
            .ce(),
            .sr(N__10217));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_10_9_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_10_9_4 .LUT_INIT=16'b0000101000001011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_10_9_4  (
            .in0(N__6295),
            .in1(N__7320),
            .in2(N__7042),
            .in3(N__7332),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8785),
            .ce(),
            .sr(N__10217));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_10_10_0 .LUT_INIT=16'b1101110101000100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_10_10_0  (
            .in0(N__6508),
            .in1(N__7266),
            .in2(_gnd_net_),
            .in3(N__6579),
            .lcout(\U712_REG_SM.N_407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_10_10_1 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_10_10_1  (
            .in0(N__7265),
            .in1(N__7237),
            .in2(_gnd_net_),
            .in3(N__6253),
            .lcout(\U712_REG_SM.DS_EN_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_RNO_0_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_RNO_0_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_RNO_0_LC_10_10_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \U712_REG_SM.ASn_RNO_0_LC_10_10_2  (
            .in0(N__6507),
            .in1(_gnd_net_),
            .in2(N__7273),
            .in3(N__6287),
            .lcout(\U712_REG_SM.N_443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_10_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_10_3  (
            .in0(N__6220),
            .in1(N__7268),
            .in2(_gnd_net_),
            .in3(N__7315),
            .lcout(\U712_REG_SM.STATE_COUNT_srsts_i_i_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_10_10_4 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_10_10_4  (
            .in0(N__6254),
            .in1(N__7267),
            .in2(N__6529),
            .in3(N__6288),
            .lcout(\U712_REG_SM.N_515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_10_10_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_2_LC_10_10_5 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_2_LC_10_10_5  (
            .in0(N__6286),
            .in1(N__6577),
            .in2(N__6530),
            .in3(N__6255),
            .lcout(\U712_REG_SM.un1_STATE_COUNT_4_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_10_10_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_10_10_6  (
            .in0(N__6506),
            .in1(N__6219),
            .in2(N__6593),
            .in3(N__6205),
            .lcout(\U712_REG_SM.START_RST_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_10_7 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_10_7  (
            .in0(N__7264),
            .in1(N__6573),
            .in2(_gnd_net_),
            .in3(N__6505),
            .lcout(\U712_REG_SM.N_480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_10_11_2 .LUT_INIT=16'b1111101100000001;
    LogicCell40 \U712_REG_SM.DS_EN_LC_10_11_2  (
            .in0(N__6184),
            .in1(N__6178),
            .in2(N__6172),
            .in3(N__9324),
            .lcout(DS_ENm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8794),
            .ce(),
            .sr(N__10214));
    defparam \U712_REG_SM.ASn_LC_10_11_7 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_LC_10_11_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_LC_10_11_7 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \U712_REG_SM.ASn_LC_10_11_7  (
            .in0(N__6607),
            .in1(N__6580),
            .in2(N__6534),
            .in3(N__6431),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8794),
            .ce(),
            .sr(N__10214));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_12_6 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_10_12_6  (
            .in0(N__11245),
            .in1(N__11324),
            .in2(_gnd_net_),
            .in3(N__7950),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8796),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_10_15_0.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_10_15_0.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_10_15_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_10_15_0 (
            .in0(N__7959),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DMA_LATCH_EN_i_i_a2_LC_10_19_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.DMA_LATCH_EN_i_i_a2_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DMA_LATCH_EN_i_i_a2_LC_10_19_0 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \U712_BUFFERS.DMA_LATCH_EN_i_i_a2_LC_10_19_0  (
            .in0(N__7179),
            .in1(N__11329),
            .in2(_gnd_net_),
            .in3(N__11256),
            .lcout(N_549),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_5_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_5_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_11_5_0  (
            .in0(_gnd_net_),
            .in1(N__6373),
            .in2(_gnd_net_),
            .in3(N__6361),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__6864),
            .ce(),
            .sr(N__6778));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_5_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_5_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__6358),
            .in2(_gnd_net_),
            .in3(N__6346),
            .lcout(\U712_CHIP_RAM.REFRESH5lto1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__6864),
            .ce(),
            .sr(N__6778));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_5_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_5_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(N__6343),
            .in2(_gnd_net_),
            .in3(N__6331),
            .lcout(\U712_CHIP_RAM.REFRESH5lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__6864),
            .ce(),
            .sr(N__6778));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_5_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_5_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__6328),
            .in2(_gnd_net_),
            .in3(N__6316),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__6864),
            .ce(),
            .sr(N__6778));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_5_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_5_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_11_5_4  (
            .in0(_gnd_net_),
            .in1(N__6312),
            .in2(_gnd_net_),
            .in3(N__6298),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__6864),
            .ce(),
            .sr(N__6778));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_5_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_5_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_11_5_5  (
            .in0(_gnd_net_),
            .in1(N__6910),
            .in2(_gnd_net_),
            .in3(N__6898),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__6864),
            .ce(),
            .sr(N__6778));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_5_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_5_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_11_5_6  (
            .in0(_gnd_net_),
            .in1(N__6895),
            .in2(_gnd_net_),
            .in3(N__6883),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__6864),
            .ce(),
            .sr(N__6778));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_5_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_5_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(N__6877),
            .in2(_gnd_net_),
            .in3(N__6880),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6864),
            .ce(),
            .sr(N__6778));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_6_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_11_6_2  (
            .in0(N__9005),
            .in1(N__6835),
            .in2(_gnd_net_),
            .in3(N__6813),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_6_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_11_6_3  (
            .in0(N__9147),
            .in1(N__9003),
            .in2(N__8296),
            .in3(N__8353),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(\U712_CHIP_RAM.REFRESH_RST_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_6_4 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_11_6_4  (
            .in0(N__9004),
            .in1(N__8354),
            .in2(N__6766),
            .in3(N__9148),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__6763),
            .in2(_gnd_net_),
            .in3(N__6669),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8775),
            .ce(N__6613),
            .sr(N__10222));
    defparam \U712_CYCLE_TERM.RAM_CYCLE_RNO_0_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.RAM_CYCLE_RNO_0_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.RAM_CYCLE_RNO_0_LC_11_8_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.RAM_CYCLE_RNO_0_LC_11_8_1  (
            .in0(N__6977),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6946),
            .lcout(\U712_CYCLE_TERM.N_566 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_8_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_8_2 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_8_2  (
            .in0(N__6947),
            .in1(N__6998),
            .in2(_gnd_net_),
            .in3(N__6978),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.TACK_EN_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_11_8_3 .LUT_INIT=16'b1100111100001111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__7585),
            .in2(N__7048),
            .in3(N__8038),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8777),
            .ce(),
            .sr(N__10218));
    defparam \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_0_a2_1_0_LC_11_8_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_0_a2_1_0_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_0_a2_1_0_LC_11_8_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_0_a2_1_0_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__6997),
            .in2(_gnd_net_),
            .in3(N__6976),
            .lcout(\U712_CYCLE_TERM.N_598 ),
            .ltout(\U712_CYCLE_TERM.N_598_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_8_5 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_11_8_5 .LUT_INIT=16'b0010001000110010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_11_8_5  (
            .in0(N__8089),
            .in1(N__8069),
            .in2(N__7045),
            .in3(N__8050),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8777),
            .ce(),
            .sr(N__10218));
    defparam \U712_REG_SM.REG_TACK_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_11_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_11_8_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_11_8_7  (
            .in0(N__7041),
            .in1(N__7015),
            .in2(N__7003),
            .in3(N__6916),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8777),
            .ce(),
            .sr(N__10218));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_9_0 .LUT_INIT=16'b0000000100110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_9_0  (
            .in0(N__7002),
            .in1(N__7349),
            .in2(N__6982),
            .in3(N__6948),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_571_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_9_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_9_1 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_11_9_1  (
            .in0(N__6949),
            .in1(N__7960),
            .in2(N__6931),
            .in3(N__8185),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8781),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_11_9_2  (
            .in0(N__7963),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7371),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8781),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_11_9_3 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_11_9_3  (
            .in0(N__7316),
            .in1(N__7236),
            .in2(_gnd_net_),
            .in3(N__6927),
            .lcout(\U712_REG_SM.REG_TACK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_9_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_11_9_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_11_9_4  (
            .in0(N__7961),
            .in1(N__8183),
            .in2(_gnd_net_),
            .in3(N__7350),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8781),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_11_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__7962),
            .in2(_gnd_net_),
            .in3(N__8070),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8781),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNI05SV_3_LC_11_9_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNI05SV_3_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNI05SV_3_LC_11_9_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNI05SV_3_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__7370),
            .in2(_gnd_net_),
            .in3(N__7348),
            .lcout(\U712_CYCLE_TERM.N_440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_10_2 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_11_10_2  (
            .in0(N__7949),
            .in1(N__7333),
            .in2(N__7321),
            .in3(N__7272),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8786),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_11_19_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_11_19_1 .LUT_INIT=16'b0000100001111111;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_11_19_1  (
            .in0(N__11325),
            .in1(N__11255),
            .in2(N__7235),
            .in3(N__7180),
            .lcout(N_483),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_3_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_3_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_3_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_12_3_0  (
            .in0(N__8888),
            .in1(N__8364),
            .in2(_gnd_net_),
            .in3(N__9073),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8759),
            .ce(N__8667),
            .sr(N__10243));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_4_0 .LUT_INIT=16'b1011001110000011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_4_0  (
            .in0(N__7675),
            .in1(N__9072),
            .in2(N__8893),
            .in3(N__7492),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8761),
            .ce(N__8677),
            .sr(N__10235));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_12_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_12_5_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(N__10277),
            .in2(_gnd_net_),
            .in3(N__7054),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_1 .LUT_INIT=16'b1100111110001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_12_5_1  (
            .in0(N__10039),
            .in1(N__8867),
            .in2(N__9086),
            .in3(N__9644),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_5_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(N__9160),
            .in2(_gnd_net_),
            .in3(N__8298),
            .lcout(\U712_CHIP_RAM.N_412 ),
            .ltout(\U712_CHIP_RAM.N_412_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_4 .LUT_INIT=16'b0010010100000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_5_4  (
            .in0(N__9075),
            .in1(N__9620),
            .in2(N__7516),
            .in3(N__10038),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_5_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_5_5  (
            .in0(N__9621),
            .in1(N__7513),
            .in2(_gnd_net_),
            .in3(N__9421),
            .lcout(\U712_CHIP_RAM.N_478 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_6  (
            .in0(N__9076),
            .in1(N__7486),
            .in2(N__9663),
            .in3(N__8428),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_5_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(N__9643),
            .in2(_gnd_net_),
            .in3(N__9074),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_1 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_6_1  (
            .in0(N__7474),
            .in1(N__9021),
            .in2(N__9659),
            .in3(N__9472),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_6_2 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_12_6_2  (
            .in0(N__8874),
            .in1(N__8927),
            .in2(N__7468),
            .in3(N__9880),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8763),
            .ce(N__8676),
            .sr(N__10221));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_6_6 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_12_6_6  (
            .in0(N__8875),
            .in1(N__8928),
            .in2(N__8419),
            .in3(N__8191),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8763),
            .ce(N__8676),
            .sr(N__10221));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_12_7_2  (
            .in0(N__7435),
            .in1(N__7401),
            .in2(_gnd_net_),
            .in3(N__9070),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_3  (
            .in0(N__9071),
            .in1(N__9636),
            .in2(N__8194),
            .in3(N__8443),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pll_RNI8MQ3_LC_12_8_0.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_12_8_0.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_12_8_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 pll_RNI8MQ3_LC_12_8_0 (
            .in0(N__8182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNIDG0M2_4_LC_12_8_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNIDG0M2_4_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNIDG0M2_4_LC_12_8_1 .LUT_INIT=16'b1111010111110100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNIDG0M2_4_LC_12_8_1  (
            .in0(N__8088),
            .in1(N__8077),
            .in2(N__8071),
            .in3(N__8049),
            .lcout(\U712_CYCLE_TERM.un13_0 ),
            .ltout(\U712_CYCLE_TERM.un13_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.RAM_CYCLE_LC_12_8_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.RAM_CYCLE_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.RAM_CYCLE_LC_12_8_2 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \U712_CYCLE_TERM.RAM_CYCLE_LC_12_8_2  (
            .in0(N__7924),
            .in1(N__7828),
            .in2(N__7822),
            .in3(N__7620),
            .lcout(\U712_CYCLE_TERM.RAM_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8769),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_8_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_8_4  (
            .in0(N__9635),
            .in1(N__9069),
            .in2(N__7819),
            .in3(N__9367),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_12_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_12_8_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_12_8_6  (
            .in0(_gnd_net_),
            .in1(N__9738),
            .in2(_gnd_net_),
            .in3(N__7807),
            .lcout(\U712_CHIP_RAM.N_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_8_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_8_7  (
            .in0(N__7710),
            .in1(N__9634),
            .in2(_gnd_net_),
            .in3(N__9976),
            .lcout(\U712_CHIP_RAM.N_455 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.RAM_CYCLE_RNILITE_LC_12_9_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.RAM_CYCLE_RNILITE_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.RAM_CYCLE_RNILITE_LC_12_9_3 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \U712_CYCLE_TERM.RAM_CYCLE_RNILITE_LC_12_9_3  (
            .in0(N__7652),
            .in1(N__7621),
            .in2(_gnd_net_),
            .in3(N__7586),
            .lcout(U712_CYCLE_TERM_TCIn_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_11_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_11_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_11_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_12_13_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_12_13_3 .LUT_INIT=16'b1011000000110000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_LC_12_13_3  (
            .in0(N__11005),
            .in1(N__11158),
            .in2(N__9667),
            .in3(N__9228),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_563_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_56_i_LC_12_13_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_56_i_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_56_i_LC_12_13_4 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \U712_BYTE_ENABLE.N_56_i_LC_12_13_4  (
            .in0(N__9781),
            .in1(N__9834),
            .in2(N__8407),
            .in3(N__11320),
            .lcout(N_56_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_o2_LC_12_15_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_o2_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_o2_LC_12_15_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_0_0_o2_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__11053),
            .in2(_gnd_net_),
            .in3(N__10869),
            .lcout(\U712_BYTE_ENABLE.N_410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WEn_LC_13_2_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_13_2_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_13_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_13_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8302),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8760),
            .ce(),
            .sr(N__10257));
    defparam \U712_CHIP_RAM.CRCSn_LC_13_2_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_2_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_13_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8365),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8760),
            .ce(),
            .sr(N__10257));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_4_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_4_0 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_4_0  (
            .in0(N__9168),
            .in1(N__9050),
            .in2(_gnd_net_),
            .in3(N__8297),
            .lcout(\U712_CHIP_RAM.CMA_5_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_4_5 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_13_4_5  (
            .in0(N__9051),
            .in1(N__8245),
            .in2(N__9664),
            .in3(N__8437),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_5_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_13_5_0  (
            .in0(N__8236),
            .in1(N__8230),
            .in2(_gnd_net_),
            .in3(N__8224),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8764),
            .ce(N__8675),
            .sr(N__10237));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_5_2 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_13_5_2  (
            .in0(N__8921),
            .in1(N__10684),
            .in2(N__8890),
            .in3(N__8617),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8764),
            .ce(N__8675),
            .sr(N__10237));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_5_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_13_5_3  (
            .in0(N__8523),
            .in1(N__8590),
            .in2(N__9658),
            .in3(N__10630),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8764),
            .ce(N__8675),
            .sr(N__10237));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_13_5_6 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_13_5_6  (
            .in0(N__8922),
            .in1(N__9478),
            .in2(N__8891),
            .in3(N__8548),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8764),
            .ce(N__8675),
            .sr(N__10237));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_6_4 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_13_6_4  (
            .in0(N__8527),
            .in1(N__8512),
            .in2(N__9665),
            .in3(N__10372),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8767),
            .ce(N__8674),
            .sr(N__10232));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_6_6 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_13_6_6  (
            .in0(N__8926),
            .in1(N__9484),
            .in2(N__8892),
            .in3(N__8473),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8767),
            .ce(N__8674),
            .sr(N__10232));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_7_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_7_1  (
            .in0(N__9460),
            .in1(N__9407),
            .in2(_gnd_net_),
            .in3(N__10594),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__10316),
            .sr(N__10223));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_7_2  (
            .in0(N__10596),
            .in1(N__10428),
            .in2(_gnd_net_),
            .in3(N__10675),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__10316),
            .sr(N__10223));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_4  (
            .in0(N__10595),
            .in1(N__10731),
            .in2(_gnd_net_),
            .in3(N__10674),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__10316),
            .sr(N__10223));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_8_5  (
            .in0(N__10587),
            .in1(N__9456),
            .in2(_gnd_net_),
            .in3(N__10018),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10355),
            .ce(N__10314),
            .sr(N__10219));
    defparam \U712_CHIP_RAM.DMA_A20_LC_13_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_13_9_5 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_13_9_5  (
            .in0(N__9289),
            .in1(N__10421),
            .in2(N__10591),
            .in3(N__9270),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__10216));
    defparam \U712_BYTE_ENABLE.N_58_i_LC_13_12_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_58_i_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_58_i_LC_13_12_1 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \U712_BYTE_ENABLE.N_58_i_LC_13_12_1  (
            .in0(N__9835),
            .in1(N__11316),
            .in2(N__9211),
            .in3(N__9783),
            .lcout(N_58_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_13_13_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_13_13_1 .LUT_INIT=16'b0111001100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_13_13_1  (
            .in0(N__11018),
            .in1(N__11157),
            .in2(N__9232),
            .in3(N__9666),
            .lcout(\U712_BYTE_ENABLE.N_559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_129_i_LC_13_20_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_129_i_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_129_i_LC_13_20_2 .LUT_INIT=16'b0000111011100000;
    LogicCell40 \U712_BYTE_ENABLE.N_129_i_LC_13_20_2  (
            .in0(N__11006),
            .in1(N__11065),
            .in2(N__10927),
            .in3(N__10841),
            .lcout(N_129_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_14_2_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_14_2_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_14_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_14_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9088),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8762),
            .ce(),
            .sr(N__10260));
    defparam \U712_CHIP_RAM.RASn_LC_14_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_14_4_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_14_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_14_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9169),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8765),
            .ce(),
            .sr(N__10252));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_5_1 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_5_1  (
            .in0(N__9648),
            .in1(N__9100),
            .in2(N__9087),
            .in3(N__10090),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_14_5_2 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_14_5_2  (
            .in0(N__8929),
            .in1(N__8889),
            .in2(N__8827),
            .in3(N__9490),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__8768),
            .ce(N__8663),
            .sr(N__10245));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_6_0  (
            .in0(N__10617),
            .in1(N__9409),
            .in2(_gnd_net_),
            .in3(N__10068),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10357),
            .ce(N__10321),
            .sr(N__10238));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_6_3  (
            .in0(N__9408),
            .in1(N__9455),
            .in2(_gnd_net_),
            .in3(N__10616),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10357),
            .ce(N__10321),
            .sr(N__10238));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_6_7  (
            .in0(N__10673),
            .in1(N__10735),
            .in2(_gnd_net_),
            .in3(N__10618),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10357),
            .ce(N__10321),
            .sr(N__10238));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_7_4  (
            .in0(N__9955),
            .in1(N__10020),
            .in2(_gnd_net_),
            .in3(N__10530),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10319),
            .sr(N__10233));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_7_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_7_7  (
            .in0(N__10531),
            .in1(_gnd_net_),
            .in2(N__10024),
            .in3(N__9448),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10319),
            .sr(N__10233));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_8_6  (
            .in0(N__10067),
            .in1(N__9398),
            .in2(_gnd_net_),
            .in3(N__10555),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__10317),
            .sr(N__10224));
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_14_20_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_14_20_4 .LUT_INIT=16'b0100100011111111;
    LogicCell40 \U712_BYTE_ENABLE.un1_UDSn_i_0_0_LC_14_20_4  (
            .in0(N__10843),
            .in1(N__11086),
            .in2(N__10929),
            .in3(N__9340),
            .lcout(un1_UDSn_i_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_14_20_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_14_20_6 .LUT_INIT=16'b0001000011111111;
    LogicCell40 \U712_BYTE_ENABLE.un1_LDSn_i_0_0_LC_14_20_6  (
            .in0(N__10842),
            .in1(N__11085),
            .in2(N__10928),
            .in3(N__9339),
            .lcout(un1_LDSn_i_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_5_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_5_2  (
            .in0(N__10615),
            .in1(N__10786),
            .in2(_gnd_net_),
            .in3(N__10730),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__10324),
            .sr(N__10253));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_15_6_0  (
            .in0(N__10614),
            .in1(N__10084),
            .in2(_gnd_net_),
            .in3(N__10778),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__10323),
            .sr(N__10246));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_7_2  (
            .in0(N__10521),
            .in1(N__10080),
            .in2(_gnd_net_),
            .in3(N__10769),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10353),
            .ce(N__10322),
            .sr(N__10239));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_6  (
            .in0(N__10019),
            .in1(N__9954),
            .in2(_gnd_net_),
            .in3(N__10599),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10352),
            .ce(N__10320),
            .sr(N__10234));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_5  (
            .in0(N__10598),
            .in1(N__9913),
            .in2(_gnd_net_),
            .in3(N__9946),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10318),
            .sr(N__10225));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_10_5  (
            .in0(N__9953),
            .in1(N__9909),
            .in2(_gnd_net_),
            .in3(N__10597),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10351),
            .ce(N__10315),
            .sr(N__10220));
    defparam \U712_BYTE_ENABLE.N_57_i_LC_15_11_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_57_i_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_57_i_LC_15_11_1 .LUT_INIT=16'b0011001100100011;
    LogicCell40 \U712_BYTE_ENABLE.N_57_i_LC_15_11_1  (
            .in0(N__11224),
            .in1(N__11167),
            .in2(N__9787),
            .in3(N__9845),
            .lcout(N_57_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_59_i_LC_15_12_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_59_i_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_59_i_LC_15_12_7 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \U712_BYTE_ENABLE.N_59_i_LC_15_12_7  (
            .in0(N__11257),
            .in1(N__9673),
            .in2(N__9850),
            .in3(N__9782),
            .lcout(N_59_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_15_13_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_15_13_0 .LUT_INIT=16'b0001111100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_15_13_0  (
            .in0(N__11084),
            .in1(N__11020),
            .in2(N__11156),
            .in3(N__9629),
            .lcout(\U712_BYTE_ENABLE.N_557 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_15_13_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_15_13_4 .LUT_INIT=16'b0100111100000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_0_a2_LC_15_13_4  (
            .in0(N__11083),
            .in1(N__11019),
            .in2(N__11155),
            .in3(N__9628),
            .lcout(\U712_BYTE_ENABLE.N_561 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_0_x2_LC_15_16_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_0_x2_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_i_o2_0_x2_LC_15_16_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_i_o2_0_x2_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(N__10942),
            .in2(_gnd_net_),
            .in3(N__10870),
            .lcout(\U712_BYTE_ENABLE.N_397_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_130_i_LC_15_20_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_130_i_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_130_i_LC_15_20_0 .LUT_INIT=16'b0000110111010000;
    LogicCell40 \U712_BYTE_ENABLE.N_130_i_LC_15_20_0  (
            .in0(N__11012),
            .in1(N__11089),
            .in2(N__10868),
            .in3(N__10936),
            .lcout(N_130_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_127_i_LC_15_20_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_127_i_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_127_i_LC_15_20_1 .LUT_INIT=16'b0000110011010000;
    LogicCell40 \U712_BYTE_ENABLE.N_127_i_LC_15_20_1  (
            .in0(N__11087),
            .in1(N__11010),
            .in2(N__10940),
            .in3(N__10857),
            .lcout(N_127_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_128_i_LC_15_20_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_128_i_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_128_i_LC_15_20_5 .LUT_INIT=16'b0000001101110000;
    LogicCell40 \U712_BYTE_ENABLE.N_128_i_LC_15_20_5  (
            .in0(N__11088),
            .in1(N__11011),
            .in2(N__10941),
            .in3(N__10858),
            .lcout(N_128_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_5_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_16_5_2  (
            .in0(N__10593),
            .in1(N__10785),
            .in2(_gnd_net_),
            .in3(N__10720),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10356),
            .ce(N__10327),
            .sr(N__10258));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_6_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_6_1  (
            .in0(N__10592),
            .in1(N__10429),
            .in2(_gnd_net_),
            .in3(N__10667),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10354),
            .ce(N__10325),
            .sr(N__10254));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_18_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_18_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_18_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_18_8_5  (
            .in0(N__10569),
            .in1(N__10438),
            .in2(_gnd_net_),
            .in3(N__10403),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10350),
            .ce(N__10326),
            .sr(N__10255));
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_19_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_19_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_19_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_19_5  (
            .in0(N__10126),
            .in1(N__11300),
            .in2(_gnd_net_),
            .in3(N__11218),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

module U400_CYCLE_TERM (

    output TACKn

);

assign TACKn = 1'bz;

endmodule

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 13 2025 09:32:57

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U111_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U111_TOP
entity U111_TOP is
port (
    D_LM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UM_AMIGA : inout std_logic_vector(7 downto 0);
    D_LL_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_AMIGA : inout std_logic_vector(7 downto 0);
    D_LL_040 : inout std_logic_vector(7 downto 0);
    D_UU_040 : inout std_logic_vector(7 downto 0);
    D_LM_040 : inout std_logic_vector(7 downto 0);
    D_UM_040 : inout std_logic_vector(7 downto 0);
    A_AMIGA : out std_logic_vector(1 downto 0);
    A_040 : in std_logic_vector(1 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    TBIn : in std_logic;
    TEAn : in std_logic;
    TSn : inout std_logic;
    RESETn : in std_logic;
    CLKRAMA : out std_logic;
    PORTSIZE : in std_logic;
    DMAAn : out std_logic;
    TEA_CPUn : out std_logic;
    LBENn : in std_logic;
    CLK40B : out std_logic;
    TBI_CPUn : out std_logic;
    TAn : inout std_logic;
    CPUBGn : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CLK80_CPU : out std_logic;
    BUFDIR : out std_logic;
    TCI_CPUn : out std_logic;
    TS_CPUn : inout std_logic;
    CLKRAMB : out std_logic;
    CLK40A : out std_logic;
    TCIn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    BBn : in std_logic;
    TACKn : inout std_logic;
    BGn : in std_logic);
end U111_TOP;

-- Architecture of U111_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U111_TOP is

signal \N__9464\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4344\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3054\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2790\ : std_logic;
signal \N__2787\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2688\ : std_logic;
signal \N__2685\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2655\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2595\ : std_logic;
signal \TCIn_c\ : std_logic;
signal \TSn_in\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \TAn_in\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U111_CYCLE_SM_A_AMIGA_0_i_1\ : std_logic;
signal \A_040_c_0\ : std_logic;
signal \A_AMIGA_c_0\ : std_logic;
signal \D_LL_AMIGA_in_4\ : std_logic;
signal \un2_D_LL_AMIGA_4\ : std_logic;
signal \D_LL_AMIGA_in_1\ : std_logic;
signal \un2_D_LL_AMIGA_1\ : std_logic;
signal \D_UM_040_in_0\ : std_logic;
signal \D_LL_040_in_0\ : std_logic;
signal \un1_D_UM_040_0\ : std_logic;
signal \D_LM_AMIGA_in_3\ : std_logic;
signal \N_119\ : std_logic;
signal \D_LM_AMIGA_in_1\ : std_logic;
signal \N_121\ : std_logic;
signal \D_LL_040_in_6\ : std_logic;
signal \D_UM_040_in_6\ : std_logic;
signal \un1_D_UM_040_6\ : std_logic;
signal \D_LM_AMIGA_in_2\ : std_logic;
signal \N_120\ : std_logic;
signal \D_LM_040_in_0\ : std_logic;
signal \D_UU_040_in_0\ : std_logic;
signal \un1_D_UU_040_0\ : std_logic;
signal \D_UU_040_in_4\ : std_logic;
signal \D_LM_040_in_4\ : std_logic;
signal \un1_D_UU_040_4\ : std_logic;
signal \D_UU_040_in_6\ : std_logic;
signal \D_LM_040_in_6\ : std_logic;
signal \un1_D_UU_040_6\ : std_logic;
signal \D_LL_AMIGA_in_2\ : std_logic;
signal \un2_D_LL_AMIGA_2\ : std_logic;
signal \D_LL_AMIGA_in_3\ : std_logic;
signal \un2_D_LL_AMIGA_3\ : std_logic;
signal \A_040_c_1\ : std_logic;
signal \D_LM_AMIGA_in_0\ : std_logic;
signal \N_122\ : std_logic;
signal \U111_CYCLE_SM.A2_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.N_151\ : std_logic;
signal \D_UM_040_in_1\ : std_logic;
signal \D_LL_040_in_1\ : std_logic;
signal \un1_D_UM_040_1\ : std_logic;
signal \D_LL_040_in_3\ : std_logic;
signal \D_UM_040_in_3\ : std_logic;
signal \un1_D_UM_040_3\ : std_logic;
signal \D_LM_AMIGA_in_7\ : std_logic;
signal \N_115\ : std_logic;
signal \D_UU_AMIGA_in_2\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\ : std_logic;
signal \N_129\ : std_logic;
signal \D_UU_040_in_2\ : std_logic;
signal \D_LM_040_in_2\ : std_logic;
signal \un1_D_UU_040_2\ : std_logic;
signal \CPUBGn_c_i_0\ : std_logic;
signal \D_LL_AMIGA_in_7\ : std_logic;
signal \un2_D_LL_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.N_112_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_144_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_142\ : std_logic;
signal \U111_CYCLE_SM.N_197\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\ : std_logic;
signal \U111_CYCLE_SM.N_195_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_1_0\ : std_logic;
signal \TBIn_c\ : std_logic;
signal \U111_CYCLE_SM.BURSTZ0\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNTZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.BURST_COUNTZ0Z_1\ : std_logic;
signal \U111_CYCLE_SM.N_109\ : std_logic;
signal \U111_CYCLE_SM.N_109_cascade_\ : std_logic;
signal \U111_CYCLE_SM.PORT_MISMATCHZ0\ : std_logic;
signal \D_LM_AMIGA_in_5\ : std_logic;
signal \N_117\ : std_logic;
signal \D_LM_AMIGA_in_4\ : std_logic;
signal \N_118\ : std_logic;
signal \D_UM_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\ : std_logic;
signal \un1_D_UM_AMIGA_1\ : std_logic;
signal \D_LM_AMIGA_in_6\ : std_logic;
signal \N_116\ : std_logic;
signal \N_102_i\ : std_logic;
signal \BUFDIR_c\ : std_logic;
signal \BBn_c\ : std_logic;
signal \N_104\ : std_logic;
signal \D_UU_AMIGA_in_3\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\ : std_logic;
signal \N_128\ : std_logic;
signal \U111_CYCLE_SM.N_195\ : std_logic;
signal \U111_CYCLE_SM.N_132\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0\ : std_logic;
signal \TS_OUT\ : std_logic;
signal \INVU111_CYCLE_SM.TS_OUTC_net\ : std_logic;
signal \PORTSIZE_c\ : std_logic;
signal \U111_CYCLE_SM_OFFBOARD_EN_0\ : std_logic;
signal \U111_CYCLE_SM.un4_TS_OUT_i_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.N_106\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U111_CYCLE_SM.N_140\ : std_logic;
signal \U111_CYCLE_SM.N_107\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U111_CYCLE_SM.LATCH_EN_5\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\ : std_logic;
signal \U111_CYCLE_SM.N_57\ : std_logic;
signal \D_UM_AMIGA_in_7\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\ : std_logic;
signal \un1_D_UM_AMIGA_7\ : std_logic;
signal \GB_BUFFER_CLK40_THRU_CO\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\ : std_logic;
signal \D_UU_AMIGA_in_6\ : std_logic;
signal \N_124\ : std_logic;
signal \D_UU_AMIGA_in_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\ : std_logic;
signal \N_126\ : std_logic;
signal \D_UU_AMIGA_in_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\ : std_logic;
signal \N_123\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\ : std_logic;
signal \D_UU_AMIGA_in_4\ : std_logic;
signal \N_127\ : std_logic;
signal \TEAn_c\ : std_logic;
signal \U111_CYCLE_SM_TEA_CPUn_0_i\ : std_logic;
signal \D_UU_040_in_1\ : std_logic;
signal \D_LM_040_in_1\ : std_logic;
signal \un1_D_UU_040_1\ : std_logic;
signal \D_UM_040_in_7\ : std_logic;
signal \D_LL_040_in_7\ : std_logic;
signal \un1_D_UM_040_7\ : std_logic;
signal \D_UM_AMIGA_in_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\ : std_logic;
signal \un1_D_UM_AMIGA_3\ : std_logic;
signal \D_LL_040_in_4\ : std_logic;
signal \D_UM_040_in_4\ : std_logic;
signal \un1_D_UM_040_4\ : std_logic;
signal \D_LL_AMIGA_in_6\ : std_logic;
signal \un2_D_LL_AMIGA_6\ : std_logic;
signal \D_LL_AMIGA_in_5\ : std_logic;
signal \un2_D_LL_AMIGA_5\ : std_logic;
signal \TS_CPUn_in\ : std_logic;
signal \U111_CYCLE_SM.TS_DELAYZ0\ : std_logic;
signal \U111_CYCLE_SM.un4_TS_OUT_i_0\ : std_logic;
signal \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.N_107_i\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\ : std_logic;
signal \U111_CYCLE_SM.LW_TRANSZ0\ : std_logic;
signal \CLK40\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \D_UU_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\ : std_logic;
signal \N_130\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\ : std_logic;
signal \D_UU_AMIGA_in_0\ : std_logic;
signal \N_131\ : std_logic;
signal \U111_CYCLE_SM.TA_DISZ0\ : std_logic;
signal \N_66\ : std_logic;
signal \D_UM_AMIGA_in_5\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\ : std_logic;
signal \un1_D_UM_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\ : std_logic;
signal \D_UM_AMIGA_in_4\ : std_logic;
signal \un1_D_UM_AMIGA_4\ : std_logic;
signal \D_UU_040_in_5\ : std_logic;
signal \D_LM_040_in_5\ : std_logic;
signal \un1_D_UU_040_5\ : std_logic;
signal \LBENn_c\ : std_logic;
signal \LBENn_c_i\ : std_logic;
signal \D_LL_AMIGA_in_0\ : std_logic;
signal \un2_D_LL_AMIGA_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_ENZ0\ : std_logic;
signal \BGn_c\ : std_logic;
signal \CPUBGn_c\ : std_logic;
signal \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\ : std_logic;
signal \CPUBGn_c_cascade_\ : std_logic;
signal \RnW_c\ : std_logic;
signal \N_62_i\ : std_logic;
signal \D_UM_AMIGA_in_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\ : std_logic;
signal \un1_D_UM_AMIGA_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\ : std_logic;
signal \D_UM_AMIGA_in_0\ : std_logic;
signal \un1_D_UM_AMIGA_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\ : std_logic;
signal \D_UM_AMIGA_in_6\ : std_logic;
signal \U111_CYCLE_SM.LATCH_ENZ0\ : std_logic;
signal \N_125\ : std_logic;
signal \D_LL_040_in_2\ : std_logic;
signal \D_UM_040_in_2\ : std_logic;
signal \un1_D_UM_040_2\ : std_logic;
signal \CLK80\ : std_logic;
signal \GB_BUFFER_CLK80_THRU_CO\ : std_logic;
signal \D_UU_040_in_3\ : std_logic;
signal \D_LM_040_in_3\ : std_logic;
signal \un1_D_UU_040_3\ : std_logic;
signal \D_UU_040_in_7\ : std_logic;
signal \D_LM_040_in_7\ : std_logic;
signal \un1_D_UU_040_7\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \D_LL_040_in_5\ : std_logic;
signal \D_UM_040_in_5\ : std_logic;
signal \U111_CYCLE_SM.FLIP_WORDZ0\ : std_logic;
signal \un1_D_UM_040_5\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \LBENn_wire\ : std_logic;
signal \CPUBGn_wire\ : std_logic;
signal \TEA_CPUn_wire\ : std_logic;
signal \A_040_wire\ : std_logic_vector(1 downto 0);
signal \A_AMIGA_wire\ : std_logic_vector(1 downto 0);
signal \CLK40B_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \BUFDIR_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \CLKRAMB_wire\ : std_logic;
signal \TEAn_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \CLK80_CPU_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \BGn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \TBI_CPUn_wire\ : std_logic;
signal \CLK40A_wire\ : std_logic;
signal \CLKRAMA_wire\ : std_logic;
signal \TCI_CPUn_wire\ : std_logic;
signal \BBn_wire\ : std_logic;
signal \DMAAn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \pll_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \LBENn_wire\ <= LBENn;
    CPUBGn <= \CPUBGn_wire\;
    TEA_CPUn <= \TEA_CPUn_wire\;
    \A_040_wire\ <= A_040;
    A_AMIGA <= \A_AMIGA_wire\;
    CLK40B <= \CLK40B_wire\;
    \TBIn_wire\ <= TBIn;
    BUFDIR <= \BUFDIR_wire\;
    \SIZ_wire\ <= SIZ;
    CLKRAMB <= \CLKRAMB_wire\;
    \TEAn_wire\ <= TEAn;
    BUFENn <= \BUFENn_wire\;
    CLK80_CPU <= \CLK80_CPU_wire\;
    \PORTSIZE_wire\ <= PORTSIZE;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    \BGn_wire\ <= BGn;
    \TCIn_wire\ <= TCIn;
    TBI_CPUn <= \TBI_CPUn_wire\;
    CLK40A <= \CLK40A_wire\;
    CLKRAMA <= \CLKRAMA_wire\;
    TCI_CPUn <= \TCI_CPUn_wire\;
    \BBn_wire\ <= BBn;
    DMAAn <= \DMAAn_wire\;
    \RnW_wire\ <= RnW;
    \pll_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_pll\ : PLL40_2F
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            SCLK => '0',
            PLLOUTGLOBALA => \CLK80\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALB => \CLK40\,
            SDI => '0',
            PLLOUTCOREA => OPEN,
            BYPASS => '0',
            RESETB => \N__7998\,
            PLLOUTCOREB => OPEN,
            LOCK => OPEN,
            SDO => OPEN,
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \pll_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__9464\
        );

    \pll_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__9464\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \LBENn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9448\,
            DIN => \N__9447\,
            DOUT => \N__9446\,
            PACKAGEPIN => \LBENn_wire\
        );

    \LBENn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9448\,
            PADOUT => \N__9447\,
            PADIN => \N__9446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \LBENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9439\,
            DIN => \N__9438\,
            DOUT => \N__9437\,
            PACKAGEPIN => D_UM_040(3)
        );

    \D_UM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9439\,
            PADOUT => \N__9438\,
            PADIN => \N__9437\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7010\,
            DIN0 => \D_UM_040_in_3\,
            DOUT0 => \N__6015\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9430\,
            DIN => \N__9429\,
            DOUT => \N__9428\,
            PACKAGEPIN => TAn
        );

    \TAn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9430\,
            PADOUT => \N__9429\,
            PADIN => \N__9428\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6105\,
            DIN0 => \TAn_in\,
            DOUT0 => \N__4548\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9421\,
            DIN => \N__9420\,
            DOUT => \N__9419\,
            PACKAGEPIN => D_LL_AMIGA(1)
        );

    \D_LL_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9421\,
            PADOUT => \N__9420\,
            PADIN => \N__9419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4910\,
            DIN0 => \D_LL_AMIGA_in_1\,
            DOUT0 => \N__3341\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9412\,
            DIN => \N__9411\,
            DOUT => \N__9410\,
            PACKAGEPIN => D_UU_AMIGA(5)
        );

    \D_UU_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9412\,
            PADOUT => \N__9411\,
            PADIN => \N__9410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4931\,
            DIN0 => \D_UU_AMIGA_in_5\,
            DOUT0 => \N__7470\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9403\,
            DIN => \N__9402\,
            DOUT => \N__9401\,
            PACKAGEPIN => D_UU_040(6)
        );

    \D_UU_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9403\,
            PADOUT => \N__9402\,
            PADIN => \N__9401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6973\,
            DIN0 => \D_UU_040_in_6\,
            DOUT0 => \N__5649\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUBGn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9394\,
            DIN => \N__9393\,
            DOUT => \N__9392\,
            PACKAGEPIN => \CPUBGn_wire\
        );

    \CPUBGn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9394\,
            PADOUT => \N__9393\,
            PADIN => \N__9392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7272\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9385\,
            DIN => \N__9384\,
            DOUT => \N__9383\,
            PACKAGEPIN => D_LL_040(7)
        );

    \D_LL_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9385\,
            PADOUT => \N__9384\,
            PADIN => \N__9383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6850\,
            DIN0 => \D_LL_040_in_7\,
            DOUT0 => \N__3567\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9376\,
            DIN => \N__9375\,
            DOUT => \N__9374\,
            PACKAGEPIN => D_LL_AMIGA(4)
        );

    \D_LL_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9376\,
            PADOUT => \N__9375\,
            PADIN => \N__9374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4909\,
            DIN0 => \D_LL_AMIGA_in_4\,
            DOUT0 => \N__5999\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9367\,
            DIN => \N__9366\,
            DOUT => \N__9365\,
            PACKAGEPIN => D_UM_AMIGA(3)
        );

    \D_UM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9367\,
            PADOUT => \N__9366\,
            PADIN => \N__9365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4918\,
            DIN0 => \D_UM_AMIGA_in_3\,
            DOUT0 => \N__3816\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9358\,
            DIN => \N__9357\,
            DOUT => \N__9356\,
            PACKAGEPIN => D_UU_040(3)
        );

    \D_UU_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9358\,
            PADOUT => \N__9357\,
            PADIN => \N__9356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7004\,
            DIN0 => \D_UU_040_in_3\,
            DOUT0 => \N__4158\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEA_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9349\,
            DIN => \N__9348\,
            DOUT => \N__9347\,
            PACKAGEPIN => \TEA_CPUn_wire\
        );

    \TEA_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9349\,
            PADOUT => \N__9348\,
            PADIN => \N__9347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5310\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9340\,
            DIN => \N__9339\,
            DOUT => \N__9338\,
            PACKAGEPIN => \A_040_wire\(1)
        );

    \A_040_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9340\,
            PADOUT => \N__9339\,
            PADIN => \N__9338\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9331\,
            DIN => \N__9330\,
            DOUT => \N__9329\,
            PACKAGEPIN => D_LM_AMIGA(3)
        );

    \D_LM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9331\,
            PADOUT => \N__9330\,
            PADIN => \N__9329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4708\,
            DIN0 => \D_LM_AMIGA_in_3\,
            DOUT0 => \N__8139\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9322\,
            DIN => \N__9321\,
            DOUT => \N__9320\,
            PACKAGEPIN => D_LM_040(0)
        );

    \D_LM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9322\,
            PADOUT => \N__9321\,
            PADIN => \N__9320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6851\,
            DIN0 => \D_LM_040_in_0\,
            DOUT0 => \N__3429\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9313\,
            DIN => \N__9312\,
            DOUT => \N__9311\,
            PACKAGEPIN => D_UM_AMIGA(6)
        );

    \D_UM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9313\,
            PADOUT => \N__9312\,
            PADIN => \N__9311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4930\,
            DIN0 => \D_UM_AMIGA_in_6\,
            DOUT0 => \N__3069\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9304\,
            DIN => \N__9303\,
            DOUT => \N__9302\,
            PACKAGEPIN => D_LM_AMIGA(4)
        );

    \D_LM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9304\,
            PADOUT => \N__9303\,
            PADIN => \N__9302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4840\,
            DIN0 => \D_LM_AMIGA_in_4\,
            DOUT0 => \N__2925\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9295\,
            DIN => \N__9294\,
            DOUT => \N__9293\,
            PACKAGEPIN => \A_AMIGA_wire\(1)
        );

    \A_AMIGA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9295\,
            PADOUT => \N__9294\,
            PADIN => \N__9293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2760\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9286\,
            DIN => \N__9285\,
            DOUT => \N__9284\,
            PACKAGEPIN => D_LM_040(7)
        );

    \D_LM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9286\,
            PADOUT => \N__9285\,
            PADIN => \N__9284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6970\,
            DIN0 => \D_LM_040_in_7\,
            DOUT0 => \N__3780\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9277\,
            DIN => \N__9276\,
            DOUT => \N__9275\,
            PACKAGEPIN => D_UM_040(4)
        );

    \D_UM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9277\,
            PADOUT => \N__9276\,
            PADIN => \N__9275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7005\,
            DIN0 => \D_UM_040_in_4\,
            DOUT0 => \N__7542\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9268\,
            DIN => \N__9267\,
            DOUT => \N__9266\,
            PACKAGEPIN => \CLK40B_wire\
        );

    \CLK40B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9268\,
            PADOUT => \N__9267\,
            PADIN => \N__9266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5764\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9259\,
            DIN => \N__9258\,
            DOUT => \N__9257\,
            PACKAGEPIN => D_UU_AMIGA(0)
        );

    \D_UU_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9259\,
            PADOUT => \N__9258\,
            PADIN => \N__9257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4878\,
            DIN0 => \D_UU_AMIGA_in_0\,
            DOUT0 => \N__2964\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9250\,
            DIN => \N__9249\,
            DOUT => \N__9248\,
            PACKAGEPIN => D_UM_040(1)
        );

    \D_UM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9250\,
            PADOUT => \N__9249\,
            PADIN => \N__9248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6849\,
            DIN0 => \D_UM_040_in_1\,
            DOUT0 => \N__4347\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9241\,
            DIN => \N__9240\,
            DOUT => \N__9239\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9241\,
            PADOUT => \N__9240\,
            PADIN => \N__9239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TBIn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9232\,
            DIN => \N__9231\,
            DOUT => \N__9230\,
            PACKAGEPIN => D_LL_040(4)
        );

    \D_LL_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9232\,
            PADOUT => \N__9231\,
            PADIN => \N__9230\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6909\,
            DIN0 => \D_LL_040_in_4\,
            DOUT0 => \N__2706\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9223\,
            DIN => \N__9222\,
            DOUT => \N__9221\,
            PACKAGEPIN => D_LL_AMIGA(7)
        );

    \D_LL_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9223\,
            PADOUT => \N__9222\,
            PADIN => \N__9221\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4863\,
            DIN0 => \D_LL_AMIGA_in_7\,
            DOUT0 => \N__5199\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9214\,
            DIN => \N__9213\,
            DOUT => \N__9212\,
            PACKAGEPIN => D_UU_AMIGA(7)
        );

    \D_UU_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9214\,
            PADOUT => \N__9213\,
            PADIN => \N__9212\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4914\,
            DIN0 => \D_UU_AMIGA_in_7\,
            DOUT0 => \N__8013\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9205\,
            DIN => \N__9204\,
            DOUT => \N__9203\,
            PACKAGEPIN => \BUFDIR_wire\
        );

    \BUFDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9205\,
            PADOUT => \N__9204\,
            PADIN => \N__9203\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4284\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9196\,
            DIN => \N__9195\,
            DOUT => \N__9194\,
            PACKAGEPIN => D_UU_040(4)
        );

    \D_UU_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9196\,
            PADOUT => \N__9195\,
            PADIN => \N__9194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6936\,
            DIN0 => \D_UU_040_in_4\,
            DOUT0 => \N__5406\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9187\,
            DIN => \N__9186\,
            DOUT => \N__9185\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9187\,
            PADOUT => \N__9186\,
            PADIN => \N__9185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9178\,
            DIN => \N__9177\,
            DOUT => \N__9176\,
            PACKAGEPIN => D_LL_040(1)
        );

    \D_LL_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9178\,
            PADOUT => \N__9177\,
            PADIN => \N__9176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6908\,
            DIN0 => \D_LL_040_in_1\,
            DOUT0 => \N__2673\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9169\,
            DIN => \N__9168\,
            DOUT => \N__9167\,
            PACKAGEPIN => D_UM_AMIGA(5)
        );

    \D_UM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9169\,
            PADOUT => \N__9168\,
            PADIN => \N__9167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4879\,
            DIN0 => \D_UM_AMIGA_in_5\,
            DOUT0 => \N__8574\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9160\,
            DIN => \N__9159\,
            DOUT => \N__9158\,
            PACKAGEPIN => D_UU_040(1)
        );

    \D_UU_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9160\,
            PADOUT => \N__9159\,
            PADIN => \N__9158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7011\,
            DIN0 => \D_UU_040_in_1\,
            DOUT0 => \N__6243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9151\,
            DIN => \N__9150\,
            DOUT => \N__9149\,
            PACKAGEPIN => D_LM_AMIGA(1)
        );

    \D_LM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9151\,
            PADOUT => \N__9150\,
            PADIN => \N__9149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4775\,
            DIN0 => \D_LM_AMIGA_in_1\,
            DOUT0 => \N__5277\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9142\,
            DIN => \N__9141\,
            DOUT => \N__9140\,
            PACKAGEPIN => D_LM_040(2)
        );

    \D_LM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9142\,
            PADOUT => \N__9141\,
            PADIN => \N__9140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6860\,
            DIN0 => \D_LM_040_in_2\,
            DOUT0 => \N__3045\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9133\,
            DIN => \N__9132\,
            DOUT => \N__9131\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9133\,
            PADOUT => \N__9132\,
            PADIN => \N__9131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7374\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__2793\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9124\,
            DIN => \N__9123\,
            DOUT => \N__9122\,
            PACKAGEPIN => D_UM_040(2)
        );

    \D_UM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9124\,
            PADOUT => \N__9123\,
            PADIN => \N__9122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6924\,
            DIN0 => \D_UM_040_in_2\,
            DOUT0 => \N__6663\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9115\,
            DIN => \N__9114\,
            DOUT => \N__9113\,
            PACKAGEPIN => \CLKRAMB_wire\
        );

    \CLKRAMB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9115\,
            PADOUT => \N__9114\,
            PADIN => \N__9113\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8189\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9106\,
            DIN => \N__9105\,
            DOUT => \N__9104\,
            PACKAGEPIN => D_LL_AMIGA(2)
        );

    \D_LL_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9106\,
            PADOUT => \N__9105\,
            PADIN => \N__9104\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4735\,
            DIN0 => \D_LL_AMIGA_in_2\,
            DOUT0 => \N__8283\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9097\,
            DIN => \N__9096\,
            DOUT => \N__9095\,
            PACKAGEPIN => D_UU_AMIGA(2)
        );

    \D_UU_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9097\,
            PADOUT => \N__9096\,
            PADIN => \N__9095\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4877\,
            DIN0 => \D_UU_AMIGA_in_2\,
            DOUT0 => \N__3609\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEAn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9088\,
            DIN => \N__9087\,
            DOUT => \N__9086\,
            PACKAGEPIN => \TEAn_wire\
        );

    \TEAn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9088\,
            PADOUT => \N__9087\,
            PADIN => \N__9086\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TEAn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9079\,
            DIN => \N__9078\,
            DOUT => \N__9077\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9079\,
            PADOUT => \N__9078\,
            PADIN => \N__9077\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4296\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9070\,
            DIN => \N__9069\,
            DOUT => \N__9068\,
            PACKAGEPIN => D_LL_040(6)
        );

    \D_LL_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9070\,
            PADOUT => \N__9069\,
            PADIN => \N__9068\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6961\,
            DIN0 => \D_LL_040_in_6\,
            DOUT0 => \N__5901\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9061\,
            DIN => \N__9060\,
            DOUT => \N__9059\,
            PACKAGEPIN => D_LL_AMIGA(5)
        );

    \D_LL_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9061\,
            PADOUT => \N__9060\,
            PADIN => \N__9059\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4866\,
            DIN0 => \D_LL_AMIGA_in_5\,
            DOUT0 => \N__7983\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9052\,
            DIN => \N__9051\,
            DOUT => \N__9050\,
            PACKAGEPIN => D_UM_AMIGA(0)
        );

    \D_UM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9052\,
            PADOUT => \N__9051\,
            PADIN => \N__9050\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4839\,
            DIN0 => \D_UM_AMIGA_in_0\,
            DOUT0 => \N__3222\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9043\,
            DIN => \N__9042\,
            DOUT => \N__9041\,
            PACKAGEPIN => D_UU_040(2)
        );

    \D_UU_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9043\,
            PADOUT => \N__9042\,
            PADIN => \N__9041\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6852\,
            DIN0 => \D_UU_040_in_2\,
            DOUT0 => \N__3696\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9034\,
            DIN => \N__9033\,
            DOUT => \N__9032\,
            PACKAGEPIN => TSn
        );

    \TSn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9034\,
            PADOUT => \N__9033\,
            PADIN => \N__9032\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3591\,
            DIN0 => \TSn_in\,
            DOUT0 => \N__4098\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9025\,
            DIN => \N__9024\,
            DOUT => \N__9023\,
            PACKAGEPIN => D_LM_AMIGA(2)
        );

    \D_LM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9025\,
            PADOUT => \N__9024\,
            PADIN => \N__9023\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4838\,
            DIN0 => \D_LM_AMIGA_in_2\,
            DOUT0 => \N__3651\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TS_CPUn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9016\,
            DIN => \N__9015\,
            DOUT => \N__9014\,
            PACKAGEPIN => TS_CPUn
        );

    \TS_CPUn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9016\,
            PADOUT => \N__9015\,
            PADIN => \N__9014\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7271\,
            DIN0 => \TS_CPUn_in\,
            DOUT0 => \N__2649\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK80_CPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9007\,
            DIN => \N__9006\,
            DOUT => \N__9005\,
            PACKAGEPIN => \CLK80_CPU_wire\
        );

    \CLK80_CPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9007\,
            PADOUT => \N__9006\,
            PADIN => \N__9005\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8193\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8998\,
            DIN => \N__8997\,
            DOUT => \N__8996\,
            PACKAGEPIN => D_LL_040(3)
        );

    \D_LL_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8998\,
            PADOUT => \N__8997\,
            PADIN => \N__8996\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6994\,
            DIN0 => \D_LL_040_in_3\,
            DOUT0 => \N__3495\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8989\,
            DIN => \N__8988\,
            DOUT => \N__8987\,
            PACKAGEPIN => D_LM_040(1)
        );

    \D_LM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8989\,
            PADOUT => \N__8988\,
            PADIN => \N__8987\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6859\,
            DIN0 => \D_LM_040_in_1\,
            DOUT0 => \N__3156\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8980\,
            DIN => \N__8979\,
            DOUT => \N__8978\,
            PACKAGEPIN => D_UM_AMIGA(7)
        );

    \D_UM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8980\,
            PADOUT => \N__8979\,
            PADIN => \N__8978\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4916\,
            DIN0 => \D_UM_AMIGA_in_7\,
            DOUT0 => \N__5151\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8971\,
            DIN => \N__8970\,
            DOUT => \N__8969\,
            PACKAGEPIN => D_LM_AMIGA(7)
        );

    \D_LM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8971\,
            PADOUT => \N__8970\,
            PADIN => \N__8969\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4891\,
            DIN0 => \D_LM_AMIGA_in_7\,
            DOUT0 => \N__8055\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8962\,
            DIN => \N__8961\,
            DOUT => \N__8960\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8962\,
            PADOUT => \N__8961\,
            PADIN => \N__8960\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PORTSIZE_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8953\,
            DIN => \N__8952\,
            DOUT => \N__8951\,
            PACKAGEPIN => \A_AMIGA_wire\(0)
        );

    \A_AMIGA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8953\,
            PADOUT => \N__8952\,
            PADIN => \N__8951\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2736\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8944\,
            DIN => \N__8943\,
            DOUT => \N__8942\,
            PACKAGEPIN => D_LM_040(4)
        );

    \D_LM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8944\,
            PADOUT => \N__8943\,
            PADIN => \N__8942\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6927\,
            DIN0 => \D_LM_040_in_4\,
            DOUT0 => \N__4431\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8935\,
            DIN => \N__8934\,
            DOUT => \N__8933\,
            PACKAGEPIN => D_UM_040(7)
        );

    \D_UM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8935\,
            PADOUT => \N__8934\,
            PADIN => \N__8933\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7009\,
            DIN0 => \D_UM_040_in_7\,
            DOUT0 => \N__4998\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8926\,
            DIN => \N__8925\,
            DOUT => \N__8924\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8926\,
            PADOUT => \N__8925\,
            PADIN => \N__8924\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8917\,
            DIN => \N__8916\,
            DOUT => \N__8915\,
            PACKAGEPIN => D_UU_AMIGA(1)
        );

    \D_UU_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8917\,
            PADOUT => \N__8916\,
            PADIN => \N__8915\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4917\,
            DIN0 => \D_UU_AMIGA_in_1\,
            DOUT0 => \N__5235\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8908\,
            DIN => \N__8907\,
            DOUT => \N__8906\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8908\,
            PADOUT => \N__8907\,
            PADIN => \N__8906\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5754\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8899\,
            DIN => \N__8898\,
            DOUT => \N__8897\,
            PACKAGEPIN => D_UM_040(0)
        );

    \D_UM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8899\,
            PADOUT => \N__8898\,
            PADIN => \N__8897\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6925\,
            DIN0 => \D_UM_040_in_0\,
            DOUT0 => \N__8499\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8890\,
            DIN => \N__8889\,
            DOUT => \N__8888\,
            PACKAGEPIN => D_LL_AMIGA(0)
        );

    \D_LL_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8890\,
            PADOUT => \N__8889\,
            PADIN => \N__8888\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4929\,
            DIN0 => \D_LL_AMIGA_in_0\,
            DOUT0 => \N__3264\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8881\,
            DIN => \N__8880\,
            DOUT => \N__8879\,
            PACKAGEPIN => D_UU_AMIGA(4)
        );

    \D_UU_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8881\,
            PADOUT => \N__8880\,
            PADIN => \N__8879\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4876\,
            DIN0 => \D_UU_AMIGA_in_4\,
            DOUT0 => \N__2886\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8872\,
            DIN => \N__8871\,
            DOUT => \N__8870\,
            PACKAGEPIN => D_UU_040(7)
        );

    \D_UU_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8872\,
            PADOUT => \N__8871\,
            PADIN => \N__8870\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6972\,
            DIN0 => \D_UU_040_in_7\,
            DOUT0 => \N__5490\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8863\,
            DIN => \N__8862\,
            DOUT => \N__8861\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8863\,
            PADOUT => \N__8862\,
            PADIN => \N__8861\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BGn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8854\,
            DIN => \N__8853\,
            DOUT => \N__8852\,
            PACKAGEPIN => \BGn_wire\
        );

    \BGn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8854\,
            PADOUT => \N__8853\,
            PADIN => \N__8852\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BGn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8845\,
            DIN => \N__8844\,
            DOUT => \N__8843\,
            PACKAGEPIN => D_LL_040(0)
        );

    \D_LL_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8845\,
            PADOUT => \N__8844\,
            PADIN => \N__8843\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6995\,
            DIN0 => \D_LL_040_in_0\,
            DOUT0 => \N__7347\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8836\,
            DIN => \N__8835\,
            DOUT => \N__8834\,
            PACKAGEPIN => D_UM_AMIGA(2)
        );

    \D_UM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8836\,
            PADOUT => \N__8835\,
            PADIN => \N__8834\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4841\,
            DIN0 => \D_UM_AMIGA_in_2\,
            DOUT0 => \N__8226\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8827\,
            DIN => \N__8826\,
            DOUT => \N__8825\,
            PACKAGEPIN => D_UU_040(0)
        );

    \D_UU_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8827\,
            PADOUT => \N__8826\,
            PADIN => \N__8825\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6971\,
            DIN0 => \D_UU_040_in_0\,
            DOUT0 => \N__6159\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8818\,
            DIN => \N__8817\,
            DOUT => \N__8816\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8818\,
            PADOUT => \N__8817\,
            PADIN => \N__8816\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TCIn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8809\,
            DIN => \N__8808\,
            DOUT => \N__8807\,
            PACKAGEPIN => \A_040_wire\(0)
        );

    \A_040_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8809\,
            PADOUT => \N__8808\,
            PADIN => \N__8807\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8800\,
            DIN => \N__8799\,
            DOUT => \N__8798\,
            PACKAGEPIN => D_LM_AMIGA(0)
        );

    \D_LM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8800\,
            PADOUT => \N__8799\,
            PADIN => \N__8798\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4864\,
            DIN0 => \D_LM_AMIGA_in_0\,
            DOUT0 => \N__3030\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8791\,
            DIN => \N__8790\,
            DOUT => \N__8789\,
            PACKAGEPIN => \TBI_CPUn_wire\
        );

    \TBI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8791\,
            PADOUT => \N__8790\,
            PADIN => \N__8789\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4070\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8782\,
            DIN => \N__8781\,
            DOUT => \N__8780\,
            PACKAGEPIN => \CLK40A_wire\
        );

    \CLK40A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8782\,
            PADOUT => \N__8781\,
            PADIN => \N__8780\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5768\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8773\,
            DIN => \N__8772\,
            DOUT => \N__8771\,
            PACKAGEPIN => D_LM_040(3)
        );

    \D_LM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8773\,
            PADOUT => \N__8772\,
            PADIN => \N__8771\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6969\,
            DIN0 => \D_LM_040_in_3\,
            DOUT0 => \N__3189\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8764\,
            DIN => \N__8763\,
            DOUT => \N__8762\,
            PACKAGEPIN => D_LM_AMIGA(5)
        );

    \D_LM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8764\,
            PADOUT => \N__8763\,
            PADIN => \N__8762\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4889\,
            DIN0 => \D_LM_AMIGA_in_5\,
            DOUT0 => \N__7506\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8755\,
            DIN => \N__8754\,
            DOUT => \N__8753\,
            PACKAGEPIN => D_LM_040(6)
        );

    \D_LM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8755\,
            PADOUT => \N__8754\,
            PADIN => \N__8753\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6932\,
            DIN0 => \D_LM_040_in_6\,
            DOUT0 => \N__4308\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8746\,
            DIN => \N__8745\,
            DOUT => \N__8744\,
            PACKAGEPIN => D_UM_040(5)
        );

    \D_UM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8746\,
            PADOUT => \N__8745\,
            PADIN => \N__8744\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6996\,
            DIN0 => \D_UM_040_in_5\,
            DOUT0 => \N__7635\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8737\,
            DIN => \N__8736\,
            DOUT => \N__8735\,
            PACKAGEPIN => D_LL_AMIGA(3)
        );

    \D_LL_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8737\,
            PADOUT => \N__8736\,
            PADIN => \N__8735\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4734\,
            DIN0 => \D_LL_AMIGA_in_3\,
            DOUT0 => \N__3878\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8728\,
            DIN => \N__8727\,
            DOUT => \N__8726\,
            PACKAGEPIN => D_UU_AMIGA(3)
        );

    \D_UU_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8728\,
            PADOUT => \N__8727\,
            PADIN => \N__8726\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4932\,
            DIN0 => \D_UU_AMIGA_in_3\,
            DOUT0 => \N__8094\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8719\,
            DIN => \N__8718\,
            DOUT => \N__8717\,
            PACKAGEPIN => D_LL_040(5)
        );

    \D_LL_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8719\,
            PADOUT => \N__8718\,
            PADIN => \N__8717\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6960\,
            DIN0 => \D_LL_040_in_5\,
            DOUT0 => \N__5862\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8710\,
            DIN => \N__8709\,
            DOUT => \N__8708\,
            PACKAGEPIN => D_LL_AMIGA(6)
        );

    \D_LL_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8710\,
            PADOUT => \N__8709\,
            PADIN => \N__8708\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4865\,
            DIN0 => \D_LL_AMIGA_in_6\,
            DOUT0 => \N__3135\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8701\,
            DIN => \N__8700\,
            DOUT => \N__8699\,
            PACKAGEPIN => D_UU_AMIGA(6)
        );

    \D_UU_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8701\,
            PADOUT => \N__8700\,
            PADIN => \N__8699\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4915\,
            DIN0 => \D_UU_AMIGA_in_6\,
            DOUT0 => \N__2811\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8692\,
            DIN => \N__8691\,
            DOUT => \N__8690\,
            PACKAGEPIN => D_UM_AMIGA(1)
        );

    \D_UM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8692\,
            PADOUT => \N__8691\,
            PADIN => \N__8690\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4890\,
            DIN0 => \D_UM_AMIGA_in_1\,
            DOUT0 => \N__3294\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8683\,
            DIN => \N__8682\,
            DOUT => \N__8681\,
            PACKAGEPIN => D_UU_040(5)
        );

    \D_UU_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8683\,
            PADOUT => \N__8682\,
            PADIN => \N__8681\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6997\,
            DIN0 => \D_UU_040_in_5\,
            DOUT0 => \N__5565\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8674\,
            DIN => \N__8673\,
            DOUT => \N__8672\,
            PACKAGEPIN => \CLKRAMA_wire\
        );

    \CLKRAMA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8674\,
            PADOUT => \N__8673\,
            PADIN => \N__8672\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5772\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8665\,
            DIN => \N__8664\,
            DOUT => \N__8663\,
            PACKAGEPIN => D_LL_040(2)
        );

    \D_LL_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8665\,
            PADOUT => \N__8664\,
            PADIN => \N__8663\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6962\,
            DIN0 => \D_LL_040_in_2\,
            DOUT0 => \N__3534\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8656\,
            DIN => \N__8655\,
            DOUT => \N__8654\,
            PACKAGEPIN => \TCI_CPUn_wire\
        );

    \TCI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8656\,
            PADOUT => \N__8655\,
            PADIN => \N__8654\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2622\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BBn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8647\,
            DIN => \N__8646\,
            DOUT => \N__8645\,
            PACKAGEPIN => \BBn_wire\
        );

    \BBn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8647\,
            PADOUT => \N__8646\,
            PADIN => \N__8645\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BBn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMAAn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8638\,
            DIN => \N__8637\,
            DOUT => \N__8636\,
            PACKAGEPIN => \DMAAn_wire\
        );

    \DMAAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8638\,
            PADOUT => \N__8637\,
            PADIN => \N__8636\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4245\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8629\,
            DIN => \N__8628\,
            DOUT => \N__8627\,
            PACKAGEPIN => D_UM_AMIGA(4)
        );

    \D_UM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8629\,
            PADOUT => \N__8628\,
            PADIN => \N__8627\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4919\,
            DIN0 => \D_UM_AMIGA_in_4\,
            DOUT0 => \N__5937\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8620\,
            DIN => \N__8619\,
            DOUT => \N__8618\,
            PACKAGEPIN => D_LM_AMIGA(6)
        );

    \D_LM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8620\,
            PADOUT => \N__8619\,
            PADIN => \N__8618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4892\,
            DIN0 => \D_LM_AMIGA_in_6\,
            DOUT0 => \N__2850\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8611\,
            DIN => \N__8610\,
            DOUT => \N__8609\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8611\,
            PADOUT => \N__8610\,
            PADIN => \N__8609\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8602\,
            DIN => \N__8601\,
            DOUT => \N__8600\,
            PACKAGEPIN => D_LM_040(5)
        );

    \D_LM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8602\,
            PADOUT => \N__8601\,
            PADIN => \N__8600\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6926\,
            DIN0 => \D_LM_040_in_5\,
            DOUT0 => \N__3957\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8593\,
            DIN => \N__8592\,
            DOUT => \N__8591\,
            PACKAGEPIN => D_UM_040(6)
        );

    \D_UM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8593\,
            PADOUT => \N__8592\,
            PADIN => \N__8591\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6931\,
            DIN0 => \D_UM_040_in_6\,
            DOUT0 => \N__8304\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2213\ : IoInMux
    port map (
            O => \N__8574\,
            I => \N__8571\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__8571\,
            I => \N__8568\
        );

    \I__2211\ : IoSpan4Mux
    port map (
            O => \N__8568\,
            I => \N__8565\
        );

    \I__2210\ : Sp12to4
    port map (
            O => \N__8565\,
            I => \N__8562\
        );

    \I__2209\ : Span12Mux_s6_v
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__2208\ : Odrv12
    port map (
            O => \N__8559\,
            I => \un1_D_UM_040_5\
        );

    \I__2207\ : InMux
    port map (
            O => \N__8556\,
            I => \N__8552\
        );

    \I__2206\ : InMux
    port map (
            O => \N__8555\,
            I => \N__8549\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__8552\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__8549\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__2203\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8541\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__8541\,
            I => \N__8537\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__8540\,
            I => \N__8534\
        );

    \I__2200\ : Span4Mux_v
    port map (
            O => \N__8537\,
            I => \N__8531\
        );

    \I__2199\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8528\
        );

    \I__2198\ : Span4Mux_v
    port map (
            O => \N__8531\,
            I => \N__8523\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__8528\,
            I => \N__8523\
        );

    \I__2196\ : Span4Mux_v
    port map (
            O => \N__8523\,
            I => \N__8520\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__8520\,
            I => \N__8516\
        );

    \I__2194\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8513\
        );

    \I__2193\ : Span4Mux_h
    port map (
            O => \N__8516\,
            I => \N__8510\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__8513\,
            I => \N__8507\
        );

    \I__2191\ : Sp12to4
    port map (
            O => \N__8510\,
            I => \N__8502\
        );

    \I__2190\ : Span12Mux_h
    port map (
            O => \N__8507\,
            I => \N__8502\
        );

    \I__2189\ : Odrv12
    port map (
            O => \N__8502\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__2188\ : IoInMux
    port map (
            O => \N__8499\,
            I => \N__8496\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__8496\,
            I => \N__8493\
        );

    \I__2186\ : IoSpan4Mux
    port map (
            O => \N__8493\,
            I => \N__8490\
        );

    \I__2185\ : Span4Mux_s2_h
    port map (
            O => \N__8490\,
            I => \N__8487\
        );

    \I__2184\ : Sp12to4
    port map (
            O => \N__8487\,
            I => \N__8484\
        );

    \I__2183\ : Span12Mux_s11_h
    port map (
            O => \N__8484\,
            I => \N__8481\
        );

    \I__2182\ : Odrv12
    port map (
            O => \N__8481\,
            I => \un1_D_UM_AMIGA_0\
        );

    \I__2181\ : InMux
    port map (
            O => \N__8478\,
            I => \N__8474\
        );

    \I__2180\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8471\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__8474\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__8471\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__2177\ : InMux
    port map (
            O => \N__8466\,
            I => \N__8462\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__8465\,
            I => \N__8459\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__8462\,
            I => \N__8456\
        );

    \I__2174\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8453\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__8456\,
            I => \N__8447\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__8453\,
            I => \N__8447\
        );

    \I__2171\ : InMux
    port map (
            O => \N__8452\,
            I => \N__8444\
        );

    \I__2170\ : Span4Mux_v
    port map (
            O => \N__8447\,
            I => \N__8441\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__8444\,
            I => \N__8436\
        );

    \I__2168\ : Sp12to4
    port map (
            O => \N__8441\,
            I => \N__8436\
        );

    \I__2167\ : Span12Mux_h
    port map (
            O => \N__8436\,
            I => \N__8433\
        );

    \I__2166\ : Span12Mux_v
    port map (
            O => \N__8433\,
            I => \N__8430\
        );

    \I__2165\ : Odrv12
    port map (
            O => \N__8430\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__2164\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8416\
        );

    \I__2163\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8416\
        );

    \I__2162\ : InMux
    port map (
            O => \N__8425\,
            I => \N__8411\
        );

    \I__2161\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8411\
        );

    \I__2160\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8408\
        );

    \I__2159\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8405\
        );

    \I__2158\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8398\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__8416\,
            I => \N__8393\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__8411\,
            I => \N__8390\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__8408\,
            I => \N__8385\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__8405\,
            I => \N__8385\
        );

    \I__2153\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8382\
        );

    \I__2152\ : InMux
    port map (
            O => \N__8403\,
            I => \N__8375\
        );

    \I__2151\ : InMux
    port map (
            O => \N__8402\,
            I => \N__8375\
        );

    \I__2150\ : InMux
    port map (
            O => \N__8401\,
            I => \N__8375\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__8398\,
            I => \N__8372\
        );

    \I__2148\ : InMux
    port map (
            O => \N__8397\,
            I => \N__8369\
        );

    \I__2147\ : InMux
    port map (
            O => \N__8396\,
            I => \N__8366\
        );

    \I__2146\ : Span4Mux_v
    port map (
            O => \N__8393\,
            I => \N__8360\
        );

    \I__2145\ : Span4Mux_h
    port map (
            O => \N__8390\,
            I => \N__8351\
        );

    \I__2144\ : Span4Mux_v
    port map (
            O => \N__8385\,
            I => \N__8351\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__8382\,
            I => \N__8351\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__8375\,
            I => \N__8351\
        );

    \I__2141\ : Span4Mux_v
    port map (
            O => \N__8372\,
            I => \N__8346\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__8369\,
            I => \N__8346\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__8366\,
            I => \N__8343\
        );

    \I__2138\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8338\
        );

    \I__2137\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8338\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__8363\,
            I => \N__8334\
        );

    \I__2135\ : Span4Mux_v
    port map (
            O => \N__8360\,
            I => \N__8331\
        );

    \I__2134\ : Span4Mux_v
    port map (
            O => \N__8351\,
            I => \N__8328\
        );

    \I__2133\ : Span4Mux_v
    port map (
            O => \N__8346\,
            I => \N__8321\
        );

    \I__2132\ : Span4Mux_v
    port map (
            O => \N__8343\,
            I => \N__8321\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__8338\,
            I => \N__8321\
        );

    \I__2130\ : InMux
    port map (
            O => \N__8337\,
            I => \N__8318\
        );

    \I__2129\ : InMux
    port map (
            O => \N__8334\,
            I => \N__8315\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__8331\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__8328\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__2126\ : Odrv4
    port map (
            O => \N__8321\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__8318\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__8315\,
            I => \U111_CYCLE_SM.LATCH_ENZ0\
        );

    \I__2123\ : IoInMux
    port map (
            O => \N__8304\,
            I => \N__8301\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__8301\,
            I => \N__8298\
        );

    \I__2121\ : IoSpan4Mux
    port map (
            O => \N__8298\,
            I => \N__8295\
        );

    \I__2120\ : Span4Mux_s0_h
    port map (
            O => \N__8295\,
            I => \N__8292\
        );

    \I__2119\ : Sp12to4
    port map (
            O => \N__8292\,
            I => \N__8289\
        );

    \I__2118\ : Span12Mux_s7_h
    port map (
            O => \N__8289\,
            I => \N__8286\
        );

    \I__2117\ : Odrv12
    port map (
            O => \N__8286\,
            I => \N_125\
        );

    \I__2116\ : IoInMux
    port map (
            O => \N__8283\,
            I => \N__8280\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__8280\,
            I => \N__8276\
        );

    \I__2114\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8273\
        );

    \I__2113\ : IoSpan4Mux
    port map (
            O => \N__8276\,
            I => \N__8270\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__8273\,
            I => \N__8267\
        );

    \I__2111\ : Span4Mux_s2_h
    port map (
            O => \N__8270\,
            I => \N__8264\
        );

    \I__2110\ : Span4Mux_v
    port map (
            O => \N__8267\,
            I => \N__8261\
        );

    \I__2109\ : Sp12to4
    port map (
            O => \N__8264\,
            I => \N__8258\
        );

    \I__2108\ : Sp12to4
    port map (
            O => \N__8261\,
            I => \N__8255\
        );

    \I__2107\ : Span12Mux_h
    port map (
            O => \N__8258\,
            I => \N__8252\
        );

    \I__2106\ : Span12Mux_h
    port map (
            O => \N__8255\,
            I => \N__8249\
        );

    \I__2105\ : Span12Mux_h
    port map (
            O => \N__8252\,
            I => \N__8246\
        );

    \I__2104\ : Span12Mux_v
    port map (
            O => \N__8249\,
            I => \N__8243\
        );

    \I__2103\ : Odrv12
    port map (
            O => \N__8246\,
            I => \D_LL_040_in_2\
        );

    \I__2102\ : Odrv12
    port map (
            O => \N__8243\,
            I => \D_LL_040_in_2\
        );

    \I__2101\ : InMux
    port map (
            O => \N__8238\,
            I => \N__8235\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__8235\,
            I => \N__8232\
        );

    \I__2099\ : Span12Mux_h
    port map (
            O => \N__8232\,
            I => \N__8229\
        );

    \I__2098\ : Odrv12
    port map (
            O => \N__8229\,
            I => \D_UM_040_in_2\
        );

    \I__2097\ : IoInMux
    port map (
            O => \N__8226\,
            I => \N__8223\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__8223\,
            I => \N__8220\
        );

    \I__2095\ : Span4Mux_s3_h
    port map (
            O => \N__8220\,
            I => \N__8217\
        );

    \I__2094\ : Sp12to4
    port map (
            O => \N__8217\,
            I => \N__8214\
        );

    \I__2093\ : Span12Mux_v
    port map (
            O => \N__8214\,
            I => \N__8211\
        );

    \I__2092\ : Span12Mux_h
    port map (
            O => \N__8211\,
            I => \N__8208\
        );

    \I__2091\ : Odrv12
    port map (
            O => \N__8208\,
            I => \un1_D_UM_040_2\
        );

    \I__2090\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8202\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__8202\,
            I => \N__8199\
        );

    \I__2088\ : Glb2LocalMux
    port map (
            O => \N__8199\,
            I => \N__8196\
        );

    \I__2087\ : GlobalMux
    port map (
            O => \N__8196\,
            I => \CLK80\
        );

    \I__2086\ : IoInMux
    port map (
            O => \N__8193\,
            I => \N__8190\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__8190\,
            I => \N__8186\
        );

    \I__2084\ : IoInMux
    port map (
            O => \N__8189\,
            I => \N__8183\
        );

    \I__2083\ : IoSpan4Mux
    port map (
            O => \N__8186\,
            I => \N__8180\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__8183\,
            I => \N__8177\
        );

    \I__2081\ : Sp12to4
    port map (
            O => \N__8180\,
            I => \N__8174\
        );

    \I__2080\ : Span12Mux_s3_v
    port map (
            O => \N__8177\,
            I => \N__8171\
        );

    \I__2079\ : Span12Mux_s7_h
    port map (
            O => \N__8174\,
            I => \N__8168\
        );

    \I__2078\ : Span12Mux_v
    port map (
            O => \N__8171\,
            I => \N__8165\
        );

    \I__2077\ : Odrv12
    port map (
            O => \N__8168\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__2076\ : Odrv12
    port map (
            O => \N__8165\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__2075\ : InMux
    port map (
            O => \N__8160\,
            I => \N__8157\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__8157\,
            I => \N__8154\
        );

    \I__2073\ : Span4Mux_v
    port map (
            O => \N__8154\,
            I => \N__8151\
        );

    \I__2072\ : Span4Mux_h
    port map (
            O => \N__8151\,
            I => \N__8148\
        );

    \I__2071\ : Sp12to4
    port map (
            O => \N__8148\,
            I => \N__8145\
        );

    \I__2070\ : Span12Mux_h
    port map (
            O => \N__8145\,
            I => \N__8142\
        );

    \I__2069\ : Odrv12
    port map (
            O => \N__8142\,
            I => \D_UU_040_in_3\
        );

    \I__2068\ : IoInMux
    port map (
            O => \N__8139\,
            I => \N__8136\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__8136\,
            I => \N__8133\
        );

    \I__2066\ : IoSpan4Mux
    port map (
            O => \N__8133\,
            I => \N__8129\
        );

    \I__2065\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8126\
        );

    \I__2064\ : IoSpan4Mux
    port map (
            O => \N__8129\,
            I => \N__8123\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__8126\,
            I => \N__8120\
        );

    \I__2062\ : Span4Mux_s2_h
    port map (
            O => \N__8123\,
            I => \N__8117\
        );

    \I__2061\ : Span4Mux_v
    port map (
            O => \N__8120\,
            I => \N__8114\
        );

    \I__2060\ : Sp12to4
    port map (
            O => \N__8117\,
            I => \N__8111\
        );

    \I__2059\ : Sp12to4
    port map (
            O => \N__8114\,
            I => \N__8108\
        );

    \I__2058\ : Span12Mux_h
    port map (
            O => \N__8111\,
            I => \N__8105\
        );

    \I__2057\ : Span12Mux_h
    port map (
            O => \N__8108\,
            I => \N__8102\
        );

    \I__2056\ : Span12Mux_h
    port map (
            O => \N__8105\,
            I => \N__8097\
        );

    \I__2055\ : Span12Mux_v
    port map (
            O => \N__8102\,
            I => \N__8097\
        );

    \I__2054\ : Odrv12
    port map (
            O => \N__8097\,
            I => \D_LM_040_in_3\
        );

    \I__2053\ : IoInMux
    port map (
            O => \N__8094\,
            I => \N__8091\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__8091\,
            I => \N__8088\
        );

    \I__2051\ : Span4Mux_s2_v
    port map (
            O => \N__8088\,
            I => \N__8085\
        );

    \I__2050\ : Span4Mux_v
    port map (
            O => \N__8085\,
            I => \N__8082\
        );

    \I__2049\ : Sp12to4
    port map (
            O => \N__8082\,
            I => \N__8079\
        );

    \I__2048\ : Span12Mux_s11_h
    port map (
            O => \N__8079\,
            I => \N__8076\
        );

    \I__2047\ : Odrv12
    port map (
            O => \N__8076\,
            I => \un1_D_UU_040_3\
        );

    \I__2046\ : InMux
    port map (
            O => \N__8073\,
            I => \N__8070\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__8070\,
            I => \N__8067\
        );

    \I__2044\ : Span4Mux_v
    port map (
            O => \N__8067\,
            I => \N__8064\
        );

    \I__2043\ : Sp12to4
    port map (
            O => \N__8064\,
            I => \N__8061\
        );

    \I__2042\ : Span12Mux_h
    port map (
            O => \N__8061\,
            I => \N__8058\
        );

    \I__2041\ : Odrv12
    port map (
            O => \N__8058\,
            I => \D_UU_040_in_7\
        );

    \I__2040\ : IoInMux
    port map (
            O => \N__8055\,
            I => \N__8052\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__8052\,
            I => \N__8049\
        );

    \I__2038\ : IoSpan4Mux
    port map (
            O => \N__8049\,
            I => \N__8045\
        );

    \I__2037\ : InMux
    port map (
            O => \N__8048\,
            I => \N__8042\
        );

    \I__2036\ : Span4Mux_s2_h
    port map (
            O => \N__8045\,
            I => \N__8039\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__8042\,
            I => \N__8036\
        );

    \I__2034\ : Sp12to4
    port map (
            O => \N__8039\,
            I => \N__8033\
        );

    \I__2033\ : Span4Mux_v
    port map (
            O => \N__8036\,
            I => \N__8030\
        );

    \I__2032\ : Span12Mux_h
    port map (
            O => \N__8033\,
            I => \N__8027\
        );

    \I__2031\ : Sp12to4
    port map (
            O => \N__8030\,
            I => \N__8024\
        );

    \I__2030\ : Span12Mux_h
    port map (
            O => \N__8027\,
            I => \N__8021\
        );

    \I__2029\ : Span12Mux_h
    port map (
            O => \N__8024\,
            I => \N__8018\
        );

    \I__2028\ : Odrv12
    port map (
            O => \N__8021\,
            I => \D_LM_040_in_7\
        );

    \I__2027\ : Odrv12
    port map (
            O => \N__8018\,
            I => \D_LM_040_in_7\
        );

    \I__2026\ : IoInMux
    port map (
            O => \N__8013\,
            I => \N__8010\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__8010\,
            I => \N__8007\
        );

    \I__2024\ : Span12Mux_s8_v
    port map (
            O => \N__8007\,
            I => \N__8004\
        );

    \I__2023\ : Span12Mux_h
    port map (
            O => \N__8004\,
            I => \N__8001\
        );

    \I__2022\ : Odrv12
    port map (
            O => \N__8001\,
            I => \un1_D_UU_040_7\
        );

    \I__2021\ : IoInMux
    port map (
            O => \N__7998\,
            I => \N__7995\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__7995\,
            I => \N__7992\
        );

    \I__2019\ : Span4Mux_s2_v
    port map (
            O => \N__7992\,
            I => \N__7989\
        );

    \I__2018\ : Span4Mux_v
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__7986\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2016\ : IoInMux
    port map (
            O => \N__7983\,
            I => \N__7980\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__7980\,
            I => \N__7977\
        );

    \I__2014\ : IoSpan4Mux
    port map (
            O => \N__7977\,
            I => \N__7973\
        );

    \I__2013\ : InMux
    port map (
            O => \N__7976\,
            I => \N__7970\
        );

    \I__2012\ : Span4Mux_s2_h
    port map (
            O => \N__7973\,
            I => \N__7967\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__7970\,
            I => \N__7964\
        );

    \I__2010\ : Span4Mux_v
    port map (
            O => \N__7967\,
            I => \N__7961\
        );

    \I__2009\ : Sp12to4
    port map (
            O => \N__7964\,
            I => \N__7958\
        );

    \I__2008\ : Sp12to4
    port map (
            O => \N__7961\,
            I => \N__7955\
        );

    \I__2007\ : Span12Mux_v
    port map (
            O => \N__7958\,
            I => \N__7952\
        );

    \I__2006\ : Span12Mux_h
    port map (
            O => \N__7955\,
            I => \N__7947\
        );

    \I__2005\ : Span12Mux_v
    port map (
            O => \N__7952\,
            I => \N__7947\
        );

    \I__2004\ : Span12Mux_h
    port map (
            O => \N__7947\,
            I => \N__7944\
        );

    \I__2003\ : Odrv12
    port map (
            O => \N__7944\,
            I => \D_LL_040_in_5\
        );

    \I__2002\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7938\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__7938\,
            I => \N__7935\
        );

    \I__2000\ : Span4Mux_v
    port map (
            O => \N__7935\,
            I => \N__7932\
        );

    \I__1999\ : Sp12to4
    port map (
            O => \N__7932\,
            I => \N__7929\
        );

    \I__1998\ : Span12Mux_h
    port map (
            O => \N__7929\,
            I => \N__7926\
        );

    \I__1997\ : Odrv12
    port map (
            O => \N__7926\,
            I => \D_UM_040_in_5\
        );

    \I__1996\ : InMux
    port map (
            O => \N__7923\,
            I => \N__7910\
        );

    \I__1995\ : InMux
    port map (
            O => \N__7922\,
            I => \N__7910\
        );

    \I__1994\ : InMux
    port map (
            O => \N__7921\,
            I => \N__7910\
        );

    \I__1993\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7904\
        );

    \I__1992\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7904\
        );

    \I__1991\ : InMux
    port map (
            O => \N__7918\,
            I => \N__7898\
        );

    \I__1990\ : InMux
    port map (
            O => \N__7917\,
            I => \N__7890\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__7910\,
            I => \N__7887\
        );

    \I__1988\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7884\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__7904\,
            I => \N__7880\
        );

    \I__1986\ : InMux
    port map (
            O => \N__7903\,
            I => \N__7877\
        );

    \I__1985\ : InMux
    port map (
            O => \N__7902\,
            I => \N__7872\
        );

    \I__1984\ : InMux
    port map (
            O => \N__7901\,
            I => \N__7872\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__7898\,
            I => \N__7868\
        );

    \I__1982\ : InMux
    port map (
            O => \N__7897\,
            I => \N__7861\
        );

    \I__1981\ : InMux
    port map (
            O => \N__7896\,
            I => \N__7861\
        );

    \I__1980\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7861\
        );

    \I__1979\ : InMux
    port map (
            O => \N__7894\,
            I => \N__7856\
        );

    \I__1978\ : InMux
    port map (
            O => \N__7893\,
            I => \N__7856\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__7890\,
            I => \N__7853\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__7887\,
            I => \N__7847\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__7884\,
            I => \N__7844\
        );

    \I__1974\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7841\
        );

    \I__1973\ : Span4Mux_v
    port map (
            O => \N__7880\,
            I => \N__7834\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__7877\,
            I => \N__7834\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__7872\,
            I => \N__7831\
        );

    \I__1970\ : InMux
    port map (
            O => \N__7871\,
            I => \N__7828\
        );

    \I__1969\ : Span4Mux_v
    port map (
            O => \N__7868\,
            I => \N__7825\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__7861\,
            I => \N__7822\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__7856\,
            I => \N__7819\
        );

    \I__1966\ : Span4Mux_v
    port map (
            O => \N__7853\,
            I => \N__7814\
        );

    \I__1965\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7809\
        );

    \I__1964\ : InMux
    port map (
            O => \N__7851\,
            I => \N__7809\
        );

    \I__1963\ : InMux
    port map (
            O => \N__7850\,
            I => \N__7802\
        );

    \I__1962\ : Span4Mux_h
    port map (
            O => \N__7847\,
            I => \N__7795\
        );

    \I__1961\ : Span4Mux_v
    port map (
            O => \N__7844\,
            I => \N__7795\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__7841\,
            I => \N__7795\
        );

    \I__1959\ : InMux
    port map (
            O => \N__7840\,
            I => \N__7790\
        );

    \I__1958\ : InMux
    port map (
            O => \N__7839\,
            I => \N__7790\
        );

    \I__1957\ : Span4Mux_v
    port map (
            O => \N__7834\,
            I => \N__7787\
        );

    \I__1956\ : Span4Mux_h
    port map (
            O => \N__7831\,
            I => \N__7782\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__7828\,
            I => \N__7782\
        );

    \I__1954\ : Span4Mux_h
    port map (
            O => \N__7825\,
            I => \N__7777\
        );

    \I__1953\ : Span4Mux_v
    port map (
            O => \N__7822\,
            I => \N__7777\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__7819\,
            I => \N__7774\
        );

    \I__1951\ : InMux
    port map (
            O => \N__7818\,
            I => \N__7769\
        );

    \I__1950\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7769\
        );

    \I__1949\ : Span4Mux_h
    port map (
            O => \N__7814\,
            I => \N__7764\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__7809\,
            I => \N__7764\
        );

    \I__1947\ : InMux
    port map (
            O => \N__7808\,
            I => \N__7757\
        );

    \I__1946\ : InMux
    port map (
            O => \N__7807\,
            I => \N__7757\
        );

    \I__1945\ : InMux
    port map (
            O => \N__7806\,
            I => \N__7757\
        );

    \I__1944\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7754\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__7802\,
            I => \N__7747\
        );

    \I__1942\ : Span4Mux_v
    port map (
            O => \N__7795\,
            I => \N__7742\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__7790\,
            I => \N__7742\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__7787\,
            I => \N__7737\
        );

    \I__1939\ : Span4Mux_v
    port map (
            O => \N__7782\,
            I => \N__7737\
        );

    \I__1938\ : Span4Mux_v
    port map (
            O => \N__7777\,
            I => \N__7730\
        );

    \I__1937\ : Span4Mux_v
    port map (
            O => \N__7774\,
            I => \N__7730\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__7769\,
            I => \N__7730\
        );

    \I__1935\ : Sp12to4
    port map (
            O => \N__7764\,
            I => \N__7723\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__7757\,
            I => \N__7723\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__7754\,
            I => \N__7723\
        );

    \I__1932\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7716\
        );

    \I__1931\ : InMux
    port map (
            O => \N__7752\,
            I => \N__7716\
        );

    \I__1930\ : InMux
    port map (
            O => \N__7751\,
            I => \N__7716\
        );

    \I__1929\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7713\
        );

    \I__1928\ : Odrv12
    port map (
            O => \N__7747\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1927\ : Odrv4
    port map (
            O => \N__7742\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__7737\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__7730\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1924\ : Odrv12
    port map (
            O => \N__7723\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__7716\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__7713\,
            I => \U111_CYCLE_SM.FLIP_WORDZ0\
        );

    \I__1921\ : InMux
    port map (
            O => \N__7698\,
            I => \N__7695\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__7695\,
            I => \N__7691\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__7694\,
            I => \N__7688\
        );

    \I__1918\ : Span4Mux_v
    port map (
            O => \N__7691\,
            I => \N__7685\
        );

    \I__1917\ : InMux
    port map (
            O => \N__7688\,
            I => \N__7682\
        );

    \I__1916\ : Span4Mux_v
    port map (
            O => \N__7685\,
            I => \N__7677\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__7682\,
            I => \N__7677\
        );

    \I__1914\ : Span4Mux_v
    port map (
            O => \N__7677\,
            I => \N__7674\
        );

    \I__1913\ : Span4Mux_v
    port map (
            O => \N__7674\,
            I => \N__7671\
        );

    \I__1912\ : Span4Mux_h
    port map (
            O => \N__7671\,
            I => \N__7667\
        );

    \I__1911\ : InMux
    port map (
            O => \N__7670\,
            I => \N__7664\
        );

    \I__1910\ : Sp12to4
    port map (
            O => \N__7667\,
            I => \N__7659\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__7664\,
            I => \N__7659\
        );

    \I__1908\ : Span12Mux_h
    port map (
            O => \N__7659\,
            I => \N__7656\
        );

    \I__1907\ : Odrv12
    port map (
            O => \N__7656\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1906\ : InMux
    port map (
            O => \N__7653\,
            I => \N__7650\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__7650\,
            I => \N__7647\
        );

    \I__1904\ : Span4Mux_v
    port map (
            O => \N__7647\,
            I => \N__7643\
        );

    \I__1903\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7640\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__7643\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__7640\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__1900\ : IoInMux
    port map (
            O => \N__7635\,
            I => \N__7632\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__7632\,
            I => \N__7629\
        );

    \I__1898\ : Span4Mux_s3_v
    port map (
            O => \N__7629\,
            I => \N__7626\
        );

    \I__1897\ : Span4Mux_h
    port map (
            O => \N__7626\,
            I => \N__7623\
        );

    \I__1896\ : Sp12to4
    port map (
            O => \N__7623\,
            I => \N__7620\
        );

    \I__1895\ : Span12Mux_s10_v
    port map (
            O => \N__7620\,
            I => \N__7617\
        );

    \I__1894\ : Span12Mux_h
    port map (
            O => \N__7617\,
            I => \N__7614\
        );

    \I__1893\ : Odrv12
    port map (
            O => \N__7614\,
            I => \un1_D_UM_AMIGA_5\
        );

    \I__1892\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7608\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__7608\,
            I => \N__7605\
        );

    \I__1890\ : Span4Mux_v
    port map (
            O => \N__7605\,
            I => \N__7602\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__7602\,
            I => \N__7598\
        );

    \I__1888\ : InMux
    port map (
            O => \N__7601\,
            I => \N__7595\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__7598\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__7595\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__7590\,
            I => \N__7587\
        );

    \I__1884\ : InMux
    port map (
            O => \N__7587\,
            I => \N__7582\
        );

    \I__1883\ : InMux
    port map (
            O => \N__7586\,
            I => \N__7579\
        );

    \I__1882\ : InMux
    port map (
            O => \N__7585\,
            I => \N__7576\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__7582\,
            I => \N__7573\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__7579\,
            I => \N__7570\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__7576\,
            I => \N__7567\
        );

    \I__1878\ : Span4Mux_h
    port map (
            O => \N__7573\,
            I => \N__7564\
        );

    \I__1877\ : Span4Mux_v
    port map (
            O => \N__7570\,
            I => \N__7561\
        );

    \I__1876\ : Span12Mux_v
    port map (
            O => \N__7567\,
            I => \N__7556\
        );

    \I__1875\ : Sp12to4
    port map (
            O => \N__7564\,
            I => \N__7556\
        );

    \I__1874\ : Sp12to4
    port map (
            O => \N__7561\,
            I => \N__7553\
        );

    \I__1873\ : Span12Mux_v
    port map (
            O => \N__7556\,
            I => \N__7550\
        );

    \I__1872\ : Span12Mux_h
    port map (
            O => \N__7553\,
            I => \N__7547\
        );

    \I__1871\ : Odrv12
    port map (
            O => \N__7550\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1870\ : Odrv12
    port map (
            O => \N__7547\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1869\ : IoInMux
    port map (
            O => \N__7542\,
            I => \N__7539\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__7539\,
            I => \N__7536\
        );

    \I__1867\ : Span12Mux_s7_v
    port map (
            O => \N__7536\,
            I => \N__7533\
        );

    \I__1866\ : Span12Mux_h
    port map (
            O => \N__7533\,
            I => \N__7530\
        );

    \I__1865\ : Odrv12
    port map (
            O => \N__7530\,
            I => \un1_D_UM_AMIGA_4\
        );

    \I__1864\ : InMux
    port map (
            O => \N__7527\,
            I => \N__7524\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__7524\,
            I => \N__7521\
        );

    \I__1862\ : Span4Mux_h
    port map (
            O => \N__7521\,
            I => \N__7518\
        );

    \I__1861\ : Sp12to4
    port map (
            O => \N__7518\,
            I => \N__7515\
        );

    \I__1860\ : Span12Mux_v
    port map (
            O => \N__7515\,
            I => \N__7512\
        );

    \I__1859\ : Span12Mux_h
    port map (
            O => \N__7512\,
            I => \N__7509\
        );

    \I__1858\ : Odrv12
    port map (
            O => \N__7509\,
            I => \D_UU_040_in_5\
        );

    \I__1857\ : IoInMux
    port map (
            O => \N__7506\,
            I => \N__7503\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__7503\,
            I => \N__7500\
        );

    \I__1855\ : IoSpan4Mux
    port map (
            O => \N__7500\,
            I => \N__7497\
        );

    \I__1854\ : IoSpan4Mux
    port map (
            O => \N__7497\,
            I => \N__7494\
        );

    \I__1853\ : Span4Mux_s2_h
    port map (
            O => \N__7494\,
            I => \N__7490\
        );

    \I__1852\ : InMux
    port map (
            O => \N__7493\,
            I => \N__7487\
        );

    \I__1851\ : Sp12to4
    port map (
            O => \N__7490\,
            I => \N__7484\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__7487\,
            I => \N__7481\
        );

    \I__1849\ : Span12Mux_h
    port map (
            O => \N__7484\,
            I => \N__7476\
        );

    \I__1848\ : Span12Mux_v
    port map (
            O => \N__7481\,
            I => \N__7476\
        );

    \I__1847\ : Span12Mux_h
    port map (
            O => \N__7476\,
            I => \N__7473\
        );

    \I__1846\ : Odrv12
    port map (
            O => \N__7473\,
            I => \D_LM_040_in_5\
        );

    \I__1845\ : IoInMux
    port map (
            O => \N__7470\,
            I => \N__7467\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__7467\,
            I => \N__7464\
        );

    \I__1843\ : IoSpan4Mux
    port map (
            O => \N__7464\,
            I => \N__7461\
        );

    \I__1842\ : Span4Mux_s2_h
    port map (
            O => \N__7461\,
            I => \N__7458\
        );

    \I__1841\ : Sp12to4
    port map (
            O => \N__7458\,
            I => \N__7455\
        );

    \I__1840\ : Span12Mux_h
    port map (
            O => \N__7455\,
            I => \N__7452\
        );

    \I__1839\ : Odrv12
    port map (
            O => \N__7452\,
            I => \un1_D_UU_040_5\
        );

    \I__1838\ : InMux
    port map (
            O => \N__7449\,
            I => \N__7446\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__7446\,
            I => \N__7442\
        );

    \I__1836\ : InMux
    port map (
            O => \N__7445\,
            I => \N__7439\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__7442\,
            I => \N__7433\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__7439\,
            I => \N__7433\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__7438\,
            I => \N__7430\
        );

    \I__1832\ : Span4Mux_h
    port map (
            O => \N__7433\,
            I => \N__7427\
        );

    \I__1831\ : InMux
    port map (
            O => \N__7430\,
            I => \N__7424\
        );

    \I__1830\ : Span4Mux_v
    port map (
            O => \N__7427\,
            I => \N__7420\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__7424\,
            I => \N__7417\
        );

    \I__1828\ : InMux
    port map (
            O => \N__7423\,
            I => \N__7414\
        );

    \I__1827\ : Span4Mux_v
    port map (
            O => \N__7420\,
            I => \N__7409\
        );

    \I__1826\ : Span4Mux_h
    port map (
            O => \N__7417\,
            I => \N__7409\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__7414\,
            I => \N__7405\
        );

    \I__1824\ : Span4Mux_v
    port map (
            O => \N__7409\,
            I => \N__7402\
        );

    \I__1823\ : InMux
    port map (
            O => \N__7408\,
            I => \N__7399\
        );

    \I__1822\ : Span12Mux_h
    port map (
            O => \N__7405\,
            I => \N__7396\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__7402\,
            I => \N__7393\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__7399\,
            I => \N__7390\
        );

    \I__1819\ : Span12Mux_v
    port map (
            O => \N__7396\,
            I => \N__7387\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__7393\,
            I => \N__7384\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__7390\,
            I => \N__7381\
        );

    \I__1816\ : Odrv12
    port map (
            O => \N__7387\,
            I => \LBENn_c\
        );

    \I__1815\ : Odrv4
    port map (
            O => \N__7384\,
            I => \LBENn_c\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__7381\,
            I => \LBENn_c\
        );

    \I__1813\ : IoInMux
    port map (
            O => \N__7374\,
            I => \N__7371\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__7371\,
            I => \N__7368\
        );

    \I__1811\ : Odrv12
    port map (
            O => \N__7368\,
            I => \LBENn_c_i\
        );

    \I__1810\ : InMux
    port map (
            O => \N__7365\,
            I => \N__7362\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__7362\,
            I => \N__7359\
        );

    \I__1808\ : Span4Mux_v
    port map (
            O => \N__7359\,
            I => \N__7356\
        );

    \I__1807\ : Sp12to4
    port map (
            O => \N__7356\,
            I => \N__7353\
        );

    \I__1806\ : Span12Mux_h
    port map (
            O => \N__7353\,
            I => \N__7350\
        );

    \I__1805\ : Odrv12
    port map (
            O => \N__7350\,
            I => \D_LL_AMIGA_in_0\
        );

    \I__1804\ : IoInMux
    port map (
            O => \N__7347\,
            I => \N__7344\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__7344\,
            I => \N__7341\
        );

    \I__1802\ : Span4Mux_s2_h
    port map (
            O => \N__7341\,
            I => \N__7338\
        );

    \I__1801\ : Span4Mux_v
    port map (
            O => \N__7338\,
            I => \N__7335\
        );

    \I__1800\ : Span4Mux_h
    port map (
            O => \N__7335\,
            I => \N__7332\
        );

    \I__1799\ : Sp12to4
    port map (
            O => \N__7332\,
            I => \N__7329\
        );

    \I__1798\ : Span12Mux_h
    port map (
            O => \N__7329\,
            I => \N__7326\
        );

    \I__1797\ : Odrv12
    port map (
            O => \N__7326\,
            I => \un2_D_LL_AMIGA_0\
        );

    \I__1796\ : InMux
    port map (
            O => \N__7323\,
            I => \N__7320\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__7320\,
            I => \N__7315\
        );

    \I__1794\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7312\
        );

    \I__1793\ : InMux
    port map (
            O => \N__7318\,
            I => \N__7309\
        );

    \I__1792\ : Odrv12
    port map (
            O => \N__7315\,
            I => \U111_CYCLE_SM.CYCLE_ENZ0\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__7312\,
            I => \U111_CYCLE_SM.CYCLE_ENZ0\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__7309\,
            I => \U111_CYCLE_SM.CYCLE_ENZ0\
        );

    \I__1789\ : InMux
    port map (
            O => \N__7302\,
            I => \N__7298\
        );

    \I__1788\ : InMux
    port map (
            O => \N__7301\,
            I => \N__7295\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__7298\,
            I => \N__7292\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__7295\,
            I => \N__7289\
        );

    \I__1785\ : Span4Mux_v
    port map (
            O => \N__7292\,
            I => \N__7286\
        );

    \I__1784\ : Span4Mux_v
    port map (
            O => \N__7289\,
            I => \N__7283\
        );

    \I__1783\ : Sp12to4
    port map (
            O => \N__7286\,
            I => \N__7278\
        );

    \I__1782\ : Sp12to4
    port map (
            O => \N__7283\,
            I => \N__7278\
        );

    \I__1781\ : Span12Mux_h
    port map (
            O => \N__7278\,
            I => \N__7275\
        );

    \I__1780\ : Odrv12
    port map (
            O => \N__7275\,
            I => \BGn_c\
        );

    \I__1779\ : IoInMux
    port map (
            O => \N__7272\,
            I => \N__7268\
        );

    \I__1778\ : IoInMux
    port map (
            O => \N__7271\,
            I => \N__7265\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__7268\,
            I => \N__7262\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__7265\,
            I => \N__7259\
        );

    \I__1775\ : IoSpan4Mux
    port map (
            O => \N__7262\,
            I => \N__7253\
        );

    \I__1774\ : IoSpan4Mux
    port map (
            O => \N__7259\,
            I => \N__7250\
        );

    \I__1773\ : InMux
    port map (
            O => \N__7258\,
            I => \N__7247\
        );

    \I__1772\ : InMux
    port map (
            O => \N__7257\,
            I => \N__7242\
        );

    \I__1771\ : InMux
    port map (
            O => \N__7256\,
            I => \N__7242\
        );

    \I__1770\ : Span4Mux_s2_h
    port map (
            O => \N__7253\,
            I => \N__7239\
        );

    \I__1769\ : Span4Mux_s1_v
    port map (
            O => \N__7250\,
            I => \N__7236\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__7247\,
            I => \N__7231\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__7242\,
            I => \N__7231\
        );

    \I__1766\ : Sp12to4
    port map (
            O => \N__7239\,
            I => \N__7227\
        );

    \I__1765\ : Span4Mux_v
    port map (
            O => \N__7236\,
            I => \N__7224\
        );

    \I__1764\ : Span4Mux_v
    port map (
            O => \N__7231\,
            I => \N__7221\
        );

    \I__1763\ : InMux
    port map (
            O => \N__7230\,
            I => \N__7218\
        );

    \I__1762\ : Span12Mux_s9_h
    port map (
            O => \N__7227\,
            I => \N__7215\
        );

    \I__1761\ : Span4Mux_v
    port map (
            O => \N__7224\,
            I => \N__7210\
        );

    \I__1760\ : Span4Mux_h
    port map (
            O => \N__7221\,
            I => \N__7210\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__7218\,
            I => \N__7207\
        );

    \I__1758\ : Span12Mux_v
    port map (
            O => \N__7215\,
            I => \N__7204\
        );

    \I__1757\ : Span4Mux_v
    port map (
            O => \N__7210\,
            I => \N__7201\
        );

    \I__1756\ : Span4Mux_h
    port map (
            O => \N__7207\,
            I => \N__7198\
        );

    \I__1755\ : Odrv12
    port map (
            O => \N__7204\,
            I => \CPUBGn_c\
        );

    \I__1754\ : Odrv4
    port map (
            O => \N__7201\,
            I => \CPUBGn_c\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__7198\,
            I => \CPUBGn_c\
        );

    \I__1752\ : InMux
    port map (
            O => \N__7191\,
            I => \N__7185\
        );

    \I__1751\ : InMux
    port map (
            O => \N__7190\,
            I => \N__7178\
        );

    \I__1750\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7178\
        );

    \I__1749\ : InMux
    port map (
            O => \N__7188\,
            I => \N__7178\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__7185\,
            I => \N__7164\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__7178\,
            I => \N__7161\
        );

    \I__1746\ : InMux
    port map (
            O => \N__7177\,
            I => \N__7148\
        );

    \I__1745\ : InMux
    port map (
            O => \N__7176\,
            I => \N__7148\
        );

    \I__1744\ : InMux
    port map (
            O => \N__7175\,
            I => \N__7148\
        );

    \I__1743\ : InMux
    port map (
            O => \N__7174\,
            I => \N__7148\
        );

    \I__1742\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7148\
        );

    \I__1741\ : InMux
    port map (
            O => \N__7172\,
            I => \N__7148\
        );

    \I__1740\ : InMux
    port map (
            O => \N__7171\,
            I => \N__7141\
        );

    \I__1739\ : InMux
    port map (
            O => \N__7170\,
            I => \N__7141\
        );

    \I__1738\ : InMux
    port map (
            O => \N__7169\,
            I => \N__7141\
        );

    \I__1737\ : InMux
    port map (
            O => \N__7168\,
            I => \N__7134\
        );

    \I__1736\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7131\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__7164\,
            I => \N__7128\
        );

    \I__1734\ : Span4Mux_h
    port map (
            O => \N__7161\,
            I => \N__7125\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__7148\,
            I => \N__7122\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__7141\,
            I => \N__7119\
        );

    \I__1731\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7112\
        );

    \I__1730\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7112\
        );

    \I__1729\ : InMux
    port map (
            O => \N__7138\,
            I => \N__7112\
        );

    \I__1728\ : InMux
    port map (
            O => \N__7137\,
            I => \N__7109\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__7134\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__7131\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1725\ : Odrv4
    port map (
            O => \N__7128\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__7125\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__7122\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1722\ : Odrv4
    port map (
            O => \N__7119\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__7112\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__7109\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__7092\,
            I => \CPUBGn_c_cascade_\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__7089\,
            I => \N__7084\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__7088\,
            I => \N__7081\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__7087\,
            I => \N__7078\
        );

    \I__1715\ : InMux
    port map (
            O => \N__7084\,
            I => \N__7075\
        );

    \I__1714\ : InMux
    port map (
            O => \N__7081\,
            I => \N__7072\
        );

    \I__1713\ : InMux
    port map (
            O => \N__7078\,
            I => \N__7069\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__7075\,
            I => \N__7064\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__7072\,
            I => \N__7059\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__7069\,
            I => \N__7059\
        );

    \I__1709\ : InMux
    port map (
            O => \N__7068\,
            I => \N__7056\
        );

    \I__1708\ : InMux
    port map (
            O => \N__7067\,
            I => \N__7053\
        );

    \I__1707\ : Span4Mux_v
    port map (
            O => \N__7064\,
            I => \N__7050\
        );

    \I__1706\ : Span4Mux_h
    port map (
            O => \N__7059\,
            I => \N__7047\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__7056\,
            I => \N__7044\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__7053\,
            I => \N__7041\
        );

    \I__1703\ : Span4Mux_v
    port map (
            O => \N__7050\,
            I => \N__7038\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__7047\,
            I => \N__7035\
        );

    \I__1701\ : Sp12to4
    port map (
            O => \N__7044\,
            I => \N__7032\
        );

    \I__1700\ : Span12Mux_s11_v
    port map (
            O => \N__7041\,
            I => \N__7029\
        );

    \I__1699\ : Sp12to4
    port map (
            O => \N__7038\,
            I => \N__7022\
        );

    \I__1698\ : Sp12to4
    port map (
            O => \N__7035\,
            I => \N__7022\
        );

    \I__1697\ : Span12Mux_v
    port map (
            O => \N__7032\,
            I => \N__7022\
        );

    \I__1696\ : Span12Mux_h
    port map (
            O => \N__7029\,
            I => \N__7019\
        );

    \I__1695\ : Span12Mux_h
    port map (
            O => \N__7022\,
            I => \N__7016\
        );

    \I__1694\ : Odrv12
    port map (
            O => \N__7019\,
            I => \RnW_c\
        );

    \I__1693\ : Odrv12
    port map (
            O => \N__7016\,
            I => \RnW_c\
        );

    \I__1692\ : IoInMux
    port map (
            O => \N__7011\,
            I => \N__7006\
        );

    \I__1691\ : IoInMux
    port map (
            O => \N__7010\,
            I => \N__7001\
        );

    \I__1690\ : IoInMux
    port map (
            O => \N__7009\,
            I => \N__6998\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__7006\,
            I => \N__6991\
        );

    \I__1688\ : IoInMux
    port map (
            O => \N__7005\,
            I => \N__6988\
        );

    \I__1687\ : IoInMux
    port map (
            O => \N__7004\,
            I => \N__6985\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__7001\,
            I => \N__6980\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__6998\,
            I => \N__6980\
        );

    \I__1684\ : IoInMux
    port map (
            O => \N__6997\,
            I => \N__6977\
        );

    \I__1683\ : IoInMux
    port map (
            O => \N__6996\,
            I => \N__6974\
        );

    \I__1682\ : IoInMux
    port map (
            O => \N__6995\,
            I => \N__6966\
        );

    \I__1681\ : IoInMux
    port map (
            O => \N__6994\,
            I => \N__6963\
        );

    \I__1680\ : IoSpan4Mux
    port map (
            O => \N__6991\,
            I => \N__6953\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__6988\,
            I => \N__6953\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__6985\,
            I => \N__6953\
        );

    \I__1677\ : Span4Mux_s2_h
    port map (
            O => \N__6980\,
            I => \N__6946\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__6977\,
            I => \N__6946\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__6974\,
            I => \N__6946\
        );

    \I__1674\ : IoInMux
    port map (
            O => \N__6973\,
            I => \N__6943\
        );

    \I__1673\ : IoInMux
    port map (
            O => \N__6972\,
            I => \N__6940\
        );

    \I__1672\ : IoInMux
    port map (
            O => \N__6971\,
            I => \N__6937\
        );

    \I__1671\ : IoInMux
    port map (
            O => \N__6970\,
            I => \N__6933\
        );

    \I__1670\ : IoInMux
    port map (
            O => \N__6969\,
            I => \N__6928\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__6966\,
            I => \N__6919\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__6963\,
            I => \N__6919\
        );

    \I__1667\ : IoInMux
    port map (
            O => \N__6962\,
            I => \N__6916\
        );

    \I__1666\ : IoInMux
    port map (
            O => \N__6961\,
            I => \N__6913\
        );

    \I__1665\ : IoInMux
    port map (
            O => \N__6960\,
            I => \N__6910\
        );

    \I__1664\ : IoSpan4Mux
    port map (
            O => \N__6953\,
            I => \N__6897\
        );

    \I__1663\ : IoSpan4Mux
    port map (
            O => \N__6946\,
            I => \N__6897\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__6943\,
            I => \N__6897\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__6940\,
            I => \N__6897\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__6937\,
            I => \N__6897\
        );

    \I__1659\ : IoInMux
    port map (
            O => \N__6936\,
            I => \N__6894\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__6933\,
            I => \N__6891\
        );

    \I__1657\ : IoInMux
    port map (
            O => \N__6932\,
            I => \N__6888\
        );

    \I__1656\ : IoInMux
    port map (
            O => \N__6931\,
            I => \N__6885\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__6928\,
            I => \N__6882\
        );

    \I__1654\ : IoInMux
    port map (
            O => \N__6927\,
            I => \N__6879\
        );

    \I__1653\ : IoInMux
    port map (
            O => \N__6926\,
            I => \N__6876\
        );

    \I__1652\ : IoInMux
    port map (
            O => \N__6925\,
            I => \N__6873\
        );

    \I__1651\ : IoInMux
    port map (
            O => \N__6924\,
            I => \N__6870\
        );

    \I__1650\ : IoSpan4Mux
    port map (
            O => \N__6919\,
            I => \N__6861\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__6916\,
            I => \N__6861\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__6913\,
            I => \N__6861\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__6910\,
            I => \N__6861\
        );

    \I__1646\ : IoInMux
    port map (
            O => \N__6909\,
            I => \N__6856\
        );

    \I__1645\ : IoInMux
    port map (
            O => \N__6908\,
            I => \N__6853\
        );

    \I__1644\ : IoSpan4Mux
    port map (
            O => \N__6897\,
            I => \N__6844\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__6894\,
            I => \N__6844\
        );

    \I__1642\ : IoSpan4Mux
    port map (
            O => \N__6891\,
            I => \N__6837\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__6888\,
            I => \N__6837\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__6885\,
            I => \N__6837\
        );

    \I__1639\ : IoSpan4Mux
    port map (
            O => \N__6882\,
            I => \N__6826\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__6879\,
            I => \N__6826\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__6876\,
            I => \N__6826\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__6873\,
            I => \N__6826\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__6870\,
            I => \N__6826\
        );

    \I__1634\ : IoSpan4Mux
    port map (
            O => \N__6861\,
            I => \N__6823\
        );

    \I__1633\ : IoInMux
    port map (
            O => \N__6860\,
            I => \N__6820\
        );

    \I__1632\ : IoInMux
    port map (
            O => \N__6859\,
            I => \N__6817\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__6856\,
            I => \N__6812\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__6853\,
            I => \N__6812\
        );

    \I__1629\ : IoInMux
    port map (
            O => \N__6852\,
            I => \N__6809\
        );

    \I__1628\ : IoInMux
    port map (
            O => \N__6851\,
            I => \N__6806\
        );

    \I__1627\ : IoInMux
    port map (
            O => \N__6850\,
            I => \N__6803\
        );

    \I__1626\ : IoInMux
    port map (
            O => \N__6849\,
            I => \N__6800\
        );

    \I__1625\ : Span4Mux_s2_v
    port map (
            O => \N__6844\,
            I => \N__6797\
        );

    \I__1624\ : IoSpan4Mux
    port map (
            O => \N__6837\,
            I => \N__6792\
        );

    \I__1623\ : IoSpan4Mux
    port map (
            O => \N__6826\,
            I => \N__6792\
        );

    \I__1622\ : Span4Mux_s3_h
    port map (
            O => \N__6823\,
            I => \N__6789\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__6820\,
            I => \N__6784\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__6817\,
            I => \N__6784\
        );

    \I__1619\ : Span12Mux_s5_h
    port map (
            O => \N__6812\,
            I => \N__6781\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__6809\,
            I => \N__6778\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__6806\,
            I => \N__6773\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__6803\,
            I => \N__6773\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__6800\,
            I => \N__6770\
        );

    \I__1614\ : Span4Mux_h
    port map (
            O => \N__6797\,
            I => \N__6767\
        );

    \I__1613\ : Span4Mux_s2_h
    port map (
            O => \N__6792\,
            I => \N__6764\
        );

    \I__1612\ : Sp12to4
    port map (
            O => \N__6789\,
            I => \N__6759\
        );

    \I__1611\ : Span12Mux_s5_h
    port map (
            O => \N__6784\,
            I => \N__6759\
        );

    \I__1610\ : Span12Mux_h
    port map (
            O => \N__6781\,
            I => \N__6756\
        );

    \I__1609\ : Span12Mux_s6_v
    port map (
            O => \N__6778\,
            I => \N__6753\
        );

    \I__1608\ : Span12Mux_s10_h
    port map (
            O => \N__6773\,
            I => \N__6750\
        );

    \I__1607\ : Span12Mux_s10_h
    port map (
            O => \N__6770\,
            I => \N__6745\
        );

    \I__1606\ : Sp12to4
    port map (
            O => \N__6767\,
            I => \N__6745\
        );

    \I__1605\ : Sp12to4
    port map (
            O => \N__6764\,
            I => \N__6742\
        );

    \I__1604\ : Span12Mux_h
    port map (
            O => \N__6759\,
            I => \N__6739\
        );

    \I__1603\ : Span12Mux_v
    port map (
            O => \N__6756\,
            I => \N__6734\
        );

    \I__1602\ : Span12Mux_h
    port map (
            O => \N__6753\,
            I => \N__6734\
        );

    \I__1601\ : Span12Mux_v
    port map (
            O => \N__6750\,
            I => \N__6727\
        );

    \I__1600\ : Span12Mux_v
    port map (
            O => \N__6745\,
            I => \N__6727\
        );

    \I__1599\ : Span12Mux_s10_h
    port map (
            O => \N__6742\,
            I => \N__6727\
        );

    \I__1598\ : Odrv12
    port map (
            O => \N__6739\,
            I => \N_62_i\
        );

    \I__1597\ : Odrv12
    port map (
            O => \N__6734\,
            I => \N_62_i\
        );

    \I__1596\ : Odrv12
    port map (
            O => \N__6727\,
            I => \N_62_i\
        );

    \I__1595\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6717\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__6717\,
            I => \N__6714\
        );

    \I__1593\ : Span4Mux_v
    port map (
            O => \N__6714\,
            I => \N__6709\
        );

    \I__1592\ : InMux
    port map (
            O => \N__6713\,
            I => \N__6706\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__6712\,
            I => \N__6703\
        );

    \I__1590\ : Span4Mux_v
    port map (
            O => \N__6709\,
            I => \N__6700\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__6706\,
            I => \N__6697\
        );

    \I__1588\ : InMux
    port map (
            O => \N__6703\,
            I => \N__6694\
        );

    \I__1587\ : Span4Mux_v
    port map (
            O => \N__6700\,
            I => \N__6689\
        );

    \I__1586\ : Span4Mux_v
    port map (
            O => \N__6697\,
            I => \N__6689\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__6694\,
            I => \N__6686\
        );

    \I__1584\ : Sp12to4
    port map (
            O => \N__6689\,
            I => \N__6681\
        );

    \I__1583\ : Span12Mux_v
    port map (
            O => \N__6686\,
            I => \N__6681\
        );

    \I__1582\ : Span12Mux_h
    port map (
            O => \N__6681\,
            I => \N__6678\
        );

    \I__1581\ : Odrv12
    port map (
            O => \N__6678\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1580\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6671\
        );

    \I__1579\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6668\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__6671\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__6668\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__1576\ : IoInMux
    port map (
            O => \N__6663\,
            I => \N__6660\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__6660\,
            I => \N__6657\
        );

    \I__1574\ : IoSpan4Mux
    port map (
            O => \N__6657\,
            I => \N__6654\
        );

    \I__1573\ : Span4Mux_s0_h
    port map (
            O => \N__6654\,
            I => \N__6651\
        );

    \I__1572\ : Span4Mux_h
    port map (
            O => \N__6651\,
            I => \N__6648\
        );

    \I__1571\ : Sp12to4
    port map (
            O => \N__6648\,
            I => \N__6645\
        );

    \I__1570\ : Odrv12
    port map (
            O => \N__6645\,
            I => \un1_D_UM_AMIGA_2\
        );

    \I__1569\ : InMux
    port map (
            O => \N__6642\,
            I => \N__6636\
        );

    \I__1568\ : InMux
    port map (
            O => \N__6641\,
            I => \N__6636\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__6636\,
            I => \N__6632\
        );

    \I__1566\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6629\
        );

    \I__1565\ : Span4Mux_v
    port map (
            O => \N__6632\,
            I => \N__6621\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__6629\,
            I => \N__6621\
        );

    \I__1563\ : InMux
    port map (
            O => \N__6628\,
            I => \N__6618\
        );

    \I__1562\ : InMux
    port map (
            O => \N__6627\,
            I => \N__6613\
        );

    \I__1561\ : InMux
    port map (
            O => \N__6626\,
            I => \N__6613\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__6621\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__6618\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__6613\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1557\ : InMux
    port map (
            O => \N__6606\,
            I => \N__6597\
        );

    \I__1556\ : InMux
    port map (
            O => \N__6605\,
            I => \N__6585\
        );

    \I__1555\ : InMux
    port map (
            O => \N__6604\,
            I => \N__6580\
        );

    \I__1554\ : InMux
    port map (
            O => \N__6603\,
            I => \N__6580\
        );

    \I__1553\ : InMux
    port map (
            O => \N__6602\,
            I => \N__6577\
        );

    \I__1552\ : InMux
    port map (
            O => \N__6601\,
            I => \N__6572\
        );

    \I__1551\ : InMux
    port map (
            O => \N__6600\,
            I => \N__6572\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__6597\,
            I => \N__6569\
        );

    \I__1549\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6556\
        );

    \I__1548\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6556\
        );

    \I__1547\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6556\
        );

    \I__1546\ : InMux
    port map (
            O => \N__6593\,
            I => \N__6556\
        );

    \I__1545\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6556\
        );

    \I__1544\ : InMux
    port map (
            O => \N__6591\,
            I => \N__6556\
        );

    \I__1543\ : InMux
    port map (
            O => \N__6590\,
            I => \N__6549\
        );

    \I__1542\ : InMux
    port map (
            O => \N__6589\,
            I => \N__6549\
        );

    \I__1541\ : InMux
    port map (
            O => \N__6588\,
            I => \N__6549\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__6585\,
            I => \U111_CYCLE_SM.N_107_i\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__6580\,
            I => \U111_CYCLE_SM.N_107_i\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__6577\,
            I => \U111_CYCLE_SM.N_107_i\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__6572\,
            I => \U111_CYCLE_SM.N_107_i\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__6569\,
            I => \U111_CYCLE_SM.N_107_i\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__6556\,
            I => \U111_CYCLE_SM.N_107_i\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__6549\,
            I => \U111_CYCLE_SM.N_107_i\
        );

    \I__1533\ : InMux
    port map (
            O => \N__6534\,
            I => \N__6530\
        );

    \I__1532\ : InMux
    port map (
            O => \N__6533\,
            I => \N__6527\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__6530\,
            I => \N__6524\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__6527\,
            I => \N__6521\
        );

    \I__1529\ : Span12Mux_h
    port map (
            O => \N__6524\,
            I => \N__6518\
        );

    \I__1528\ : Sp12to4
    port map (
            O => \N__6521\,
            I => \N__6515\
        );

    \I__1527\ : Span12Mux_h
    port map (
            O => \N__6518\,
            I => \N__6512\
        );

    \I__1526\ : Span12Mux_v
    port map (
            O => \N__6515\,
            I => \N__6509\
        );

    \I__1525\ : Span12Mux_v
    port map (
            O => \N__6512\,
            I => \N__6506\
        );

    \I__1524\ : Span12Mux_h
    port map (
            O => \N__6509\,
            I => \N__6503\
        );

    \I__1523\ : Odrv12
    port map (
            O => \N__6506\,
            I => \SIZ_c_1\
        );

    \I__1522\ : Odrv12
    port map (
            O => \N__6503\,
            I => \SIZ_c_1\
        );

    \I__1521\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6494\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__6497\,
            I => \N__6491\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__6494\,
            I => \N__6488\
        );

    \I__1518\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6485\
        );

    \I__1517\ : Span4Mux_h
    port map (
            O => \N__6488\,
            I => \N__6480\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__6485\,
            I => \N__6480\
        );

    \I__1515\ : Span4Mux_v
    port map (
            O => \N__6480\,
            I => \N__6477\
        );

    \I__1514\ : Span4Mux_v
    port map (
            O => \N__6477\,
            I => \N__6474\
        );

    \I__1513\ : Sp12to4
    port map (
            O => \N__6474\,
            I => \N__6471\
        );

    \I__1512\ : Span12Mux_h
    port map (
            O => \N__6471\,
            I => \N__6468\
        );

    \I__1511\ : Odrv12
    port map (
            O => \N__6468\,
            I => \SIZ_c_0\
        );

    \I__1510\ : CascadeMux
    port map (
            O => \N__6465\,
            I => \N__6459\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__6464\,
            I => \N__6454\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__6463\,
            I => \N__6450\
        );

    \I__1507\ : InMux
    port map (
            O => \N__6462\,
            I => \N__6447\
        );

    \I__1506\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6444\
        );

    \I__1505\ : InMux
    port map (
            O => \N__6458\,
            I => \N__6441\
        );

    \I__1504\ : InMux
    port map (
            O => \N__6457\,
            I => \N__6438\
        );

    \I__1503\ : InMux
    port map (
            O => \N__6454\,
            I => \N__6433\
        );

    \I__1502\ : InMux
    port map (
            O => \N__6453\,
            I => \N__6433\
        );

    \I__1501\ : InMux
    port map (
            O => \N__6450\,
            I => \N__6430\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__6447\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__6444\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__6441\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__6438\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__6433\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__6430\,
            I => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\
        );

    \I__1494\ : InMux
    port map (
            O => \N__6417\,
            I => \N__6414\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__6414\,
            I => \N__6410\
        );

    \I__1492\ : InMux
    port map (
            O => \N__6413\,
            I => \N__6406\
        );

    \I__1491\ : Span4Mux_h
    port map (
            O => \N__6410\,
            I => \N__6403\
        );

    \I__1490\ : InMux
    port map (
            O => \N__6409\,
            I => \N__6400\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__6406\,
            I => \N__6397\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__6403\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__6400\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__6397\,
            I => \U111_CYCLE_SM.LW_TRANSZ0\
        );

    \I__1485\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6387\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__6387\,
            I => \N__6371\
        );

    \I__1483\ : ClkMux
    port map (
            O => \N__6386\,
            I => \N__6342\
        );

    \I__1482\ : ClkMux
    port map (
            O => \N__6385\,
            I => \N__6342\
        );

    \I__1481\ : ClkMux
    port map (
            O => \N__6384\,
            I => \N__6342\
        );

    \I__1480\ : ClkMux
    port map (
            O => \N__6383\,
            I => \N__6342\
        );

    \I__1479\ : ClkMux
    port map (
            O => \N__6382\,
            I => \N__6342\
        );

    \I__1478\ : ClkMux
    port map (
            O => \N__6381\,
            I => \N__6342\
        );

    \I__1477\ : ClkMux
    port map (
            O => \N__6380\,
            I => \N__6342\
        );

    \I__1476\ : ClkMux
    port map (
            O => \N__6379\,
            I => \N__6342\
        );

    \I__1475\ : ClkMux
    port map (
            O => \N__6378\,
            I => \N__6342\
        );

    \I__1474\ : ClkMux
    port map (
            O => \N__6377\,
            I => \N__6342\
        );

    \I__1473\ : ClkMux
    port map (
            O => \N__6376\,
            I => \N__6342\
        );

    \I__1472\ : ClkMux
    port map (
            O => \N__6375\,
            I => \N__6342\
        );

    \I__1471\ : ClkMux
    port map (
            O => \N__6374\,
            I => \N__6342\
        );

    \I__1470\ : Glb2LocalMux
    port map (
            O => \N__6371\,
            I => \N__6342\
        );

    \I__1469\ : GlobalMux
    port map (
            O => \N__6342\,
            I => \CLK40\
        );

    \I__1468\ : SRMux
    port map (
            O => \N__6339\,
            I => \N__6312\
        );

    \I__1467\ : SRMux
    port map (
            O => \N__6338\,
            I => \N__6312\
        );

    \I__1466\ : SRMux
    port map (
            O => \N__6337\,
            I => \N__6312\
        );

    \I__1465\ : SRMux
    port map (
            O => \N__6336\,
            I => \N__6312\
        );

    \I__1464\ : SRMux
    port map (
            O => \N__6335\,
            I => \N__6312\
        );

    \I__1463\ : SRMux
    port map (
            O => \N__6334\,
            I => \N__6312\
        );

    \I__1462\ : SRMux
    port map (
            O => \N__6333\,
            I => \N__6312\
        );

    \I__1461\ : SRMux
    port map (
            O => \N__6332\,
            I => \N__6312\
        );

    \I__1460\ : SRMux
    port map (
            O => \N__6331\,
            I => \N__6312\
        );

    \I__1459\ : GlobalMux
    port map (
            O => \N__6312\,
            I => \N__6309\
        );

    \I__1458\ : gio2CtrlBuf
    port map (
            O => \N__6309\,
            I => \RESETn_c_i_g\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__6306\,
            I => \N__6303\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6303\,
            I => \N__6300\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__6300\,
            I => \N__6296\
        );

    \I__1454\ : InMux
    port map (
            O => \N__6299\,
            I => \N__6293\
        );

    \I__1453\ : Span4Mux_v
    port map (
            O => \N__6296\,
            I => \N__6289\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__6293\,
            I => \N__6286\
        );

    \I__1451\ : InMux
    port map (
            O => \N__6292\,
            I => \N__6283\
        );

    \I__1450\ : Span4Mux_h
    port map (
            O => \N__6289\,
            I => \N__6278\
        );

    \I__1449\ : Span4Mux_v
    port map (
            O => \N__6286\,
            I => \N__6278\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__6283\,
            I => \N__6275\
        );

    \I__1447\ : Span4Mux_v
    port map (
            O => \N__6278\,
            I => \N__6272\
        );

    \I__1446\ : Span4Mux_v
    port map (
            O => \N__6275\,
            I => \N__6269\
        );

    \I__1445\ : Span4Mux_v
    port map (
            O => \N__6272\,
            I => \N__6264\
        );

    \I__1444\ : Span4Mux_h
    port map (
            O => \N__6269\,
            I => \N__6264\
        );

    \I__1443\ : Sp12to4
    port map (
            O => \N__6264\,
            I => \N__6261\
        );

    \I__1442\ : Odrv12
    port map (
            O => \N__6261\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__1441\ : InMux
    port map (
            O => \N__6258\,
            I => \N__6255\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__6255\,
            I => \N__6251\
        );

    \I__1439\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6248\
        );

    \I__1438\ : Odrv12
    port map (
            O => \N__6251\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__6248\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__1436\ : IoInMux
    port map (
            O => \N__6243\,
            I => \N__6240\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__6240\,
            I => \N__6237\
        );

    \I__1434\ : IoSpan4Mux
    port map (
            O => \N__6237\,
            I => \N__6234\
        );

    \I__1433\ : Span4Mux_s1_h
    port map (
            O => \N__6234\,
            I => \N__6231\
        );

    \I__1432\ : Span4Mux_v
    port map (
            O => \N__6231\,
            I => \N__6228\
        );

    \I__1431\ : Sp12to4
    port map (
            O => \N__6228\,
            I => \N__6225\
        );

    \I__1430\ : Span12Mux_s10_h
    port map (
            O => \N__6225\,
            I => \N__6222\
        );

    \I__1429\ : Odrv12
    port map (
            O => \N__6222\,
            I => \N_130\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6219\,
            I => \N__6216\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__6216\,
            I => \N__6212\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6209\
        );

    \I__1425\ : Odrv12
    port map (
            O => \N__6212\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__6209\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1423\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6201\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__6201\,
            I => \N__6197\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__6200\,
            I => \N__6194\
        );

    \I__1420\ : Span4Mux_v
    port map (
            O => \N__6197\,
            I => \N__6191\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6188\
        );

    \I__1418\ : Span4Mux_h
    port map (
            O => \N__6191\,
            I => \N__6183\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6188\,
            I => \N__6183\
        );

    \I__1416\ : Span4Mux_v
    port map (
            O => \N__6183\,
            I => \N__6179\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6176\
        );

    \I__1414\ : Span4Mux_v
    port map (
            O => \N__6179\,
            I => \N__6171\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__6176\,
            I => \N__6171\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__6171\,
            I => \N__6168\
        );

    \I__1411\ : Sp12to4
    port map (
            O => \N__6168\,
            I => \N__6165\
        );

    \I__1410\ : Span12Mux_h
    port map (
            O => \N__6165\,
            I => \N__6162\
        );

    \I__1409\ : Odrv12
    port map (
            O => \N__6162\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1408\ : IoInMux
    port map (
            O => \N__6159\,
            I => \N__6156\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__6156\,
            I => \N__6153\
        );

    \I__1406\ : Span4Mux_s3_v
    port map (
            O => \N__6153\,
            I => \N__6150\
        );

    \I__1405\ : Span4Mux_v
    port map (
            O => \N__6150\,
            I => \N__6147\
        );

    \I__1404\ : Sp12to4
    port map (
            O => \N__6147\,
            I => \N__6144\
        );

    \I__1403\ : Span12Mux_h
    port map (
            O => \N__6144\,
            I => \N__6141\
        );

    \I__1402\ : Odrv12
    port map (
            O => \N__6141\,
            I => \N_131\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6138\,
            I => \N__6134\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6137\,
            I => \N__6131\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6134\,
            I => \N__6127\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6131\,
            I => \N__6124\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__6130\,
            I => \N__6121\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__6127\,
            I => \N__6118\
        );

    \I__1395\ : Span4Mux_v
    port map (
            O => \N__6124\,
            I => \N__6115\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6121\,
            I => \N__6112\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__6118\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__6115\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6112\,
            I => \U111_CYCLE_SM.TA_DISZ0\
        );

    \I__1390\ : IoInMux
    port map (
            O => \N__6105\,
            I => \N__6102\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__6102\,
            I => \N__6099\
        );

    \I__1388\ : IoSpan4Mux
    port map (
            O => \N__6099\,
            I => \N__6096\
        );

    \I__1387\ : Span4Mux_s0_v
    port map (
            O => \N__6096\,
            I => \N__6093\
        );

    \I__1386\ : Span4Mux_v
    port map (
            O => \N__6093\,
            I => \N__6090\
        );

    \I__1385\ : Span4Mux_v
    port map (
            O => \N__6090\,
            I => \N__6087\
        );

    \I__1384\ : Odrv4
    port map (
            O => \N__6087\,
            I => \N_66\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__6084\,
            I => \N__6081\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6077\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6080\,
            I => \N__6074\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__6077\,
            I => \N__6071\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6074\,
            I => \N__6067\
        );

    \I__1378\ : Span4Mux_v
    port map (
            O => \N__6071\,
            I => \N__6064\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6070\,
            I => \N__6061\
        );

    \I__1376\ : Span4Mux_h
    port map (
            O => \N__6067\,
            I => \N__6058\
        );

    \I__1375\ : Span4Mux_v
    port map (
            O => \N__6064\,
            I => \N__6053\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__6061\,
            I => \N__6053\
        );

    \I__1373\ : Span4Mux_v
    port map (
            O => \N__6058\,
            I => \N__6050\
        );

    \I__1372\ : Span4Mux_v
    port map (
            O => \N__6053\,
            I => \N__6047\
        );

    \I__1371\ : Sp12to4
    port map (
            O => \N__6050\,
            I => \N__6044\
        );

    \I__1370\ : Span4Mux_h
    port map (
            O => \N__6047\,
            I => \N__6041\
        );

    \I__1369\ : Span12Mux_v
    port map (
            O => \N__6044\,
            I => \N__6036\
        );

    \I__1368\ : Sp12to4
    port map (
            O => \N__6041\,
            I => \N__6036\
        );

    \I__1367\ : Odrv12
    port map (
            O => \N__6036\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6033\,
            I => \N__6030\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__6030\,
            I => \N__6027\
        );

    \I__1364\ : Span4Mux_v
    port map (
            O => \N__6027\,
            I => \N__6023\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6026\,
            I => \N__6020\
        );

    \I__1362\ : Odrv4
    port map (
            O => \N__6023\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6020\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__1360\ : IoInMux
    port map (
            O => \N__6015\,
            I => \N__6012\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__6012\,
            I => \N__6009\
        );

    \I__1358\ : Span12Mux_s7_h
    port map (
            O => \N__6009\,
            I => \N__6006\
        );

    \I__1357\ : Span12Mux_h
    port map (
            O => \N__6006\,
            I => \N__6003\
        );

    \I__1356\ : Odrv12
    port map (
            O => \N__6003\,
            I => \un1_D_UM_AMIGA_3\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6000\,
            I => \N__5996\
        );

    \I__1354\ : IoInMux
    port map (
            O => \N__5999\,
            I => \N__5993\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__5996\,
            I => \N__5990\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__5993\,
            I => \N__5987\
        );

    \I__1351\ : Span4Mux_v
    port map (
            O => \N__5990\,
            I => \N__5984\
        );

    \I__1350\ : Span4Mux_s2_h
    port map (
            O => \N__5987\,
            I => \N__5981\
        );

    \I__1349\ : Sp12to4
    port map (
            O => \N__5984\,
            I => \N__5978\
        );

    \I__1348\ : Span4Mux_v
    port map (
            O => \N__5981\,
            I => \N__5975\
        );

    \I__1347\ : Span12Mux_v
    port map (
            O => \N__5978\,
            I => \N__5972\
        );

    \I__1346\ : Sp12to4
    port map (
            O => \N__5975\,
            I => \N__5969\
        );

    \I__1345\ : Span12Mux_v
    port map (
            O => \N__5972\,
            I => \N__5964\
        );

    \I__1344\ : Span12Mux_h
    port map (
            O => \N__5969\,
            I => \N__5964\
        );

    \I__1343\ : Span12Mux_h
    port map (
            O => \N__5964\,
            I => \N__5961\
        );

    \I__1342\ : Odrv12
    port map (
            O => \N__5961\,
            I => \D_LL_040_in_4\
        );

    \I__1341\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5955\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__5955\,
            I => \N__5952\
        );

    \I__1339\ : Span4Mux_v
    port map (
            O => \N__5952\,
            I => \N__5949\
        );

    \I__1338\ : Span4Mux_h
    port map (
            O => \N__5949\,
            I => \N__5946\
        );

    \I__1337\ : Sp12to4
    port map (
            O => \N__5946\,
            I => \N__5943\
        );

    \I__1336\ : Span12Mux_h
    port map (
            O => \N__5943\,
            I => \N__5940\
        );

    \I__1335\ : Odrv12
    port map (
            O => \N__5940\,
            I => \D_UM_040_in_4\
        );

    \I__1334\ : IoInMux
    port map (
            O => \N__5937\,
            I => \N__5934\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__5934\,
            I => \N__5931\
        );

    \I__1332\ : IoSpan4Mux
    port map (
            O => \N__5931\,
            I => \N__5928\
        );

    \I__1331\ : Sp12to4
    port map (
            O => \N__5928\,
            I => \N__5925\
        );

    \I__1330\ : Span12Mux_h
    port map (
            O => \N__5925\,
            I => \N__5922\
        );

    \I__1329\ : Odrv12
    port map (
            O => \N__5922\,
            I => \un1_D_UM_040_4\
        );

    \I__1328\ : InMux
    port map (
            O => \N__5919\,
            I => \N__5916\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__5916\,
            I => \N__5913\
        );

    \I__1326\ : Span4Mux_v
    port map (
            O => \N__5913\,
            I => \N__5910\
        );

    \I__1325\ : Sp12to4
    port map (
            O => \N__5910\,
            I => \N__5907\
        );

    \I__1324\ : Span12Mux_h
    port map (
            O => \N__5907\,
            I => \N__5904\
        );

    \I__1323\ : Odrv12
    port map (
            O => \N__5904\,
            I => \D_LL_AMIGA_in_6\
        );

    \I__1322\ : IoInMux
    port map (
            O => \N__5901\,
            I => \N__5898\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__5898\,
            I => \N__5895\
        );

    \I__1320\ : Span4Mux_s2_h
    port map (
            O => \N__5895\,
            I => \N__5892\
        );

    \I__1319\ : Span4Mux_h
    port map (
            O => \N__5892\,
            I => \N__5889\
        );

    \I__1318\ : Sp12to4
    port map (
            O => \N__5889\,
            I => \N__5886\
        );

    \I__1317\ : Span12Mux_s10_v
    port map (
            O => \N__5886\,
            I => \N__5883\
        );

    \I__1316\ : Span12Mux_h
    port map (
            O => \N__5883\,
            I => \N__5880\
        );

    \I__1315\ : Odrv12
    port map (
            O => \N__5880\,
            I => \un2_D_LL_AMIGA_6\
        );

    \I__1314\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5874\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5874\,
            I => \N__5871\
        );

    \I__1312\ : Span12Mux_v
    port map (
            O => \N__5871\,
            I => \N__5868\
        );

    \I__1311\ : Span12Mux_h
    port map (
            O => \N__5868\,
            I => \N__5865\
        );

    \I__1310\ : Odrv12
    port map (
            O => \N__5865\,
            I => \D_LL_AMIGA_in_5\
        );

    \I__1309\ : IoInMux
    port map (
            O => \N__5862\,
            I => \N__5859\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__5859\,
            I => \N__5856\
        );

    \I__1307\ : Span4Mux_s3_h
    port map (
            O => \N__5856\,
            I => \N__5853\
        );

    \I__1306\ : Span4Mux_v
    port map (
            O => \N__5853\,
            I => \N__5850\
        );

    \I__1305\ : Span4Mux_v
    port map (
            O => \N__5850\,
            I => \N__5847\
        );

    \I__1304\ : Span4Mux_h
    port map (
            O => \N__5847\,
            I => \N__5844\
        );

    \I__1303\ : Sp12to4
    port map (
            O => \N__5844\,
            I => \N__5841\
        );

    \I__1302\ : Odrv12
    port map (
            O => \N__5841\,
            I => \un2_D_LL_AMIGA_5\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5835\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__5835\,
            I => \N__5832\
        );

    \I__1299\ : Span4Mux_v
    port map (
            O => \N__5832\,
            I => \N__5829\
        );

    \I__1298\ : Span4Mux_h
    port map (
            O => \N__5829\,
            I => \N__5826\
        );

    \I__1297\ : Sp12to4
    port map (
            O => \N__5826\,
            I => \N__5823\
        );

    \I__1296\ : Span12Mux_v
    port map (
            O => \N__5823\,
            I => \N__5820\
        );

    \I__1295\ : Odrv12
    port map (
            O => \N__5820\,
            I => \TS_CPUn_in\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__5817\,
            I => \N__5813\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5810\
        );

    \I__1292\ : InMux
    port map (
            O => \N__5813\,
            I => \N__5807\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5810\,
            I => \U111_CYCLE_SM.TS_DELAYZ0\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__5807\,
            I => \U111_CYCLE_SM.TS_DELAYZ0\
        );

    \I__1289\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5797\
        );

    \I__1288\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5794\
        );

    \I__1287\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5791\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__5797\,
            I => \U111_CYCLE_SM.un4_TS_OUT_i_0\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__5794\,
            I => \U111_CYCLE_SM.un4_TS_OUT_i_0\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__5791\,
            I => \U111_CYCLE_SM.un4_TS_OUT_i_0\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5780\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5777\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__5780\,
            I => \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__5777\,
            I => \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0\
        );

    \I__1279\ : IoInMux
    port map (
            O => \N__5772\,
            I => \N__5769\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5769\,
            I => \N__5765\
        );

    \I__1277\ : IoInMux
    port map (
            O => \N__5768\,
            I => \N__5761\
        );

    \I__1276\ : IoSpan4Mux
    port map (
            O => \N__5765\,
            I => \N__5758\
        );

    \I__1275\ : IoInMux
    port map (
            O => \N__5764\,
            I => \N__5755\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5761\,
            I => \N__5751\
        );

    \I__1273\ : IoSpan4Mux
    port map (
            O => \N__5758\,
            I => \N__5746\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__5755\,
            I => \N__5746\
        );

    \I__1271\ : IoInMux
    port map (
            O => \N__5754\,
            I => \N__5743\
        );

    \I__1270\ : IoSpan4Mux
    port map (
            O => \N__5751\,
            I => \N__5740\
        );

    \I__1269\ : IoSpan4Mux
    port map (
            O => \N__5746\,
            I => \N__5737\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__5743\,
            I => \N__5734\
        );

    \I__1267\ : Sp12to4
    port map (
            O => \N__5740\,
            I => \N__5731\
        );

    \I__1266\ : Span4Mux_s0_v
    port map (
            O => \N__5737\,
            I => \N__5728\
        );

    \I__1265\ : Span4Mux_s1_h
    port map (
            O => \N__5734\,
            I => \N__5725\
        );

    \I__1264\ : Span12Mux_s7_h
    port map (
            O => \N__5731\,
            I => \N__5722\
        );

    \I__1263\ : Sp12to4
    port map (
            O => \N__5728\,
            I => \N__5719\
        );

    \I__1262\ : Sp12to4
    port map (
            O => \N__5725\,
            I => \N__5716\
        );

    \I__1261\ : Span12Mux_h
    port map (
            O => \N__5722\,
            I => \N__5711\
        );

    \I__1260\ : Span12Mux_v
    port map (
            O => \N__5719\,
            I => \N__5711\
        );

    \I__1259\ : Span12Mux_v
    port map (
            O => \N__5716\,
            I => \N__5708\
        );

    \I__1258\ : Odrv12
    port map (
            O => \N__5711\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__1257\ : Odrv12
    port map (
            O => \N__5708\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5700\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5700\,
            I => \N__5696\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5693\
        );

    \I__1253\ : Odrv12
    port map (
            O => \N__5696\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__5693\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__5688\,
            I => \N__5685\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5685\,
            I => \N__5682\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5682\,
            I => \N__5678\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5681\,
            I => \N__5675\
        );

    \I__1247\ : Span4Mux_v
    port map (
            O => \N__5678\,
            I => \N__5672\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__5675\,
            I => \N__5669\
        );

    \I__1245\ : Span4Mux_v
    port map (
            O => \N__5672\,
            I => \N__5663\
        );

    \I__1244\ : Span4Mux_v
    port map (
            O => \N__5669\,
            I => \N__5663\
        );

    \I__1243\ : InMux
    port map (
            O => \N__5668\,
            I => \N__5660\
        );

    \I__1242\ : Sp12to4
    port map (
            O => \N__5663\,
            I => \N__5655\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5660\,
            I => \N__5655\
        );

    \I__1240\ : Span12Mux_h
    port map (
            O => \N__5655\,
            I => \N__5652\
        );

    \I__1239\ : Odrv12
    port map (
            O => \N__5652\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__1238\ : IoInMux
    port map (
            O => \N__5649\,
            I => \N__5646\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__5646\,
            I => \N__5643\
        );

    \I__1236\ : Span4Mux_s3_v
    port map (
            O => \N__5643\,
            I => \N__5640\
        );

    \I__1235\ : Span4Mux_h
    port map (
            O => \N__5640\,
            I => \N__5637\
        );

    \I__1234\ : Sp12to4
    port map (
            O => \N__5637\,
            I => \N__5634\
        );

    \I__1233\ : Span12Mux_s11_v
    port map (
            O => \N__5634\,
            I => \N__5631\
        );

    \I__1232\ : Span12Mux_h
    port map (
            O => \N__5631\,
            I => \N__5628\
        );

    \I__1231\ : Odrv12
    port map (
            O => \N__5628\,
            I => \N_124\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__5625\,
            I => \N__5622\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5619\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5619\,
            I => \N__5615\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5612\
        );

    \I__1226\ : Span4Mux_v
    port map (
            O => \N__5615\,
            I => \N__5606\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__5612\,
            I => \N__5606\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5603\
        );

    \I__1223\ : Span4Mux_v
    port map (
            O => \N__5606\,
            I => \N__5600\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__5603\,
            I => \N__5597\
        );

    \I__1221\ : Span4Mux_v
    port map (
            O => \N__5600\,
            I => \N__5592\
        );

    \I__1220\ : Span4Mux_v
    port map (
            O => \N__5597\,
            I => \N__5592\
        );

    \I__1219\ : Span4Mux_v
    port map (
            O => \N__5592\,
            I => \N__5589\
        );

    \I__1218\ : Span4Mux_h
    port map (
            O => \N__5589\,
            I => \N__5586\
        );

    \I__1217\ : Sp12to4
    port map (
            O => \N__5586\,
            I => \N__5583\
        );

    \I__1216\ : Odrv12
    port map (
            O => \N__5583\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5577\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__5577\,
            I => \N__5573\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5570\
        );

    \I__1212\ : Odrv12
    port map (
            O => \N__5573\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5570\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__1210\ : IoInMux
    port map (
            O => \N__5565\,
            I => \N__5562\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__5562\,
            I => \N__5559\
        );

    \I__1208\ : Span4Mux_s1_v
    port map (
            O => \N__5559\,
            I => \N__5556\
        );

    \I__1207\ : Span4Mux_h
    port map (
            O => \N__5556\,
            I => \N__5553\
        );

    \I__1206\ : Span4Mux_v
    port map (
            O => \N__5553\,
            I => \N__5550\
        );

    \I__1205\ : Span4Mux_v
    port map (
            O => \N__5550\,
            I => \N__5547\
        );

    \I__1204\ : Sp12to4
    port map (
            O => \N__5547\,
            I => \N__5544\
        );

    \I__1203\ : Odrv12
    port map (
            O => \N__5544\,
            I => \N_126\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5537\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5534\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5537\,
            I => \N__5531\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5534\,
            I => \N__5528\
        );

    \I__1198\ : Span4Mux_v
    port map (
            O => \N__5531\,
            I => \N__5522\
        );

    \I__1197\ : Span4Mux_v
    port map (
            O => \N__5528\,
            I => \N__5522\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5519\
        );

    \I__1195\ : Sp12to4
    port map (
            O => \N__5522\,
            I => \N__5514\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5519\,
            I => \N__5514\
        );

    \I__1193\ : Span12Mux_h
    port map (
            O => \N__5514\,
            I => \N__5511\
        );

    \I__1192\ : Odrv12
    port map (
            O => \N__5511\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5508\,
            I => \N__5504\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__5507\,
            I => \N__5501\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5504\,
            I => \N__5498\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5501\,
            I => \N__5495\
        );

    \I__1187\ : Odrv12
    port map (
            O => \N__5498\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5495\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__1185\ : IoInMux
    port map (
            O => \N__5490\,
            I => \N__5487\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__5487\,
            I => \N__5484\
        );

    \I__1183\ : IoSpan4Mux
    port map (
            O => \N__5484\,
            I => \N__5481\
        );

    \I__1182\ : IoSpan4Mux
    port map (
            O => \N__5481\,
            I => \N__5478\
        );

    \I__1181\ : Span4Mux_s1_v
    port map (
            O => \N__5478\,
            I => \N__5475\
        );

    \I__1180\ : Sp12to4
    port map (
            O => \N__5475\,
            I => \N__5472\
        );

    \I__1179\ : Span12Mux_s9_v
    port map (
            O => \N__5472\,
            I => \N__5469\
        );

    \I__1178\ : Odrv12
    port map (
            O => \N__5469\,
            I => \N_123\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5463\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__5463\,
            I => \N__5459\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5462\,
            I => \N__5456\
        );

    \I__1174\ : Odrv12
    port map (
            O => \N__5459\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5456\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__5451\,
            I => \N__5448\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5445\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5445\,
            I => \N__5441\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5437\
        );

    \I__1168\ : Span4Mux_v
    port map (
            O => \N__5441\,
            I => \N__5434\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5440\,
            I => \N__5431\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5437\,
            I => \N__5428\
        );

    \I__1165\ : Span4Mux_h
    port map (
            O => \N__5434\,
            I => \N__5423\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5431\,
            I => \N__5423\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__5428\,
            I => \N__5420\
        );

    \I__1162\ : Span4Mux_v
    port map (
            O => \N__5423\,
            I => \N__5417\
        );

    \I__1161\ : Sp12to4
    port map (
            O => \N__5420\,
            I => \N__5412\
        );

    \I__1160\ : Sp12to4
    port map (
            O => \N__5417\,
            I => \N__5412\
        );

    \I__1159\ : Span12Mux_h
    port map (
            O => \N__5412\,
            I => \N__5409\
        );

    \I__1158\ : Odrv12
    port map (
            O => \N__5409\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1157\ : IoInMux
    port map (
            O => \N__5406\,
            I => \N__5403\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5403\,
            I => \N__5400\
        );

    \I__1155\ : Span4Mux_s0_v
    port map (
            O => \N__5400\,
            I => \N__5397\
        );

    \I__1154\ : Sp12to4
    port map (
            O => \N__5397\,
            I => \N__5394\
        );

    \I__1153\ : Span12Mux_h
    port map (
            O => \N__5394\,
            I => \N__5391\
        );

    \I__1152\ : Odrv12
    port map (
            O => \N__5391\,
            I => \N_127\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5388\,
            I => \N__5385\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5385\,
            I => \N__5377\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5370\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5383\,
            I => \N__5370\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5382\,
            I => \N__5370\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5381\,
            I => \N__5367\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5364\
        );

    \I__1144\ : Span4Mux_v
    port map (
            O => \N__5377\,
            I => \N__5361\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5370\,
            I => \N__5358\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__5367\,
            I => \N__5355\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5364\,
            I => \N__5352\
        );

    \I__1140\ : Sp12to4
    port map (
            O => \N__5361\,
            I => \N__5347\
        );

    \I__1139\ : Span4Mux_h
    port map (
            O => \N__5358\,
            I => \N__5344\
        );

    \I__1138\ : Span4Mux_v
    port map (
            O => \N__5355\,
            I => \N__5339\
        );

    \I__1137\ : Span4Mux_v
    port map (
            O => \N__5352\,
            I => \N__5339\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5351\,
            I => \N__5334\
        );

    \I__1135\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5334\
        );

    \I__1134\ : Span12Mux_h
    port map (
            O => \N__5347\,
            I => \N__5331\
        );

    \I__1133\ : Span4Mux_v
    port map (
            O => \N__5344\,
            I => \N__5328\
        );

    \I__1132\ : Sp12to4
    port map (
            O => \N__5339\,
            I => \N__5323\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__5334\,
            I => \N__5323\
        );

    \I__1130\ : Span12Mux_v
    port map (
            O => \N__5331\,
            I => \N__5316\
        );

    \I__1129\ : Sp12to4
    port map (
            O => \N__5328\,
            I => \N__5316\
        );

    \I__1128\ : Span12Mux_h
    port map (
            O => \N__5323\,
            I => \N__5316\
        );

    \I__1127\ : Span12Mux_v
    port map (
            O => \N__5316\,
            I => \N__5313\
        );

    \I__1126\ : Odrv12
    port map (
            O => \N__5313\,
            I => \TEAn_c\
        );

    \I__1125\ : IoInMux
    port map (
            O => \N__5310\,
            I => \N__5307\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5307\,
            I => \N__5304\
        );

    \I__1123\ : Span12Mux_s8_v
    port map (
            O => \N__5304\,
            I => \N__5301\
        );

    \I__1122\ : Odrv12
    port map (
            O => \N__5301\,
            I => \U111_CYCLE_SM_TEA_CPUn_0_i\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5298\,
            I => \N__5295\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__5295\,
            I => \N__5292\
        );

    \I__1119\ : Span4Mux_v
    port map (
            O => \N__5292\,
            I => \N__5289\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__5289\,
            I => \N__5286\
        );

    \I__1117\ : Sp12to4
    port map (
            O => \N__5286\,
            I => \N__5283\
        );

    \I__1116\ : Span12Mux_h
    port map (
            O => \N__5283\,
            I => \N__5280\
        );

    \I__1115\ : Odrv12
    port map (
            O => \N__5280\,
            I => \D_UU_040_in_1\
        );

    \I__1114\ : IoInMux
    port map (
            O => \N__5277\,
            I => \N__5273\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5270\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__5273\,
            I => \N__5267\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__5270\,
            I => \N__5264\
        );

    \I__1110\ : Span4Mux_s3_h
    port map (
            O => \N__5267\,
            I => \N__5261\
        );

    \I__1109\ : Span4Mux_h
    port map (
            O => \N__5264\,
            I => \N__5258\
        );

    \I__1108\ : Sp12to4
    port map (
            O => \N__5261\,
            I => \N__5255\
        );

    \I__1107\ : Sp12to4
    port map (
            O => \N__5258\,
            I => \N__5252\
        );

    \I__1106\ : Span12Mux_v
    port map (
            O => \N__5255\,
            I => \N__5249\
        );

    \I__1105\ : Span12Mux_v
    port map (
            O => \N__5252\,
            I => \N__5246\
        );

    \I__1104\ : Span12Mux_h
    port map (
            O => \N__5249\,
            I => \N__5241\
        );

    \I__1103\ : Span12Mux_v
    port map (
            O => \N__5246\,
            I => \N__5241\
        );

    \I__1102\ : Span12Mux_h
    port map (
            O => \N__5241\,
            I => \N__5238\
        );

    \I__1101\ : Odrv12
    port map (
            O => \N__5238\,
            I => \D_LM_040_in_1\
        );

    \I__1100\ : IoInMux
    port map (
            O => \N__5235\,
            I => \N__5232\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5232\,
            I => \N__5229\
        );

    \I__1098\ : Span12Mux_s0_h
    port map (
            O => \N__5229\,
            I => \N__5226\
        );

    \I__1097\ : Span12Mux_h
    port map (
            O => \N__5226\,
            I => \N__5223\
        );

    \I__1096\ : Odrv12
    port map (
            O => \N__5223\,
            I => \un1_D_UU_040_1\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5217\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__5217\,
            I => \N__5214\
        );

    \I__1093\ : Span4Mux_v
    port map (
            O => \N__5214\,
            I => \N__5211\
        );

    \I__1092\ : Span4Mux_v
    port map (
            O => \N__5211\,
            I => \N__5208\
        );

    \I__1091\ : Sp12to4
    port map (
            O => \N__5208\,
            I => \N__5205\
        );

    \I__1090\ : Span12Mux_h
    port map (
            O => \N__5205\,
            I => \N__5202\
        );

    \I__1089\ : Odrv12
    port map (
            O => \N__5202\,
            I => \D_UM_040_in_7\
        );

    \I__1088\ : IoInMux
    port map (
            O => \N__5199\,
            I => \N__5195\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5198\,
            I => \N__5192\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5195\,
            I => \N__5189\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5192\,
            I => \N__5186\
        );

    \I__1084\ : IoSpan4Mux
    port map (
            O => \N__5189\,
            I => \N__5183\
        );

    \I__1083\ : Span4Mux_h
    port map (
            O => \N__5186\,
            I => \N__5180\
        );

    \I__1082\ : Span4Mux_s3_h
    port map (
            O => \N__5183\,
            I => \N__5177\
        );

    \I__1081\ : Sp12to4
    port map (
            O => \N__5180\,
            I => \N__5174\
        );

    \I__1080\ : Sp12to4
    port map (
            O => \N__5177\,
            I => \N__5171\
        );

    \I__1079\ : Span12Mux_v
    port map (
            O => \N__5174\,
            I => \N__5168\
        );

    \I__1078\ : Span12Mux_v
    port map (
            O => \N__5171\,
            I => \N__5165\
        );

    \I__1077\ : Span12Mux_h
    port map (
            O => \N__5168\,
            I => \N__5162\
        );

    \I__1076\ : Span12Mux_h
    port map (
            O => \N__5165\,
            I => \N__5159\
        );

    \I__1075\ : Span12Mux_v
    port map (
            O => \N__5162\,
            I => \N__5154\
        );

    \I__1074\ : Span12Mux_h
    port map (
            O => \N__5159\,
            I => \N__5154\
        );

    \I__1073\ : Odrv12
    port map (
            O => \N__5154\,
            I => \D_LL_040_in_7\
        );

    \I__1072\ : IoInMux
    port map (
            O => \N__5151\,
            I => \N__5148\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__5148\,
            I => \N__5145\
        );

    \I__1070\ : IoSpan4Mux
    port map (
            O => \N__5145\,
            I => \N__5142\
        );

    \I__1069\ : Sp12to4
    port map (
            O => \N__5142\,
            I => \N__5139\
        );

    \I__1068\ : Span12Mux_s6_h
    port map (
            O => \N__5139\,
            I => \N__5136\
        );

    \I__1067\ : Odrv12
    port map (
            O => \N__5136\,
            I => \un1_D_UM_040_7\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5130\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5130\,
            I => \N__5127\
        );

    \I__1064\ : Odrv4
    port map (
            O => \N__5127\,
            I => \U111_CYCLE_SM.LATCH_EN_5\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5124\,
            I => \N__5116\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5123\,
            I => \N__5116\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5109\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5109\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5116\,
            I => \N__5106\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5101\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5101\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__5109\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1055\ : Odrv4
    port map (
            O => \N__5106\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5101\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5090\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5093\,
            I => \N__5083\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5090\,
            I => \N__5080\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5089\,
            I => \N__5075\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5075\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5072\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5069\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__5083\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__5080\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__5075\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5072\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5069\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1041\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5055\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5055\,
            I => \N__5052\
        );

    \I__1039\ : Odrv4
    port map (
            O => \N__5052\,
            I => \U111_CYCLE_SM.N_57\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5046\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__5046\,
            I => \N__5041\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5045\,
            I => \N__5038\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5035\
        );

    \I__1034\ : Span4Mux_v
    port map (
            O => \N__5041\,
            I => \N__5028\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__5038\,
            I => \N__5028\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5035\,
            I => \N__5028\
        );

    \I__1031\ : Span4Mux_v
    port map (
            O => \N__5028\,
            I => \N__5025\
        );

    \I__1030\ : Span4Mux_v
    port map (
            O => \N__5025\,
            I => \N__5022\
        );

    \I__1029\ : Span4Mux_v
    port map (
            O => \N__5022\,
            I => \N__5019\
        );

    \I__1028\ : Sp12to4
    port map (
            O => \N__5019\,
            I => \N__5016\
        );

    \I__1027\ : Odrv12
    port map (
            O => \N__5016\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__5013\,
            I => \N__5009\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5012\,
            I => \N__5006\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5009\,
            I => \N__5003\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5006\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__5003\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__1021\ : IoInMux
    port map (
            O => \N__4998\,
            I => \N__4995\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__4995\,
            I => \N__4992\
        );

    \I__1019\ : Span4Mux_s0_h
    port map (
            O => \N__4992\,
            I => \N__4989\
        );

    \I__1018\ : Sp12to4
    port map (
            O => \N__4989\,
            I => \N__4986\
        );

    \I__1017\ : Span12Mux_v
    port map (
            O => \N__4986\,
            I => \N__4983\
        );

    \I__1016\ : Span12Mux_h
    port map (
            O => \N__4983\,
            I => \N__4980\
        );

    \I__1015\ : Odrv12
    port map (
            O => \N__4980\,
            I => \un1_D_UM_AMIGA_7\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__4977\,
            I => \N__4974\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4974\,
            I => \N__4970\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4967\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4970\,
            I => \N__4964\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4967\,
            I => \N__4961\
        );

    \I__1009\ : Span4Mux_v
    port map (
            O => \N__4964\,
            I => \N__4957\
        );

    \I__1008\ : Span4Mux_v
    port map (
            O => \N__4961\,
            I => \N__4954\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4951\
        );

    \I__1006\ : Span4Mux_h
    port map (
            O => \N__4957\,
            I => \N__4948\
        );

    \I__1005\ : Sp12to4
    port map (
            O => \N__4954\,
            I => \N__4943\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__4951\,
            I => \N__4943\
        );

    \I__1003\ : Sp12to4
    port map (
            O => \N__4948\,
            I => \N__4938\
        );

    \I__1002\ : Span12Mux_h
    port map (
            O => \N__4943\,
            I => \N__4938\
        );

    \I__1001\ : Span12Mux_v
    port map (
            O => \N__4938\,
            I => \N__4935\
        );

    \I__1000\ : Odrv12
    port map (
            O => \N__4935\,
            I => \PORTSIZE_c\
        );

    \I__999\ : IoInMux
    port map (
            O => \N__4932\,
            I => \N__4926\
        );

    \I__998\ : IoInMux
    port map (
            O => \N__4931\,
            I => \N__4923\
        );

    \I__997\ : IoInMux
    port map (
            O => \N__4930\,
            I => \N__4920\
        );

    \I__996\ : IoInMux
    port map (
            O => \N__4929\,
            I => \N__4911\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4926\,
            I => \N__4902\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4923\,
            I => \N__4902\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4920\,
            I => \N__4902\
        );

    \I__992\ : IoInMux
    port map (
            O => \N__4919\,
            I => \N__4899\
        );

    \I__991\ : IoInMux
    port map (
            O => \N__4918\,
            I => \N__4896\
        );

    \I__990\ : IoInMux
    port map (
            O => \N__4917\,
            I => \N__4893\
        );

    \I__989\ : IoInMux
    port map (
            O => \N__4916\,
            I => \N__4886\
        );

    \I__988\ : IoInMux
    port map (
            O => \N__4915\,
            I => \N__4883\
        );

    \I__987\ : IoInMux
    port map (
            O => \N__4914\,
            I => \N__4880\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__4911\,
            I => \N__4873\
        );

    \I__985\ : IoInMux
    port map (
            O => \N__4910\,
            I => \N__4870\
        );

    \I__984\ : IoInMux
    port map (
            O => \N__4909\,
            I => \N__4867\
        );

    \I__983\ : IoSpan4Mux
    port map (
            O => \N__4902\,
            I => \N__4854\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4899\,
            I => \N__4854\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__4896\,
            I => \N__4854\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4893\,
            I => \N__4854\
        );

    \I__979\ : IoInMux
    port map (
            O => \N__4892\,
            I => \N__4851\
        );

    \I__978\ : IoInMux
    port map (
            O => \N__4891\,
            I => \N__4848\
        );

    \I__977\ : IoInMux
    port map (
            O => \N__4890\,
            I => \N__4845\
        );

    \I__976\ : IoInMux
    port map (
            O => \N__4889\,
            I => \N__4842\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__4886\,
            I => \N__4835\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4883\,
            I => \N__4830\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__4880\,
            I => \N__4830\
        );

    \I__972\ : IoInMux
    port map (
            O => \N__4879\,
            I => \N__4827\
        );

    \I__971\ : IoInMux
    port map (
            O => \N__4878\,
            I => \N__4824\
        );

    \I__970\ : IoInMux
    port map (
            O => \N__4877\,
            I => \N__4821\
        );

    \I__969\ : IoInMux
    port map (
            O => \N__4876\,
            I => \N__4818\
        );

    \I__968\ : IoSpan4Mux
    port map (
            O => \N__4873\,
            I => \N__4811\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4870\,
            I => \N__4811\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4867\,
            I => \N__4811\
        );

    \I__965\ : IoInMux
    port map (
            O => \N__4866\,
            I => \N__4808\
        );

    \I__964\ : IoInMux
    port map (
            O => \N__4865\,
            I => \N__4805\
        );

    \I__963\ : IoInMux
    port map (
            O => \N__4864\,
            I => \N__4802\
        );

    \I__962\ : IoInMux
    port map (
            O => \N__4863\,
            I => \N__4799\
        );

    \I__961\ : IoSpan4Mux
    port map (
            O => \N__4854\,
            I => \N__4788\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4851\,
            I => \N__4788\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4848\,
            I => \N__4788\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4845\,
            I => \N__4788\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4842\,
            I => \N__4788\
        );

    \I__956\ : IoInMux
    port map (
            O => \N__4841\,
            I => \N__4785\
        );

    \I__955\ : IoInMux
    port map (
            O => \N__4840\,
            I => \N__4782\
        );

    \I__954\ : IoInMux
    port map (
            O => \N__4839\,
            I => \N__4779\
        );

    \I__953\ : IoInMux
    port map (
            O => \N__4838\,
            I => \N__4776\
        );

    \I__952\ : IoSpan4Mux
    port map (
            O => \N__4835\,
            I => \N__4772\
        );

    \I__951\ : IoSpan4Mux
    port map (
            O => \N__4830\,
            I => \N__4761\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__4827\,
            I => \N__4761\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4824\,
            I => \N__4761\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4821\,
            I => \N__4761\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4818\,
            I => \N__4761\
        );

    \I__946\ : IoSpan4Mux
    port map (
            O => \N__4811\,
            I => \N__4750\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4808\,
            I => \N__4750\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4805\,
            I => \N__4750\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4802\,
            I => \N__4750\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4799\,
            I => \N__4750\
        );

    \I__941\ : IoSpan4Mux
    port map (
            O => \N__4788\,
            I => \N__4739\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4785\,
            I => \N__4739\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4782\,
            I => \N__4739\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4779\,
            I => \N__4739\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4776\,
            I => \N__4739\
        );

    \I__936\ : IoInMux
    port map (
            O => \N__4775\,
            I => \N__4736\
        );

    \I__935\ : Span4Mux_s0_h
    port map (
            O => \N__4772\,
            I => \N__4731\
        );

    \I__934\ : IoSpan4Mux
    port map (
            O => \N__4761\,
            I => \N__4728\
        );

    \I__933\ : IoSpan4Mux
    port map (
            O => \N__4750\,
            I => \N__4721\
        );

    \I__932\ : IoSpan4Mux
    port map (
            O => \N__4739\,
            I => \N__4721\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4736\,
            I => \N__4721\
        );

    \I__930\ : IoInMux
    port map (
            O => \N__4735\,
            I => \N__4718\
        );

    \I__929\ : IoInMux
    port map (
            O => \N__4734\,
            I => \N__4715\
        );

    \I__928\ : Span4Mux_h
    port map (
            O => \N__4731\,
            I => \N__4712\
        );

    \I__927\ : Span4Mux_s3_v
    port map (
            O => \N__4728\,
            I => \N__4709\
        );

    \I__926\ : IoSpan4Mux
    port map (
            O => \N__4721\,
            I => \N__4705\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4718\,
            I => \N__4700\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4715\,
            I => \N__4700\
        );

    \I__923\ : Span4Mux_h
    port map (
            O => \N__4712\,
            I => \N__4695\
        );

    \I__922\ : Span4Mux_v
    port map (
            O => \N__4709\,
            I => \N__4695\
        );

    \I__921\ : IoInMux
    port map (
            O => \N__4708\,
            I => \N__4692\
        );

    \I__920\ : Sp12to4
    port map (
            O => \N__4705\,
            I => \N__4689\
        );

    \I__919\ : Span12Mux_s8_h
    port map (
            O => \N__4700\,
            I => \N__4686\
        );

    \I__918\ : Sp12to4
    port map (
            O => \N__4695\,
            I => \N__4683\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4692\,
            I => \N__4680\
        );

    \I__916\ : Span12Mux_h
    port map (
            O => \N__4689\,
            I => \N__4677\
        );

    \I__915\ : Span12Mux_v
    port map (
            O => \N__4686\,
            I => \N__4670\
        );

    \I__914\ : Span12Mux_v
    port map (
            O => \N__4683\,
            I => \N__4670\
        );

    \I__913\ : Span12Mux_s8_h
    port map (
            O => \N__4680\,
            I => \N__4670\
        );

    \I__912\ : Odrv12
    port map (
            O => \N__4677\,
            I => \U111_CYCLE_SM_OFFBOARD_EN_0\
        );

    \I__911\ : Odrv12
    port map (
            O => \N__4670\,
            I => \U111_CYCLE_SM_OFFBOARD_EN_0\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__4665\,
            I => \U111_CYCLE_SM.un4_TS_OUT_i_0_cascade_\
        );

    \I__909\ : InMux
    port map (
            O => \N__4662\,
            I => \N__4659\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4659\,
            I => \U111_CYCLE_SM.N_106\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__4656\,
            I => \N__4653\
        );

    \I__906\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4650\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4650\,
            I => \N__4647\
        );

    \I__904\ : Span4Mux_v
    port map (
            O => \N__4647\,
            I => \N__4637\
        );

    \I__903\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4634\
        );

    \I__902\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4631\
        );

    \I__901\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4624\
        );

    \I__900\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4624\
        );

    \I__899\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4624\
        );

    \I__898\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4619\
        );

    \I__897\ : InMux
    port map (
            O => \N__4640\,
            I => \N__4619\
        );

    \I__896\ : Sp12to4
    port map (
            O => \N__4637\,
            I => \N__4612\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4634\,
            I => \N__4612\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4631\,
            I => \N__4612\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4624\,
            I => \N__4607\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4619\,
            I => \N__4607\
        );

    \I__891\ : Span12Mux_h
    port map (
            O => \N__4612\,
            I => \N__4604\
        );

    \I__890\ : Span12Mux_v
    port map (
            O => \N__4607\,
            I => \N__4601\
        );

    \I__889\ : Span12Mux_v
    port map (
            O => \N__4604\,
            I => \N__4598\
        );

    \I__888\ : Odrv12
    port map (
            O => \N__4601\,
            I => \RESETn_c\
        );

    \I__887\ : Odrv12
    port map (
            O => \N__4598\,
            I => \RESETn_c\
        );

    \I__886\ : InMux
    port map (
            O => \N__4593\,
            I => \N__4590\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4590\,
            I => \U111_CYCLE_SM.N_140\
        );

    \I__884\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4582\
        );

    \I__883\ : InMux
    port map (
            O => \N__4586\,
            I => \N__4579\
        );

    \I__882\ : InMux
    port map (
            O => \N__4585\,
            I => \N__4576\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__4582\,
            I => \U111_CYCLE_SM.N_107\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4579\,
            I => \U111_CYCLE_SM.N_107\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4576\,
            I => \U111_CYCLE_SM.N_107\
        );

    \I__878\ : InMux
    port map (
            O => \N__4569\,
            I => \N__4560\
        );

    \I__877\ : InMux
    port map (
            O => \N__4568\,
            I => \N__4560\
        );

    \I__876\ : InMux
    port map (
            O => \N__4567\,
            I => \N__4553\
        );

    \I__875\ : InMux
    port map (
            O => \N__4566\,
            I => \N__4553\
        );

    \I__874\ : InMux
    port map (
            O => \N__4565\,
            I => \N__4553\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4560\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4553\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\
        );

    \I__871\ : IoInMux
    port map (
            O => \N__4548\,
            I => \N__4544\
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__4547\,
            I => \N__4539\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4544\,
            I => \N__4534\
        );

    \I__868\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4531\
        );

    \I__867\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4524\
        );

    \I__866\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4524\
        );

    \I__865\ : InMux
    port map (
            O => \N__4538\,
            I => \N__4524\
        );

    \I__864\ : CascadeMux
    port map (
            O => \N__4537\,
            I => \N__4521\
        );

    \I__863\ : Span4Mux_s1_v
    port map (
            O => \N__4534\,
            I => \N__4516\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4531\,
            I => \N__4511\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4524\,
            I => \N__4511\
        );

    \I__860\ : InMux
    port map (
            O => \N__4521\,
            I => \N__4506\
        );

    \I__859\ : InMux
    port map (
            O => \N__4520\,
            I => \N__4506\
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__4519\,
            I => \N__4503\
        );

    \I__857\ : Span4Mux_v
    port map (
            O => \N__4516\,
            I => \N__4500\
        );

    \I__856\ : Span4Mux_v
    port map (
            O => \N__4511\,
            I => \N__4497\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4506\,
            I => \N__4494\
        );

    \I__854\ : InMux
    port map (
            O => \N__4503\,
            I => \N__4491\
        );

    \I__853\ : Sp12to4
    port map (
            O => \N__4500\,
            I => \N__4487\
        );

    \I__852\ : Span4Mux_h
    port map (
            O => \N__4497\,
            I => \N__4484\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__4494\,
            I => \N__4481\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4491\,
            I => \N__4478\
        );

    \I__849\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4475\
        );

    \I__848\ : Span12Mux_h
    port map (
            O => \N__4487\,
            I => \N__4472\
        );

    \I__847\ : Sp12to4
    port map (
            O => \N__4484\,
            I => \N__4469\
        );

    \I__846\ : Span4Mux_v
    port map (
            O => \N__4481\,
            I => \N__4466\
        );

    \I__845\ : Span4Mux_h
    port map (
            O => \N__4478\,
            I => \N__4463\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4475\,
            I => \N__4460\
        );

    \I__843\ : Span12Mux_v
    port map (
            O => \N__4472\,
            I => \N__4449\
        );

    \I__842\ : Span12Mux_h
    port map (
            O => \N__4469\,
            I => \N__4449\
        );

    \I__841\ : Sp12to4
    port map (
            O => \N__4466\,
            I => \N__4449\
        );

    \I__840\ : Sp12to4
    port map (
            O => \N__4463\,
            I => \N__4449\
        );

    \I__839\ : Span12Mux_h
    port map (
            O => \N__4460\,
            I => \N__4449\
        );

    \I__838\ : Span12Mux_v
    port map (
            O => \N__4449\,
            I => \N__4446\
        );

    \I__837\ : Odrv12
    port map (
            O => \N__4446\,
            I => \TACKn_in\
        );

    \I__836\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4440\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4440\,
            I => \N__4437\
        );

    \I__834\ : Span12Mux_v
    port map (
            O => \N__4437\,
            I => \N__4434\
        );

    \I__833\ : Odrv12
    port map (
            O => \N__4434\,
            I => \D_LM_AMIGA_in_4\
        );

    \I__832\ : IoInMux
    port map (
            O => \N__4431\,
            I => \N__4428\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4428\,
            I => \N__4425\
        );

    \I__830\ : IoSpan4Mux
    port map (
            O => \N__4425\,
            I => \N__4422\
        );

    \I__829\ : Span4Mux_s3_h
    port map (
            O => \N__4422\,
            I => \N__4419\
        );

    \I__828\ : Span4Mux_v
    port map (
            O => \N__4419\,
            I => \N__4416\
        );

    \I__827\ : Span4Mux_h
    port map (
            O => \N__4416\,
            I => \N__4413\
        );

    \I__826\ : Sp12to4
    port map (
            O => \N__4413\,
            I => \N__4410\
        );

    \I__825\ : Odrv12
    port map (
            O => \N__4410\,
            I => \N_118\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__4407\,
            I => \N__4404\
        );

    \I__823\ : InMux
    port map (
            O => \N__4404\,
            I => \N__4401\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4401\,
            I => \N__4396\
        );

    \I__821\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4393\
        );

    \I__820\ : InMux
    port map (
            O => \N__4399\,
            I => \N__4390\
        );

    \I__819\ : Span4Mux_h
    port map (
            O => \N__4396\,
            I => \N__4385\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__4393\,
            I => \N__4385\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4390\,
            I => \N__4382\
        );

    \I__816\ : Span4Mux_v
    port map (
            O => \N__4385\,
            I => \N__4379\
        );

    \I__815\ : Sp12to4
    port map (
            O => \N__4382\,
            I => \N__4376\
        );

    \I__814\ : Sp12to4
    port map (
            O => \N__4379\,
            I => \N__4373\
        );

    \I__813\ : Span12Mux_v
    port map (
            O => \N__4376\,
            I => \N__4370\
        );

    \I__812\ : Span12Mux_h
    port map (
            O => \N__4373\,
            I => \N__4367\
        );

    \I__811\ : Odrv12
    port map (
            O => \N__4370\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__810\ : Odrv12
    port map (
            O => \N__4367\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__809\ : InMux
    port map (
            O => \N__4362\,
            I => \N__4359\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4359\,
            I => \N__4355\
        );

    \I__807\ : InMux
    port map (
            O => \N__4358\,
            I => \N__4352\
        );

    \I__806\ : Odrv12
    port map (
            O => \N__4355\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4352\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__804\ : IoInMux
    port map (
            O => \N__4347\,
            I => \N__4344\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4344\,
            I => \N__4341\
        );

    \I__802\ : IoSpan4Mux
    port map (
            O => \N__4341\,
            I => \N__4338\
        );

    \I__801\ : IoSpan4Mux
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__800\ : Sp12to4
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__799\ : Span12Mux_s9_h
    port map (
            O => \N__4332\,
            I => \N__4329\
        );

    \I__798\ : Odrv12
    port map (
            O => \N__4329\,
            I => \un1_D_UM_AMIGA_1\
        );

    \I__797\ : InMux
    port map (
            O => \N__4326\,
            I => \N__4323\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4323\,
            I => \N__4320\
        );

    \I__795\ : Span4Mux_h
    port map (
            O => \N__4320\,
            I => \N__4317\
        );

    \I__794\ : Span4Mux_v
    port map (
            O => \N__4317\,
            I => \N__4314\
        );

    \I__793\ : Sp12to4
    port map (
            O => \N__4314\,
            I => \N__4311\
        );

    \I__792\ : Odrv12
    port map (
            O => \N__4311\,
            I => \D_LM_AMIGA_in_6\
        );

    \I__791\ : IoInMux
    port map (
            O => \N__4308\,
            I => \N__4305\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4305\,
            I => \N__4302\
        );

    \I__789\ : Span12Mux_s10_h
    port map (
            O => \N__4302\,
            I => \N__4299\
        );

    \I__788\ : Odrv12
    port map (
            O => \N__4299\,
            I => \N_116\
        );

    \I__787\ : IoInMux
    port map (
            O => \N__4296\,
            I => \N__4293\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4293\,
            I => \N__4290\
        );

    \I__785\ : Span12Mux_s6_v
    port map (
            O => \N__4290\,
            I => \N__4287\
        );

    \I__784\ : Odrv12
    port map (
            O => \N__4287\,
            I => \N_102_i\
        );

    \I__783\ : IoInMux
    port map (
            O => \N__4284\,
            I => \N__4281\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__4281\,
            I => \N__4278\
        );

    \I__781\ : IoSpan4Mux
    port map (
            O => \N__4278\,
            I => \N__4275\
        );

    \I__780\ : Span4Mux_s3_v
    port map (
            O => \N__4275\,
            I => \N__4272\
        );

    \I__779\ : Span4Mux_h
    port map (
            O => \N__4272\,
            I => \N__4269\
        );

    \I__778\ : Odrv4
    port map (
            O => \N__4269\,
            I => \BUFDIR_c\
        );

    \I__777\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4257\
        );

    \I__776\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4257\
        );

    \I__775\ : InMux
    port map (
            O => \N__4264\,
            I => \N__4257\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4257\,
            I => \N__4254\
        );

    \I__773\ : Span4Mux_h
    port map (
            O => \N__4254\,
            I => \N__4251\
        );

    \I__772\ : Span4Mux_v
    port map (
            O => \N__4251\,
            I => \N__4248\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__4248\,
            I => \BBn_c\
        );

    \I__770\ : IoInMux
    port map (
            O => \N__4245\,
            I => \N__4242\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4242\,
            I => \N__4239\
        );

    \I__768\ : Span4Mux_s3_v
    port map (
            O => \N__4239\,
            I => \N__4236\
        );

    \I__767\ : Span4Mux_h
    port map (
            O => \N__4236\,
            I => \N__4233\
        );

    \I__766\ : Odrv4
    port map (
            O => \N__4233\,
            I => \N_104\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__4230\,
            I => \N__4226\
        );

    \I__764\ : InMux
    port map (
            O => \N__4229\,
            I => \N__4223\
        );

    \I__763\ : InMux
    port map (
            O => \N__4226\,
            I => \N__4220\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4223\,
            I => \N__4217\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4220\,
            I => \N__4214\
        );

    \I__760\ : Span4Mux_v
    port map (
            O => \N__4217\,
            I => \N__4210\
        );

    \I__759\ : Span4Mux_v
    port map (
            O => \N__4214\,
            I => \N__4207\
        );

    \I__758\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4204\
        );

    \I__757\ : Span4Mux_v
    port map (
            O => \N__4210\,
            I => \N__4201\
        );

    \I__756\ : Span4Mux_v
    port map (
            O => \N__4207\,
            I => \N__4196\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4204\,
            I => \N__4196\
        );

    \I__754\ : Span4Mux_v
    port map (
            O => \N__4201\,
            I => \N__4193\
        );

    \I__753\ : Span4Mux_v
    port map (
            O => \N__4196\,
            I => \N__4190\
        );

    \I__752\ : Sp12to4
    port map (
            O => \N__4193\,
            I => \N__4185\
        );

    \I__751\ : Sp12to4
    port map (
            O => \N__4190\,
            I => \N__4185\
        );

    \I__750\ : Span12Mux_h
    port map (
            O => \N__4185\,
            I => \N__4182\
        );

    \I__749\ : Odrv12
    port map (
            O => \N__4182\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__748\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4176\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4176\,
            I => \N__4173\
        );

    \I__746\ : Span4Mux_v
    port map (
            O => \N__4173\,
            I => \N__4170\
        );

    \I__745\ : Span4Mux_v
    port map (
            O => \N__4170\,
            I => \N__4166\
        );

    \I__744\ : InMux
    port map (
            O => \N__4169\,
            I => \N__4163\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__4166\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4163\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__741\ : IoInMux
    port map (
            O => \N__4158\,
            I => \N__4155\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4155\,
            I => \N__4152\
        );

    \I__739\ : Span4Mux_s2_v
    port map (
            O => \N__4152\,
            I => \N__4149\
        );

    \I__738\ : Span4Mux_v
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__737\ : Sp12to4
    port map (
            O => \N__4146\,
            I => \N__4143\
        );

    \I__736\ : Span12Mux_s10_h
    port map (
            O => \N__4143\,
            I => \N__4140\
        );

    \I__735\ : Odrv12
    port map (
            O => \N__4140\,
            I => \N_128\
        );

    \I__734\ : InMux
    port map (
            O => \N__4137\,
            I => \N__4134\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4134\,
            I => \U111_CYCLE_SM.N_195\
        );

    \I__732\ : InMux
    port map (
            O => \N__4131\,
            I => \N__4128\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4128\,
            I => \U111_CYCLE_SM.N_132\
        );

    \I__730\ : CascadeMux
    port map (
            O => \N__4125\,
            I => \N__4121\
        );

    \I__729\ : InMux
    port map (
            O => \N__4124\,
            I => \N__4118\
        );

    \I__728\ : InMux
    port map (
            O => \N__4121\,
            I => \N__4115\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__4118\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4115\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\
        );

    \I__725\ : InMux
    port map (
            O => \N__4110\,
            I => \N__4106\
        );

    \I__724\ : InMux
    port map (
            O => \N__4109\,
            I => \N__4103\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4106\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4103\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__721\ : IoInMux
    port map (
            O => \N__4098\,
            I => \N__4095\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4095\,
            I => \N__4092\
        );

    \I__719\ : Span4Mux_s3_v
    port map (
            O => \N__4092\,
            I => \N__4089\
        );

    \I__718\ : Sp12to4
    port map (
            O => \N__4089\,
            I => \N__4086\
        );

    \I__717\ : Span12Mux_h
    port map (
            O => \N__4086\,
            I => \N__4083\
        );

    \I__716\ : Odrv12
    port map (
            O => \N__4083\,
            I => \TS_OUT\
        );

    \I__715\ : InMux
    port map (
            O => \N__4080\,
            I => \N__4077\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__4077\,
            I => \N__4074\
        );

    \I__713\ : Span4Mux_v
    port map (
            O => \N__4074\,
            I => \N__4071\
        );

    \I__712\ : Sp12to4
    port map (
            O => \N__4071\,
            I => \N__4067\
        );

    \I__711\ : IoInMux
    port map (
            O => \N__4070\,
            I => \N__4064\
        );

    \I__710\ : Span12Mux_h
    port map (
            O => \N__4067\,
            I => \N__4061\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__4064\,
            I => \N__4058\
        );

    \I__708\ : Span12Mux_v
    port map (
            O => \N__4061\,
            I => \N__4055\
        );

    \I__707\ : IoSpan4Mux
    port map (
            O => \N__4058\,
            I => \N__4052\
        );

    \I__706\ : Odrv12
    port map (
            O => \N__4055\,
            I => \TBIn_c\
        );

    \I__705\ : Odrv4
    port map (
            O => \N__4052\,
            I => \TBIn_c\
        );

    \I__704\ : InMux
    port map (
            O => \N__4047\,
            I => \N__4039\
        );

    \I__703\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4039\
        );

    \I__702\ : InMux
    port map (
            O => \N__4045\,
            I => \N__4034\
        );

    \I__701\ : InMux
    port map (
            O => \N__4044\,
            I => \N__4034\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4039\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__4034\,
            I => \U111_CYCLE_SM.BURSTZ0\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__4029\,
            I => \N__4024\
        );

    \I__697\ : InMux
    port map (
            O => \N__4028\,
            I => \N__4019\
        );

    \I__696\ : InMux
    port map (
            O => \N__4027\,
            I => \N__4019\
        );

    \I__695\ : InMux
    port map (
            O => \N__4024\,
            I => \N__4016\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4019\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__4016\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\
        );

    \I__692\ : InMux
    port map (
            O => \N__4011\,
            I => \N__4007\
        );

    \I__691\ : InMux
    port map (
            O => \N__4010\,
            I => \N__4004\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4007\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4004\,
            I => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\
        );

    \I__688\ : InMux
    port map (
            O => \N__3999\,
            I => \N__3996\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3996\,
            I => \U111_CYCLE_SM.N_109\
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__3993\,
            I => \U111_CYCLE_SM.N_109_cascade_\
        );

    \I__685\ : InMux
    port map (
            O => \N__3990\,
            I => \N__3984\
        );

    \I__684\ : InMux
    port map (
            O => \N__3989\,
            I => \N__3979\
        );

    \I__683\ : InMux
    port map (
            O => \N__3988\,
            I => \N__3979\
        );

    \I__682\ : InMux
    port map (
            O => \N__3987\,
            I => \N__3976\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3984\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3979\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3976\,
            I => \U111_CYCLE_SM.PORT_MISMATCHZ0\
        );

    \I__678\ : InMux
    port map (
            O => \N__3969\,
            I => \N__3966\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3966\,
            I => \N__3963\
        );

    \I__676\ : Span12Mux_v
    port map (
            O => \N__3963\,
            I => \N__3960\
        );

    \I__675\ : Odrv12
    port map (
            O => \N__3960\,
            I => \D_LM_AMIGA_in_5\
        );

    \I__674\ : IoInMux
    port map (
            O => \N__3957\,
            I => \N__3954\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__3954\,
            I => \N__3951\
        );

    \I__672\ : Span4Mux_s3_h
    port map (
            O => \N__3951\,
            I => \N__3948\
        );

    \I__671\ : Span4Mux_v
    port map (
            O => \N__3948\,
            I => \N__3945\
        );

    \I__670\ : Sp12to4
    port map (
            O => \N__3945\,
            I => \N__3942\
        );

    \I__669\ : Span12Mux_h
    port map (
            O => \N__3942\,
            I => \N__3939\
        );

    \I__668\ : Odrv12
    port map (
            O => \N__3939\,
            I => \N_117\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__3936\,
            I => \U111_CYCLE_SM.N_144_cascade_\
        );

    \I__666\ : InMux
    port map (
            O => \N__3933\,
            I => \N__3930\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3930\,
            I => \U111_CYCLE_SM.N_142\
        );

    \I__664\ : InMux
    port map (
            O => \N__3927\,
            I => \N__3923\
        );

    \I__663\ : InMux
    port map (
            O => \N__3926\,
            I => \N__3920\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3923\,
            I => \U111_CYCLE_SM.N_197\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3920\,
            I => \U111_CYCLE_SM.N_197\
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__3915\,
            I => \N__3908\
        );

    \I__659\ : InMux
    port map (
            O => \N__3914\,
            I => \N__3903\
        );

    \I__658\ : InMux
    port map (
            O => \N__3913\,
            I => \N__3903\
        );

    \I__657\ : InMux
    port map (
            O => \N__3912\,
            I => \N__3896\
        );

    \I__656\ : InMux
    port map (
            O => \N__3911\,
            I => \N__3896\
        );

    \I__655\ : InMux
    port map (
            O => \N__3908\,
            I => \N__3896\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3903\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3896\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__3891\,
            I => \U111_CYCLE_SM.N_195_cascade_\
        );

    \I__651\ : InMux
    port map (
            O => \N__3888\,
            I => \N__3885\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3885\,
            I => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_1_0\
        );

    \I__649\ : InMux
    port map (
            O => \N__3882\,
            I => \N__3879\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__3879\,
            I => \N__3875\
        );

    \I__647\ : IoInMux
    port map (
            O => \N__3878\,
            I => \N__3872\
        );

    \I__646\ : Span4Mux_v
    port map (
            O => \N__3875\,
            I => \N__3869\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3872\,
            I => \N__3866\
        );

    \I__644\ : Span4Mux_h
    port map (
            O => \N__3869\,
            I => \N__3863\
        );

    \I__643\ : Span4Mux_s3_h
    port map (
            O => \N__3866\,
            I => \N__3860\
        );

    \I__642\ : Span4Mux_v
    port map (
            O => \N__3863\,
            I => \N__3857\
        );

    \I__641\ : Sp12to4
    port map (
            O => \N__3860\,
            I => \N__3854\
        );

    \I__640\ : Sp12to4
    port map (
            O => \N__3857\,
            I => \N__3851\
        );

    \I__639\ : Span12Mux_v
    port map (
            O => \N__3854\,
            I => \N__3848\
        );

    \I__638\ : Span12Mux_v
    port map (
            O => \N__3851\,
            I => \N__3843\
        );

    \I__637\ : Span12Mux_h
    port map (
            O => \N__3848\,
            I => \N__3843\
        );

    \I__636\ : Span12Mux_h
    port map (
            O => \N__3843\,
            I => \N__3840\
        );

    \I__635\ : Odrv12
    port map (
            O => \N__3840\,
            I => \D_LL_040_in_3\
        );

    \I__634\ : InMux
    port map (
            O => \N__3837\,
            I => \N__3834\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3834\,
            I => \N__3831\
        );

    \I__632\ : Span4Mux_v
    port map (
            O => \N__3831\,
            I => \N__3828\
        );

    \I__631\ : Sp12to4
    port map (
            O => \N__3828\,
            I => \N__3825\
        );

    \I__630\ : Span12Mux_h
    port map (
            O => \N__3825\,
            I => \N__3822\
        );

    \I__629\ : Span12Mux_v
    port map (
            O => \N__3822\,
            I => \N__3819\
        );

    \I__628\ : Odrv12
    port map (
            O => \N__3819\,
            I => \D_UM_040_in_3\
        );

    \I__627\ : IoInMux
    port map (
            O => \N__3816\,
            I => \N__3813\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3813\,
            I => \N__3810\
        );

    \I__625\ : IoSpan4Mux
    port map (
            O => \N__3810\,
            I => \N__3807\
        );

    \I__624\ : Span4Mux_s2_h
    port map (
            O => \N__3807\,
            I => \N__3804\
        );

    \I__623\ : Span4Mux_h
    port map (
            O => \N__3804\,
            I => \N__3801\
        );

    \I__622\ : Span4Mux_h
    port map (
            O => \N__3801\,
            I => \N__3798\
        );

    \I__621\ : Odrv4
    port map (
            O => \N__3798\,
            I => \un1_D_UM_040_3\
        );

    \I__620\ : InMux
    port map (
            O => \N__3795\,
            I => \N__3792\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3792\,
            I => \N__3789\
        );

    \I__618\ : Sp12to4
    port map (
            O => \N__3789\,
            I => \N__3786\
        );

    \I__617\ : Span12Mux_v
    port map (
            O => \N__3786\,
            I => \N__3783\
        );

    \I__616\ : Odrv12
    port map (
            O => \N__3783\,
            I => \D_LM_AMIGA_in_7\
        );

    \I__615\ : IoInMux
    port map (
            O => \N__3780\,
            I => \N__3777\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3777\,
            I => \N__3774\
        );

    \I__613\ : IoSpan4Mux
    port map (
            O => \N__3774\,
            I => \N__3771\
        );

    \I__612\ : Span4Mux_s2_h
    port map (
            O => \N__3771\,
            I => \N__3768\
        );

    \I__611\ : Sp12to4
    port map (
            O => \N__3768\,
            I => \N__3765\
        );

    \I__610\ : Span12Mux_s9_h
    port map (
            O => \N__3765\,
            I => \N__3762\
        );

    \I__609\ : Odrv12
    port map (
            O => \N__3762\,
            I => \N_115\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__3759\,
            I => \N__3756\
        );

    \I__607\ : InMux
    port map (
            O => \N__3756\,
            I => \N__3753\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3753\,
            I => \N__3748\
        );

    \I__605\ : InMux
    port map (
            O => \N__3752\,
            I => \N__3745\
        );

    \I__604\ : InMux
    port map (
            O => \N__3751\,
            I => \N__3742\
        );

    \I__603\ : Span4Mux_h
    port map (
            O => \N__3748\,
            I => \N__3737\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3745\,
            I => \N__3737\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3742\,
            I => \N__3734\
        );

    \I__600\ : Span4Mux_v
    port map (
            O => \N__3737\,
            I => \N__3731\
        );

    \I__599\ : Span4Mux_v
    port map (
            O => \N__3734\,
            I => \N__3728\
        );

    \I__598\ : Span4Mux_h
    port map (
            O => \N__3731\,
            I => \N__3725\
        );

    \I__597\ : IoSpan4Mux
    port map (
            O => \N__3728\,
            I => \N__3722\
        );

    \I__596\ : Sp12to4
    port map (
            O => \N__3725\,
            I => \N__3719\
        );

    \I__595\ : IoSpan4Mux
    port map (
            O => \N__3722\,
            I => \N__3716\
        );

    \I__594\ : Odrv12
    port map (
            O => \N__3719\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__593\ : Odrv4
    port map (
            O => \N__3716\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__592\ : InMux
    port map (
            O => \N__3711\,
            I => \N__3708\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3708\,
            I => \N__3704\
        );

    \I__590\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3701\
        );

    \I__589\ : Odrv12
    port map (
            O => \N__3704\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3701\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__587\ : IoInMux
    port map (
            O => \N__3696\,
            I => \N__3693\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3693\,
            I => \N__3690\
        );

    \I__585\ : Span4Mux_s3_v
    port map (
            O => \N__3690\,
            I => \N__3687\
        );

    \I__584\ : Span4Mux_h
    port map (
            O => \N__3687\,
            I => \N__3684\
        );

    \I__583\ : Span4Mux_h
    port map (
            O => \N__3684\,
            I => \N__3681\
        );

    \I__582\ : Span4Mux_h
    port map (
            O => \N__3681\,
            I => \N__3678\
        );

    \I__581\ : Span4Mux_h
    port map (
            O => \N__3678\,
            I => \N__3675\
        );

    \I__580\ : Odrv4
    port map (
            O => \N__3675\,
            I => \N_129\
        );

    \I__579\ : InMux
    port map (
            O => \N__3672\,
            I => \N__3669\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3669\,
            I => \N__3666\
        );

    \I__577\ : Span4Mux_v
    port map (
            O => \N__3666\,
            I => \N__3663\
        );

    \I__576\ : Span4Mux_h
    port map (
            O => \N__3663\,
            I => \N__3660\
        );

    \I__575\ : Sp12to4
    port map (
            O => \N__3660\,
            I => \N__3657\
        );

    \I__574\ : Span12Mux_h
    port map (
            O => \N__3657\,
            I => \N__3654\
        );

    \I__573\ : Odrv12
    port map (
            O => \N__3654\,
            I => \D_UU_040_in_2\
        );

    \I__572\ : IoInMux
    port map (
            O => \N__3651\,
            I => \N__3647\
        );

    \I__571\ : InMux
    port map (
            O => \N__3650\,
            I => \N__3644\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3647\,
            I => \N__3641\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3644\,
            I => \N__3638\
        );

    \I__568\ : Span4Mux_s1_h
    port map (
            O => \N__3641\,
            I => \N__3635\
        );

    \I__567\ : Span4Mux_h
    port map (
            O => \N__3638\,
            I => \N__3632\
        );

    \I__566\ : Sp12to4
    port map (
            O => \N__3635\,
            I => \N__3629\
        );

    \I__565\ : Sp12to4
    port map (
            O => \N__3632\,
            I => \N__3626\
        );

    \I__564\ : Span12Mux_v
    port map (
            O => \N__3629\,
            I => \N__3623\
        );

    \I__563\ : Span12Mux_v
    port map (
            O => \N__3626\,
            I => \N__3620\
        );

    \I__562\ : Span12Mux_h
    port map (
            O => \N__3623\,
            I => \N__3615\
        );

    \I__561\ : Span12Mux_v
    port map (
            O => \N__3620\,
            I => \N__3615\
        );

    \I__560\ : Span12Mux_h
    port map (
            O => \N__3615\,
            I => \N__3612\
        );

    \I__559\ : Odrv12
    port map (
            O => \N__3612\,
            I => \D_LM_040_in_2\
        );

    \I__558\ : IoInMux
    port map (
            O => \N__3609\,
            I => \N__3606\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3606\,
            I => \N__3603\
        );

    \I__556\ : IoSpan4Mux
    port map (
            O => \N__3603\,
            I => \N__3600\
        );

    \I__555\ : Span4Mux_s2_v
    port map (
            O => \N__3600\,
            I => \N__3597\
        );

    \I__554\ : Span4Mux_v
    port map (
            O => \N__3597\,
            I => \N__3594\
        );

    \I__553\ : Odrv4
    port map (
            O => \N__3594\,
            I => \un1_D_UU_040_2\
        );

    \I__552\ : IoInMux
    port map (
            O => \N__3591\,
            I => \N__3588\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3588\,
            I => \N__3585\
        );

    \I__550\ : Span12Mux_s11_v
    port map (
            O => \N__3585\,
            I => \N__3582\
        );

    \I__549\ : Odrv12
    port map (
            O => \N__3582\,
            I => \CPUBGn_c_i_0\
        );

    \I__548\ : InMux
    port map (
            O => \N__3579\,
            I => \N__3576\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3576\,
            I => \N__3573\
        );

    \I__546\ : Span12Mux_v
    port map (
            O => \N__3573\,
            I => \N__3570\
        );

    \I__545\ : Odrv12
    port map (
            O => \N__3570\,
            I => \D_LL_AMIGA_in_7\
        );

    \I__544\ : IoInMux
    port map (
            O => \N__3567\,
            I => \N__3564\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3564\,
            I => \N__3561\
        );

    \I__542\ : Span12Mux_s8_h
    port map (
            O => \N__3561\,
            I => \N__3558\
        );

    \I__541\ : Span12Mux_h
    port map (
            O => \N__3558\,
            I => \N__3555\
        );

    \I__540\ : Odrv12
    port map (
            O => \N__3555\,
            I => \un2_D_LL_AMIGA_7\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__3552\,
            I => \U111_CYCLE_SM.N_112_cascade_\
        );

    \I__538\ : InMux
    port map (
            O => \N__3549\,
            I => \N__3546\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3546\,
            I => \N__3543\
        );

    \I__536\ : Span4Mux_v
    port map (
            O => \N__3543\,
            I => \N__3540\
        );

    \I__535\ : Sp12to4
    port map (
            O => \N__3540\,
            I => \N__3537\
        );

    \I__534\ : Odrv12
    port map (
            O => \N__3537\,
            I => \D_LL_AMIGA_in_2\
        );

    \I__533\ : IoInMux
    port map (
            O => \N__3534\,
            I => \N__3531\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3531\,
            I => \N__3528\
        );

    \I__531\ : IoSpan4Mux
    port map (
            O => \N__3528\,
            I => \N__3525\
        );

    \I__530\ : IoSpan4Mux
    port map (
            O => \N__3525\,
            I => \N__3522\
        );

    \I__529\ : Sp12to4
    port map (
            O => \N__3522\,
            I => \N__3519\
        );

    \I__528\ : Span12Mux_s9_h
    port map (
            O => \N__3519\,
            I => \N__3516\
        );

    \I__527\ : Span12Mux_h
    port map (
            O => \N__3516\,
            I => \N__3513\
        );

    \I__526\ : Odrv12
    port map (
            O => \N__3513\,
            I => \un2_D_LL_AMIGA_2\
        );

    \I__525\ : InMux
    port map (
            O => \N__3510\,
            I => \N__3507\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3507\,
            I => \N__3504\
        );

    \I__523\ : Span4Mux_v
    port map (
            O => \N__3504\,
            I => \N__3501\
        );

    \I__522\ : Sp12to4
    port map (
            O => \N__3501\,
            I => \N__3498\
        );

    \I__521\ : Odrv12
    port map (
            O => \N__3498\,
            I => \D_LL_AMIGA_in_3\
        );

    \I__520\ : IoInMux
    port map (
            O => \N__3495\,
            I => \N__3492\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3492\,
            I => \N__3489\
        );

    \I__518\ : Span4Mux_s2_h
    port map (
            O => \N__3489\,
            I => \N__3486\
        );

    \I__517\ : Span4Mux_v
    port map (
            O => \N__3486\,
            I => \N__3483\
        );

    \I__516\ : Span4Mux_v
    port map (
            O => \N__3483\,
            I => \N__3480\
        );

    \I__515\ : Sp12to4
    port map (
            O => \N__3480\,
            I => \N__3477\
        );

    \I__514\ : Span12Mux_s11_h
    port map (
            O => \N__3477\,
            I => \N__3474\
        );

    \I__513\ : Odrv12
    port map (
            O => \N__3474\,
            I => \un2_D_LL_AMIGA_3\
        );

    \I__512\ : InMux
    port map (
            O => \N__3471\,
            I => \N__3468\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3468\,
            I => \N__3465\
        );

    \I__510\ : Span4Mux_v
    port map (
            O => \N__3465\,
            I => \N__3462\
        );

    \I__509\ : Span4Mux_v
    port map (
            O => \N__3462\,
            I => \N__3458\
        );

    \I__508\ : InMux
    port map (
            O => \N__3461\,
            I => \N__3455\
        );

    \I__507\ : Sp12to4
    port map (
            O => \N__3458\,
            I => \N__3450\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3455\,
            I => \N__3450\
        );

    \I__505\ : Span12Mux_h
    port map (
            O => \N__3450\,
            I => \N__3447\
        );

    \I__504\ : Odrv12
    port map (
            O => \N__3447\,
            I => \A_040_c_1\
        );

    \I__503\ : InMux
    port map (
            O => \N__3444\,
            I => \N__3441\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3441\,
            I => \N__3438\
        );

    \I__501\ : Span4Mux_v
    port map (
            O => \N__3438\,
            I => \N__3435\
        );

    \I__500\ : Sp12to4
    port map (
            O => \N__3435\,
            I => \N__3432\
        );

    \I__499\ : Odrv12
    port map (
            O => \N__3432\,
            I => \D_LM_AMIGA_in_0\
        );

    \I__498\ : IoInMux
    port map (
            O => \N__3429\,
            I => \N__3426\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3426\,
            I => \N__3423\
        );

    \I__496\ : Span4Mux_s2_h
    port map (
            O => \N__3423\,
            I => \N__3420\
        );

    \I__495\ : Span4Mux_v
    port map (
            O => \N__3420\,
            I => \N__3417\
        );

    \I__494\ : Span4Mux_v
    port map (
            O => \N__3417\,
            I => \N__3414\
        );

    \I__493\ : Sp12to4
    port map (
            O => \N__3414\,
            I => \N__3411\
        );

    \I__492\ : Span12Mux_s11_h
    port map (
            O => \N__3411\,
            I => \N__3408\
        );

    \I__491\ : Odrv12
    port map (
            O => \N__3408\,
            I => \N_122\
        );

    \I__490\ : InMux
    port map (
            O => \N__3405\,
            I => \N__3399\
        );

    \I__489\ : InMux
    port map (
            O => \N__3404\,
            I => \N__3399\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3399\,
            I => \N__3396\
        );

    \I__487\ : Span4Mux_v
    port map (
            O => \N__3396\,
            I => \N__3393\
        );

    \I__486\ : Span4Mux_v
    port map (
            O => \N__3393\,
            I => \N__3390\
        );

    \I__485\ : Span4Mux_h
    port map (
            O => \N__3390\,
            I => \N__3386\
        );

    \I__484\ : InMux
    port map (
            O => \N__3389\,
            I => \N__3383\
        );

    \I__483\ : Odrv4
    port map (
            O => \N__3386\,
            I => \U111_CYCLE_SM.A2_ENZ0\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3383\,
            I => \U111_CYCLE_SM.A2_ENZ0\
        );

    \I__481\ : CascadeMux
    port map (
            O => \N__3378\,
            I => \N__3375\
        );

    \I__480\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3372\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3372\,
            I => \N__3369\
        );

    \I__478\ : Odrv4
    port map (
            O => \N__3369\,
            I => \U111_CYCLE_SM.N_151\
        );

    \I__477\ : InMux
    port map (
            O => \N__3366\,
            I => \N__3363\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3363\,
            I => \N__3360\
        );

    \I__475\ : Span4Mux_v
    port map (
            O => \N__3360\,
            I => \N__3357\
        );

    \I__474\ : Sp12to4
    port map (
            O => \N__3357\,
            I => \N__3354\
        );

    \I__473\ : Span12Mux_h
    port map (
            O => \N__3354\,
            I => \N__3351\
        );

    \I__472\ : Span12Mux_h
    port map (
            O => \N__3351\,
            I => \N__3348\
        );

    \I__471\ : Span12Mux_v
    port map (
            O => \N__3348\,
            I => \N__3345\
        );

    \I__470\ : Odrv12
    port map (
            O => \N__3345\,
            I => \D_UM_040_in_1\
        );

    \I__469\ : InMux
    port map (
            O => \N__3342\,
            I => \N__3338\
        );

    \I__468\ : IoInMux
    port map (
            O => \N__3341\,
            I => \N__3335\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3338\,
            I => \N__3332\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3335\,
            I => \N__3329\
        );

    \I__465\ : Span4Mux_v
    port map (
            O => \N__3332\,
            I => \N__3326\
        );

    \I__464\ : Span4Mux_s3_h
    port map (
            O => \N__3329\,
            I => \N__3323\
        );

    \I__463\ : Span4Mux_v
    port map (
            O => \N__3326\,
            I => \N__3320\
        );

    \I__462\ : Sp12to4
    port map (
            O => \N__3323\,
            I => \N__3317\
        );

    \I__461\ : Sp12to4
    port map (
            O => \N__3320\,
            I => \N__3314\
        );

    \I__460\ : Span12Mux_v
    port map (
            O => \N__3317\,
            I => \N__3311\
        );

    \I__459\ : Span12Mux_v
    port map (
            O => \N__3314\,
            I => \N__3308\
        );

    \I__458\ : Span12Mux_h
    port map (
            O => \N__3311\,
            I => \N__3305\
        );

    \I__457\ : Span12Mux_h
    port map (
            O => \N__3308\,
            I => \N__3302\
        );

    \I__456\ : Span12Mux_h
    port map (
            O => \N__3305\,
            I => \N__3299\
        );

    \I__455\ : Odrv12
    port map (
            O => \N__3302\,
            I => \D_LL_040_in_1\
        );

    \I__454\ : Odrv12
    port map (
            O => \N__3299\,
            I => \D_LL_040_in_1\
        );

    \I__453\ : IoInMux
    port map (
            O => \N__3294\,
            I => \N__3291\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3291\,
            I => \N__3288\
        );

    \I__451\ : Span12Mux_s10_h
    port map (
            O => \N__3288\,
            I => \N__3285\
        );

    \I__450\ : Odrv12
    port map (
            O => \N__3285\,
            I => \un1_D_UM_040_1\
        );

    \I__449\ : InMux
    port map (
            O => \N__3282\,
            I => \N__3279\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3279\,
            I => \N__3276\
        );

    \I__447\ : Span4Mux_v
    port map (
            O => \N__3276\,
            I => \N__3273\
        );

    \I__446\ : Sp12to4
    port map (
            O => \N__3273\,
            I => \N__3270\
        );

    \I__445\ : Span12Mux_h
    port map (
            O => \N__3270\,
            I => \N__3267\
        );

    \I__444\ : Odrv12
    port map (
            O => \N__3267\,
            I => \D_UM_040_in_0\
        );

    \I__443\ : IoInMux
    port map (
            O => \N__3264\,
            I => \N__3261\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__3261\,
            I => \N__3257\
        );

    \I__441\ : InMux
    port map (
            O => \N__3260\,
            I => \N__3254\
        );

    \I__440\ : IoSpan4Mux
    port map (
            O => \N__3257\,
            I => \N__3251\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3254\,
            I => \N__3248\
        );

    \I__438\ : Span4Mux_s2_h
    port map (
            O => \N__3251\,
            I => \N__3245\
        );

    \I__437\ : Span12Mux_v
    port map (
            O => \N__3248\,
            I => \N__3242\
        );

    \I__436\ : Sp12to4
    port map (
            O => \N__3245\,
            I => \N__3239\
        );

    \I__435\ : Span12Mux_v
    port map (
            O => \N__3242\,
            I => \N__3236\
        );

    \I__434\ : Span12Mux_h
    port map (
            O => \N__3239\,
            I => \N__3233\
        );

    \I__433\ : Span12Mux_h
    port map (
            O => \N__3236\,
            I => \N__3230\
        );

    \I__432\ : Span12Mux_h
    port map (
            O => \N__3233\,
            I => \N__3227\
        );

    \I__431\ : Odrv12
    port map (
            O => \N__3230\,
            I => \D_LL_040_in_0\
        );

    \I__430\ : Odrv12
    port map (
            O => \N__3227\,
            I => \D_LL_040_in_0\
        );

    \I__429\ : IoInMux
    port map (
            O => \N__3222\,
            I => \N__3219\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3219\,
            I => \N__3216\
        );

    \I__427\ : IoSpan4Mux
    port map (
            O => \N__3216\,
            I => \N__3213\
        );

    \I__426\ : Span4Mux_s3_h
    port map (
            O => \N__3213\,
            I => \N__3210\
        );

    \I__425\ : Span4Mux_h
    port map (
            O => \N__3210\,
            I => \N__3207\
        );

    \I__424\ : Odrv4
    port map (
            O => \N__3207\,
            I => \un1_D_UM_040_0\
        );

    \I__423\ : InMux
    port map (
            O => \N__3204\,
            I => \N__3201\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3201\,
            I => \N__3198\
        );

    \I__421\ : Span4Mux_v
    port map (
            O => \N__3198\,
            I => \N__3195\
        );

    \I__420\ : Sp12to4
    port map (
            O => \N__3195\,
            I => \N__3192\
        );

    \I__419\ : Odrv12
    port map (
            O => \N__3192\,
            I => \D_LM_AMIGA_in_3\
        );

    \I__418\ : IoInMux
    port map (
            O => \N__3189\,
            I => \N__3186\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3186\,
            I => \N__3183\
        );

    \I__416\ : IoSpan4Mux
    port map (
            O => \N__3183\,
            I => \N__3180\
        );

    \I__415\ : Span4Mux_s1_h
    port map (
            O => \N__3180\,
            I => \N__3177\
        );

    \I__414\ : Span4Mux_v
    port map (
            O => \N__3177\,
            I => \N__3174\
        );

    \I__413\ : Sp12to4
    port map (
            O => \N__3174\,
            I => \N__3171\
        );

    \I__412\ : Span12Mux_s10_h
    port map (
            O => \N__3171\,
            I => \N__3168\
        );

    \I__411\ : Odrv12
    port map (
            O => \N__3168\,
            I => \N_119\
        );

    \I__410\ : InMux
    port map (
            O => \N__3165\,
            I => \N__3162\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3162\,
            I => \N__3159\
        );

    \I__408\ : Odrv12
    port map (
            O => \N__3159\,
            I => \D_LM_AMIGA_in_1\
        );

    \I__407\ : IoInMux
    port map (
            O => \N__3156\,
            I => \N__3153\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3153\,
            I => \N__3150\
        );

    \I__405\ : Span4Mux_s0_h
    port map (
            O => \N__3150\,
            I => \N__3147\
        );

    \I__404\ : Sp12to4
    port map (
            O => \N__3147\,
            I => \N__3144\
        );

    \I__403\ : Span12Mux_v
    port map (
            O => \N__3144\,
            I => \N__3141\
        );

    \I__402\ : Span12Mux_h
    port map (
            O => \N__3141\,
            I => \N__3138\
        );

    \I__401\ : Odrv12
    port map (
            O => \N__3138\,
            I => \N_121\
        );

    \I__400\ : IoInMux
    port map (
            O => \N__3135\,
            I => \N__3132\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3132\,
            I => \N__3128\
        );

    \I__398\ : InMux
    port map (
            O => \N__3131\,
            I => \N__3125\
        );

    \I__397\ : IoSpan4Mux
    port map (
            O => \N__3128\,
            I => \N__3122\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3125\,
            I => \N__3119\
        );

    \I__395\ : Span4Mux_s0_h
    port map (
            O => \N__3122\,
            I => \N__3116\
        );

    \I__394\ : Span4Mux_v
    port map (
            O => \N__3119\,
            I => \N__3113\
        );

    \I__393\ : Span4Mux_v
    port map (
            O => \N__3116\,
            I => \N__3110\
        );

    \I__392\ : Sp12to4
    port map (
            O => \N__3113\,
            I => \N__3107\
        );

    \I__391\ : Sp12to4
    port map (
            O => \N__3110\,
            I => \N__3104\
        );

    \I__390\ : Span12Mux_h
    port map (
            O => \N__3107\,
            I => \N__3101\
        );

    \I__389\ : Span12Mux_h
    port map (
            O => \N__3104\,
            I => \N__3098\
        );

    \I__388\ : Span12Mux_v
    port map (
            O => \N__3101\,
            I => \N__3095\
        );

    \I__387\ : Span12Mux_h
    port map (
            O => \N__3098\,
            I => \N__3092\
        );

    \I__386\ : Span12Mux_h
    port map (
            O => \N__3095\,
            I => \N__3089\
        );

    \I__385\ : Odrv12
    port map (
            O => \N__3092\,
            I => \D_LL_040_in_6\
        );

    \I__384\ : Odrv12
    port map (
            O => \N__3089\,
            I => \D_LL_040_in_6\
        );

    \I__383\ : InMux
    port map (
            O => \N__3084\,
            I => \N__3081\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3081\,
            I => \N__3078\
        );

    \I__381\ : Span12Mux_v
    port map (
            O => \N__3078\,
            I => \N__3075\
        );

    \I__380\ : Span12Mux_h
    port map (
            O => \N__3075\,
            I => \N__3072\
        );

    \I__379\ : Odrv12
    port map (
            O => \N__3072\,
            I => \D_UM_040_in_6\
        );

    \I__378\ : IoInMux
    port map (
            O => \N__3069\,
            I => \N__3066\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__3066\,
            I => \N__3063\
        );

    \I__376\ : Span12Mux_s4_h
    port map (
            O => \N__3063\,
            I => \N__3060\
        );

    \I__375\ : Span12Mux_v
    port map (
            O => \N__3060\,
            I => \N__3057\
        );

    \I__374\ : Odrv12
    port map (
            O => \N__3057\,
            I => \un1_D_UM_040_6\
        );

    \I__373\ : InMux
    port map (
            O => \N__3054\,
            I => \N__3051\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3051\,
            I => \N__3048\
        );

    \I__371\ : Odrv12
    port map (
            O => \N__3048\,
            I => \D_LM_AMIGA_in_2\
        );

    \I__370\ : IoInMux
    port map (
            O => \N__3045\,
            I => \N__3042\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3042\,
            I => \N__3039\
        );

    \I__368\ : Span12Mux_s11_h
    port map (
            O => \N__3039\,
            I => \N__3036\
        );

    \I__367\ : Span12Mux_v
    port map (
            O => \N__3036\,
            I => \N__3033\
        );

    \I__366\ : Odrv12
    port map (
            O => \N__3033\,
            I => \N_120\
        );

    \I__365\ : IoInMux
    port map (
            O => \N__3030\,
            I => \N__3027\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3027\,
            I => \N__3024\
        );

    \I__363\ : IoSpan4Mux
    port map (
            O => \N__3024\,
            I => \N__3020\
        );

    \I__362\ : InMux
    port map (
            O => \N__3023\,
            I => \N__3017\
        );

    \I__361\ : IoSpan4Mux
    port map (
            O => \N__3020\,
            I => \N__3014\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3017\,
            I => \N__3011\
        );

    \I__359\ : Span4Mux_s2_h
    port map (
            O => \N__3014\,
            I => \N__3008\
        );

    \I__358\ : Span12Mux_v
    port map (
            O => \N__3011\,
            I => \N__3005\
        );

    \I__357\ : Sp12to4
    port map (
            O => \N__3008\,
            I => \N__3002\
        );

    \I__356\ : Span12Mux_v
    port map (
            O => \N__3005\,
            I => \N__2999\
        );

    \I__355\ : Span12Mux_h
    port map (
            O => \N__3002\,
            I => \N__2996\
        );

    \I__354\ : Span12Mux_h
    port map (
            O => \N__2999\,
            I => \N__2993\
        );

    \I__353\ : Span12Mux_h
    port map (
            O => \N__2996\,
            I => \N__2990\
        );

    \I__352\ : Odrv12
    port map (
            O => \N__2993\,
            I => \D_LM_040_in_0\
        );

    \I__351\ : Odrv12
    port map (
            O => \N__2990\,
            I => \D_LM_040_in_0\
        );

    \I__350\ : InMux
    port map (
            O => \N__2985\,
            I => \N__2982\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2982\,
            I => \N__2979\
        );

    \I__348\ : Span4Mux_v
    port map (
            O => \N__2979\,
            I => \N__2976\
        );

    \I__347\ : Span4Mux_h
    port map (
            O => \N__2976\,
            I => \N__2973\
        );

    \I__346\ : Sp12to4
    port map (
            O => \N__2973\,
            I => \N__2970\
        );

    \I__345\ : Span12Mux_h
    port map (
            O => \N__2970\,
            I => \N__2967\
        );

    \I__344\ : Odrv12
    port map (
            O => \N__2967\,
            I => \D_UU_040_in_0\
        );

    \I__343\ : IoInMux
    port map (
            O => \N__2964\,
            I => \N__2961\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2961\,
            I => \N__2958\
        );

    \I__341\ : IoSpan4Mux
    port map (
            O => \N__2958\,
            I => \N__2955\
        );

    \I__340\ : Span4Mux_s2_v
    port map (
            O => \N__2955\,
            I => \N__2952\
        );

    \I__339\ : Span4Mux_v
    port map (
            O => \N__2952\,
            I => \N__2949\
        );

    \I__338\ : Odrv4
    port map (
            O => \N__2949\,
            I => \un1_D_UU_040_0\
        );

    \I__337\ : InMux
    port map (
            O => \N__2946\,
            I => \N__2943\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2943\,
            I => \N__2940\
        );

    \I__335\ : Span4Mux_v
    port map (
            O => \N__2940\,
            I => \N__2937\
        );

    \I__334\ : Span4Mux_h
    port map (
            O => \N__2937\,
            I => \N__2934\
        );

    \I__333\ : Sp12to4
    port map (
            O => \N__2934\,
            I => \N__2931\
        );

    \I__332\ : Span12Mux_h
    port map (
            O => \N__2931\,
            I => \N__2928\
        );

    \I__331\ : Odrv12
    port map (
            O => \N__2928\,
            I => \D_UU_040_in_4\
        );

    \I__330\ : IoInMux
    port map (
            O => \N__2925\,
            I => \N__2922\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2922\,
            I => \N__2919\
        );

    \I__328\ : Span4Mux_s1_h
    port map (
            O => \N__2919\,
            I => \N__2916\
        );

    \I__327\ : Sp12to4
    port map (
            O => \N__2916\,
            I => \N__2912\
        );

    \I__326\ : InMux
    port map (
            O => \N__2915\,
            I => \N__2909\
        );

    \I__325\ : Span12Mux_v
    port map (
            O => \N__2912\,
            I => \N__2906\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__2909\,
            I => \N__2903\
        );

    \I__323\ : Span12Mux_h
    port map (
            O => \N__2906\,
            I => \N__2900\
        );

    \I__322\ : Span12Mux_v
    port map (
            O => \N__2903\,
            I => \N__2897\
        );

    \I__321\ : Span12Mux_h
    port map (
            O => \N__2900\,
            I => \N__2894\
        );

    \I__320\ : Span12Mux_h
    port map (
            O => \N__2897\,
            I => \N__2891\
        );

    \I__319\ : Odrv12
    port map (
            O => \N__2894\,
            I => \D_LM_040_in_4\
        );

    \I__318\ : Odrv12
    port map (
            O => \N__2891\,
            I => \D_LM_040_in_4\
        );

    \I__317\ : IoInMux
    port map (
            O => \N__2886\,
            I => \N__2883\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2883\,
            I => \N__2880\
        );

    \I__315\ : IoSpan4Mux
    port map (
            O => \N__2880\,
            I => \N__2877\
        );

    \I__314\ : Span4Mux_s3_v
    port map (
            O => \N__2877\,
            I => \N__2874\
        );

    \I__313\ : Odrv4
    port map (
            O => \N__2874\,
            I => \un1_D_UU_040_4\
        );

    \I__312\ : InMux
    port map (
            O => \N__2871\,
            I => \N__2868\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2868\,
            I => \N__2865\
        );

    \I__310\ : Span4Mux_v
    port map (
            O => \N__2865\,
            I => \N__2862\
        );

    \I__309\ : Sp12to4
    port map (
            O => \N__2862\,
            I => \N__2859\
        );

    \I__308\ : Span12Mux_h
    port map (
            O => \N__2859\,
            I => \N__2856\
        );

    \I__307\ : Span12Mux_h
    port map (
            O => \N__2856\,
            I => \N__2853\
        );

    \I__306\ : Odrv12
    port map (
            O => \N__2853\,
            I => \D_UU_040_in_6\
        );

    \I__305\ : IoInMux
    port map (
            O => \N__2850\,
            I => \N__2847\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2847\,
            I => \N__2844\
        );

    \I__303\ : Span4Mux_s2_h
    port map (
            O => \N__2844\,
            I => \N__2840\
        );

    \I__302\ : InMux
    port map (
            O => \N__2843\,
            I => \N__2837\
        );

    \I__301\ : Span4Mux_h
    port map (
            O => \N__2840\,
            I => \N__2834\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2837\,
            I => \N__2831\
        );

    \I__299\ : Span4Mux_h
    port map (
            O => \N__2834\,
            I => \N__2826\
        );

    \I__298\ : Span4Mux_v
    port map (
            O => \N__2831\,
            I => \N__2826\
        );

    \I__297\ : Span4Mux_v
    port map (
            O => \N__2826\,
            I => \N__2823\
        );

    \I__296\ : Sp12to4
    port map (
            O => \N__2823\,
            I => \N__2820\
        );

    \I__295\ : Span12Mux_h
    port map (
            O => \N__2820\,
            I => \N__2817\
        );

    \I__294\ : Span12Mux_h
    port map (
            O => \N__2817\,
            I => \N__2814\
        );

    \I__293\ : Odrv12
    port map (
            O => \N__2814\,
            I => \D_LM_040_in_6\
        );

    \I__292\ : IoInMux
    port map (
            O => \N__2811\,
            I => \N__2808\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2808\,
            I => \N__2805\
        );

    \I__290\ : Span4Mux_s2_v
    port map (
            O => \N__2805\,
            I => \N__2802\
        );

    \I__289\ : Span4Mux_h
    port map (
            O => \N__2802\,
            I => \N__2799\
        );

    \I__288\ : Span4Mux_v
    port map (
            O => \N__2799\,
            I => \N__2796\
        );

    \I__287\ : Odrv4
    port map (
            O => \N__2796\,
            I => \un1_D_UU_040_6\
        );

    \I__286\ : IoInMux
    port map (
            O => \N__2793\,
            I => \N__2790\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2790\,
            I => \N__2787\
        );

    \I__284\ : Span4Mux_s0_v
    port map (
            O => \N__2787\,
            I => \N__2784\
        );

    \I__283\ : Sp12to4
    port map (
            O => \N__2784\,
            I => \N__2781\
        );

    \I__282\ : Span12Mux_h
    port map (
            O => \N__2781\,
            I => \N__2778\
        );

    \I__281\ : Span12Mux_v
    port map (
            O => \N__2778\,
            I => \N__2775\
        );

    \I__280\ : Span12Mux_v
    port map (
            O => \N__2775\,
            I => \N__2772\
        );

    \I__279\ : Odrv12
    port map (
            O => \N__2772\,
            I => \TAn_in\
        );

    \I__278\ : IoInMux
    port map (
            O => \N__2769\,
            I => \N__2766\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2766\,
            I => \N__2763\
        );

    \I__276\ : Odrv12
    port map (
            O => \N__2763\,
            I => \RESETn_c_i\
        );

    \I__275\ : IoInMux
    port map (
            O => \N__2760\,
            I => \N__2757\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2757\,
            I => \N__2754\
        );

    \I__273\ : Odrv12
    port map (
            O => \N__2754\,
            I => \U111_CYCLE_SM_A_AMIGA_0_i_1\
        );

    \I__272\ : InMux
    port map (
            O => \N__2751\,
            I => \N__2748\
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2748\,
            I => \N__2745\
        );

    \I__270\ : Span4Mux_h
    port map (
            O => \N__2745\,
            I => \N__2742\
        );

    \I__269\ : Span4Mux_v
    port map (
            O => \N__2742\,
            I => \N__2739\
        );

    \I__268\ : Odrv4
    port map (
            O => \N__2739\,
            I => \A_040_c_0\
        );

    \I__267\ : IoInMux
    port map (
            O => \N__2736\,
            I => \N__2733\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2733\,
            I => \N__2730\
        );

    \I__265\ : Span4Mux_s2_v
    port map (
            O => \N__2730\,
            I => \N__2727\
        );

    \I__264\ : Span4Mux_v
    port map (
            O => \N__2727\,
            I => \N__2724\
        );

    \I__263\ : Odrv4
    port map (
            O => \N__2724\,
            I => \A_AMIGA_c_0\
        );

    \I__262\ : InMux
    port map (
            O => \N__2721\,
            I => \N__2718\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2718\,
            I => \N__2715\
        );

    \I__260\ : Span4Mux_v
    port map (
            O => \N__2715\,
            I => \N__2712\
        );

    \I__259\ : Sp12to4
    port map (
            O => \N__2712\,
            I => \N__2709\
        );

    \I__258\ : Odrv12
    port map (
            O => \N__2709\,
            I => \D_LL_AMIGA_in_4\
        );

    \I__257\ : IoInMux
    port map (
            O => \N__2706\,
            I => \N__2703\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__2703\,
            I => \N__2700\
        );

    \I__255\ : Span4Mux_s3_h
    port map (
            O => \N__2700\,
            I => \N__2697\
        );

    \I__254\ : Sp12to4
    port map (
            O => \N__2697\,
            I => \N__2694\
        );

    \I__253\ : Span12Mux_s8_v
    port map (
            O => \N__2694\,
            I => \N__2691\
        );

    \I__252\ : Span12Mux_h
    port map (
            O => \N__2691\,
            I => \N__2688\
        );

    \I__251\ : Odrv12
    port map (
            O => \N__2688\,
            I => \un2_D_LL_AMIGA_4\
        );

    \I__250\ : InMux
    port map (
            O => \N__2685\,
            I => \N__2682\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2682\,
            I => \N__2679\
        );

    \I__248\ : Span12Mux_v
    port map (
            O => \N__2679\,
            I => \N__2676\
        );

    \I__247\ : Odrv12
    port map (
            O => \N__2676\,
            I => \D_LL_AMIGA_in_1\
        );

    \I__246\ : IoInMux
    port map (
            O => \N__2673\,
            I => \N__2670\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2670\,
            I => \N__2667\
        );

    \I__244\ : IoSpan4Mux
    port map (
            O => \N__2667\,
            I => \N__2664\
        );

    \I__243\ : Span4Mux_s1_h
    port map (
            O => \N__2664\,
            I => \N__2661\
        );

    \I__242\ : Span4Mux_v
    port map (
            O => \N__2661\,
            I => \N__2658\
        );

    \I__241\ : Sp12to4
    port map (
            O => \N__2658\,
            I => \N__2655\
        );

    \I__240\ : Span12Mux_s10_h
    port map (
            O => \N__2655\,
            I => \N__2652\
        );

    \I__239\ : Odrv12
    port map (
            O => \N__2652\,
            I => \un2_D_LL_AMIGA_1\
        );

    \I__238\ : IoInMux
    port map (
            O => \N__2649\,
            I => \N__2646\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__2646\,
            I => \N__2643\
        );

    \I__236\ : Span4Mux_s1_v
    port map (
            O => \N__2643\,
            I => \N__2640\
        );

    \I__235\ : Span4Mux_v
    port map (
            O => \N__2640\,
            I => \N__2637\
        );

    \I__234\ : Sp12to4
    port map (
            O => \N__2637\,
            I => \N__2634\
        );

    \I__233\ : Span12Mux_h
    port map (
            O => \N__2634\,
            I => \N__2631\
        );

    \I__232\ : Span12Mux_v
    port map (
            O => \N__2631\,
            I => \N__2628\
        );

    \I__231\ : Span12Mux_v
    port map (
            O => \N__2628\,
            I => \N__2625\
        );

    \I__230\ : Odrv12
    port map (
            O => \N__2625\,
            I => \TSn_in\
        );

    \I__229\ : IoInMux
    port map (
            O => \N__2622\,
            I => \N__2619\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__2619\,
            I => \N__2616\
        );

    \I__227\ : Span4Mux_s0_h
    port map (
            O => \N__2616\,
            I => \N__2613\
        );

    \I__226\ : Span4Mux_h
    port map (
            O => \N__2613\,
            I => \N__2610\
        );

    \I__225\ : Span4Mux_h
    port map (
            O => \N__2610\,
            I => \N__2607\
        );

    \I__224\ : Sp12to4
    port map (
            O => \N__2607\,
            I => \N__2604\
        );

    \I__223\ : Span12Mux_s11_v
    port map (
            O => \N__2604\,
            I => \N__2601\
        );

    \I__222\ : Span12Mux_v
    port map (
            O => \N__2601\,
            I => \N__2598\
        );

    \I__221\ : Span12Mux_h
    port map (
            O => \N__2598\,
            I => \N__2595\
        );

    \I__220\ : Odrv12
    port map (
            O => \N__2595\,
            I => \TCIn_c\
        );

    \INVU111_CYCLE_SM.TS_OUTC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TS_OUTC_net\,
            I => \N__6381\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2769\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4645\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_RNIB97G_LC_3_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3461\,
            in2 => \_gnd_net_\,
            in3 => \N__3405\,
            lcout => \U111_CYCLE_SM_A_AMIGA_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_RNIA87G_LC_3_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__2751\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3404\,
            lcout => \A_AMIGA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI6HT71_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2721\,
            in1 => \N__7585\,
            in2 => \_gnd_net_\,
            in3 => \N__7894\,
            lcout => \un2_D_LL_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI0BT71_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7893\,
            in1 => \N__4399\,
            in2 => \_gnd_net_\,
            in3 => \N__2685\,
            lcout => \un2_D_LL_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI8QN01_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3282\,
            in1 => \N__3260\,
            in2 => \_gnd_net_\,
            in3 => \N__7751\,
            lcout => \un1_D_UM_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIDMI41_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7753\,
            in1 => \N__4229\,
            in2 => \_gnd_net_\,
            in3 => \N__3204\,
            lcout => \N_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI9II41_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7752\,
            in1 => \N__6299\,
            in2 => \_gnd_net_\,
            in3 => \N__3165\,
            lcout => \N_121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIK6O01_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7818\,
            in1 => \N__3131\,
            in2 => \_gnd_net_\,
            in3 => \N__3084\,
            lcout => \un1_D_UM_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIBKI41_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7817\,
            in1 => \N__3752\,
            in2 => \_gnd_net_\,
            in3 => \N__3054\,
            lcout => \N_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIHFPK_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__3023\,
            in1 => \N__2985\,
            in2 => \_gnd_net_\,
            in3 => \N__7895\,
            lcout => \un1_D_UU_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIPNPK_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7896\,
            in1 => \N__2946\,
            in2 => \_gnd_net_\,
            in3 => \N__2915\,
            lcout => \un1_D_UU_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNITRPK_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2871\,
            in1 => \N__2843\,
            in2 => \_gnd_net_\,
            in3 => \N__7897\,
            lcout => \un1_D_UU_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI2DT71_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3549\,
            in1 => \N__6720\,
            in2 => \_gnd_net_\,
            in3 => \N__7851\,
            lcout => \un2_D_LL_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI4FT71_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7852\,
            in1 => \N__6080\,
            in2 => \_gnd_net_\,
            in3 => \N__3510\,
            lcout => \un2_D_LL_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNO_0_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4960\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3471\,
            lcout => \U111_CYCLE_SM.N_151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI7GI41_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7805\,
            in1 => \N__6204\,
            in2 => \_gnd_net_\,
            in3 => \N__3444\,
            lcout => \N_122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A2_EN_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__3389\,
            in1 => \N__3927\,
            in2 => \_gnd_net_\,
            in3 => \N__5121\,
            lcout => \U111_CYCLE_SM.A2_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6385\,
            ce => 'H',
            sr => \N__6331\
        );

    \U111_CYCLE_SM.PORT_MISMATCH_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__3990\,
            in1 => \N__6417\,
            in2 => \N__4977\,
            in3 => \N__5089\,
            lcout => \U111_CYCLE_SM.PORT_MISMATCHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6385\,
            ce => 'H',
            sr => \N__6331\
        );

    \U111_CYCLE_SM.FLIP_WORD_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__5122\,
            in1 => \N__7750\,
            in2 => \N__3378\,
            in3 => \N__5088\,
            lcout => \U111_CYCLE_SM.FLIP_WORDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6385\,
            ce => 'H',
            sr => \N__6331\
        );

    \U111_CYCLE_SM.UU_LATCHED_2_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__3707\,
            in1 => \N__6606\,
            in2 => \N__3759\,
            in3 => \N__7191\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6382\,
            ce => 'H',
            sr => \N__6332\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIASN01_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3366\,
            in1 => \N__3342\,
            in2 => \_gnd_net_\,
            in3 => \N__7806\,
            lcout => \un1_D_UM_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIE0O01_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7807\,
            in1 => \N__3882\,
            in2 => \_gnd_net_\,
            in3 => \N__3837\,
            lcout => \un1_D_UM_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNILUI41_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7808\,
            in1 => \N__5527\,
            in2 => \_gnd_net_\,
            in3 => \N__3795\,
            lcout => \N_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNINJKT_2_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8421\,
            in1 => \N__3751\,
            in2 => \_gnd_net_\,
            in3 => \N__3711\,
            lcout => \N_129\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNILJPK_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3672\,
            in1 => \N__3650\,
            in2 => \_gnd_net_\,
            in3 => \N__7909\,
            lcout => \un1_D_UU_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TSn_iobuf_RNO_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7230\,
            lcout => \CPUBGn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNICNT71_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7871\,
            in1 => \N__5049\,
            in2 => \_gnd_net_\,
            in3 => \N__3579\,
            lcout => \un2_D_LL_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_5_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5350\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3914\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_5_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__4490\,
            in1 => \N__4641\,
            in2 => \N__3552\,
            in3 => \N__4124\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_0_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__5351\,
            in1 => \N__5114\,
            in2 => \N__4519\,
            in3 => \N__3913\,
            lcout => \U111_CYCLE_SM.N_132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_4_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5115\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4640\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_1_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__4643\,
            in1 => \N__3926\,
            in2 => \N__6465\,
            in3 => \N__4045\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_1_0_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__3988\,
            in1 => \N__4569\,
            in2 => \N__4547\,
            in3 => \N__3999\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_0_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__4642\,
            in1 => \N__3933\,
            in2 => \N__3936\,
            in3 => \N__3888\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__5381\,
            in1 => \N__4568\,
            in2 => \_gnd_net_\,
            in3 => \N__3912\,
            lcout => \U111_CYCLE_SM.N_142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_3_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4644\,
            in1 => \N__3989\,
            in2 => \_gnd_net_\,
            in3 => \N__4587\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIJG6K_5_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__4538\,
            in1 => \N__5380\,
            in2 => \_gnd_net_\,
            in3 => \N__3911\,
            lcout => \U111_CYCLE_SM.N_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_RNILNBJ_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3915\,
            in3 => \N__4044\,
            lcout => \U111_CYCLE_SM.N_195\,
            ltout => \U111_CYCLE_SM.N_195_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_2_0_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__4542\,
            in1 => \N__6628\,
            in2 => \N__3891\,
            in3 => \N__5800\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_srsts_0_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.BURST_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__6534\,
            in1 => \N__6498\,
            in2 => \N__6464\,
            in3 => \N__4047\,
            lcout => \U111_CYCLE_SM.BURSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6380\,
            ce => 'H',
            sr => \N__6333\
        );

    \U111_CYCLE_SM.BURST_COUNT_1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100000010"
        )
    port map (
            in0 => \N__4027\,
            in1 => \N__4586\,
            in2 => \N__6463\,
            in3 => \N__4011\,
            lcout => \U111_CYCLE_SM.BURST_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6380\,
            ce => 'H',
            sr => \N__6333\
        );

    \U111_CYCLE_SM.BURST_COUNT_0_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__6453\,
            in1 => \N__4585\,
            in2 => \_gnd_net_\,
            in3 => \N__4028\,
            lcout => \U111_CYCLE_SM.BURST_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6380\,
            ce => 'H',
            sr => \N__6333\
        );

    \U111_CYCLE_SM.BURST_COUNT_RNIFDQV_1_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101110111"
        )
    port map (
            in0 => \N__4080\,
            in1 => \N__4046\,
            in2 => \N__4029\,
            in3 => \N__4010\,
            lcout => \U111_CYCLE_SM.N_109\,
            ltout => \U111_CYCLE_SM.N_109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_1_2_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010000"
        )
    port map (
            in0 => \N__4543\,
            in1 => \N__5087\,
            in2 => \N__3993\,
            in3 => \N__3987\,
            lcout => \U111_CYCLE_SM.N_140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_1_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__4358\,
            in1 => \N__6600\,
            in2 => \N__4407\,
            in3 => \N__7188\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6377\,
            ce => 'H',
            sr => \N__6335\
        );

    \U111_CYCLE_SM.UM_LATCHED_4_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7189\,
            in1 => \N__7601\,
            in2 => \N__7590\,
            in3 => \N__6602\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6377\,
            ce => 'H',
            sr => \N__6335\
        );

    \U111_CYCLE_SM.UU_LATCHED_3_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__4169\,
            in1 => \N__6601\,
            in2 => \N__4230\,
            in3 => \N__7190\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6377\,
            ce => 'H',
            sr => \N__6335\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIHQI41_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7840\,
            in1 => \N__5618\,
            in2 => \_gnd_net_\,
            in3 => \N__3969\,
            lcout => \N_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIFOI41_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4443\,
            in1 => \N__5444\,
            in2 => \_gnd_net_\,
            in3 => \N__7839\,
            lcout => \N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_RNI51EL_1_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4400\,
            in1 => \N__4362\,
            in2 => \_gnd_net_\,
            in3 => \N__8397\,
            lcout => \un1_D_UM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIJSI41_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4326\,
            in1 => \N__5681\,
            in2 => \_gnd_net_\,
            in3 => \N__7883\,
            lcout => \N_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_BUFFERS.N_102_i_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__7258\,
            in1 => \N__4265\,
            in2 => \_gnd_net_\,
            in3 => \N__7449\,
            lcout => \N_102_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_BUFFERS.un1_DMA_EN_0_0_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__7067\,
            in1 => \N__7257\,
            in2 => \_gnd_net_\,
            in3 => \N__4266\,
            lcout => \BUFDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_BUFFERS.DMA_EN_i_0_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7256\,
            in2 => \_gnd_net_\,
            in3 => \N__4264\,
            lcout => \N_104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNIPLKT_3_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8423\,
            in1 => \N__4213\,
            in2 => \_gnd_net_\,
            in3 => \N__4179\,
            lcout => \N_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100000100"
        )
    port map (
            in0 => \N__4137\,
            in1 => \N__4131\,
            in2 => \N__4125\,
            in3 => \N__4110\,
            lcout => \U111_CYCLE_SM.TS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6384\,
            ce => 'H',
            sr => \N__6336\
        );

    \U111_CYCLE_SM.TS_OUT_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101010111"
        )
    port map (
            in0 => \N__4646\,
            in1 => \N__4109\,
            in2 => \N__7438\,
            in3 => \N__5816\,
            lcout => \TS_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TS_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_RNO_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__4973\,
            in1 => \N__5086\,
            in2 => \_gnd_net_\,
            in3 => \N__6413\,
            lcout => \U111_CYCLE_SM.N_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_RNINRNR_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__5784\,
            in1 => \N__7302\,
            in2 => \N__7088\,
            in3 => \N__7323\,
            lcout => \U111_CYCLE_SM_OFFBOARD_EN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LATCH_EN_RNO_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6627\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7137\,
            lcout => \U111_CYCLE_SM.LATCH_EN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_2_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__5384\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4566\,
            lcout => \U111_CYCLE_SM.N_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_DELAY_RNIDR7G_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5817\,
            in3 => \N__7423\,
            lcout => \U111_CYCLE_SM.un4_TS_OUT_i_0\,
            ltout => \U111_CYCLE_SM.un4_TS_OUT_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNI9UTM_0_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4665\,
            in3 => \N__6626\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVE_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_2_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010110000"
        )
    port map (
            in0 => \N__5093\,
            in1 => \N__4662\,
            in2 => \N__4656\,
            in3 => \N__4593\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6378\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_2_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__5383\,
            in1 => \_gnd_net_\,
            in2 => \N__4537\,
            in3 => \N__4565\,
            lcout => \U111_CYCLE_SM.N_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGD6K_0_2_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4567\,
            in1 => \N__5382\,
            in2 => \_gnd_net_\,
            in3 => \N__4520\,
            lcout => \U111_CYCLE_SM.N_107_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_4_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__6593\,
            in1 => \N__5462\,
            in2 => \N__5451\,
            in3 => \N__7174\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6375\,
            ce => 'H',
            sr => \N__6337\
        );

    \U111_CYCLE_SM.LATCH_EN_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111000"
        )
    port map (
            in0 => \N__5133\,
            in1 => \N__5123\,
            in2 => \N__8363\,
            in3 => \N__6458\,
            lcout => \U111_CYCLE_SM.LATCH_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6375\,
            ce => 'H',
            sr => \N__6337\
        );

    \U111_CYCLE_SM.UU_LATCHED_6_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__6595\,
            in1 => \N__5699\,
            in2 => \N__5688\,
            in3 => \N__7176\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6375\,
            ce => 'H',
            sr => \N__6337\
        );

    \U111_CYCLE_SM.UM_LATCHED_7_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__7173\,
            in1 => \N__5045\,
            in2 => \N__5013\,
            in3 => \N__6592\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6375\,
            ce => 'H',
            sr => \N__6337\
        );

    \U111_CYCLE_SM.TA_DIS_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000011111110"
        )
    port map (
            in0 => \N__5124\,
            in1 => \N__5094\,
            in2 => \N__6130\,
            in3 => \N__5058\,
            lcout => \U111_CYCLE_SM.TA_DISZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6375\,
            ce => 'H',
            sr => \N__6337\
        );

    \U111_CYCLE_SM.UM_LATCHED_3_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7172\,
            in1 => \N__6026\,
            in2 => \N__6084\,
            in3 => \N__6591\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6375\,
            ce => 'H',
            sr => \N__6337\
        );

    \U111_CYCLE_SM.UU_LATCHED_7_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__6596\,
            in1 => \N__5541\,
            in2 => \N__5507\,
            in3 => \N__7177\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6375\,
            ce => 'H',
            sr => \N__6337\
        );

    \U111_CYCLE_SM.UU_LATCHED_5_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7175\,
            in1 => \N__5576\,
            in2 => \N__5625\,
            in3 => \N__6594\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6375\,
            ce => 'H',
            sr => \N__6337\
        );

    \U111_CYCLE_SM.UM_LATCHED_RNIHDEL_7_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8337\,
            in1 => \N__5044\,
            in2 => \_gnd_net_\,
            in3 => \N__5012\,
            lcout => \un1_D_UM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_THRU_LUT4_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6390\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_CLK40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNIVRKT_6_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5703\,
            in1 => \N__5668\,
            in2 => \_gnd_net_\,
            in3 => \N__8403\,
            lcout => \N_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNITPKT_5_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8402\,
            in1 => \N__5611\,
            in2 => \_gnd_net_\,
            in3 => \N__5580\,
            lcout => \N_126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNI1UKT_7_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5540\,
            in1 => \N__5508\,
            in2 => \_gnd_net_\,
            in3 => \N__8401\,
            lcout => \N_123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNIRNKT_4_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5466\,
            in1 => \N__5440\,
            in2 => \_gnd_net_\,
            in3 => \N__8404\,
            lcout => \N_127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_RNI576J_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__5388\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6137\,
            lcout => \U111_CYCLE_SM_TEA_CPUn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIJHPK_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5298\,
            in1 => \N__5276\,
            in2 => \_gnd_net_\,
            in3 => \N__7903\,
            lcout => \un1_D_UU_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIM8O01_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5220\,
            in1 => \N__5198\,
            in2 => \_gnd_net_\,
            in3 => \N__7920\,
            lcout => \un1_D_UM_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_RNI95EL_3_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6070\,
            in1 => \N__6033\,
            in2 => \_gnd_net_\,
            in3 => \N__8422\,
            lcout => \un1_D_UM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIG2O01_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6000\,
            in1 => \N__5958\,
            in2 => \_gnd_net_\,
            in3 => \N__7919\,
            lcout => \un1_D_UM_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIALT71_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7902\,
            in1 => \N__8466\,
            in2 => \_gnd_net_\,
            in3 => \N__5919\,
            lcout => \un2_D_LL_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNI8JT71_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5877\,
            in1 => \N__7698\,
            in2 => \_gnd_net_\,
            in3 => \N__7901\,
            lcout => \un2_D_LL_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_DELAY_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5838\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.TS_DELAYZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6379\,
            ce => 'H',
            sr => \N__6334\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__7167\,
            in1 => \N__6635\,
            in2 => \N__7089\,
            in3 => \N__5802\,
            lcout => \U111_CYCLE_SM.READ_CYCLE_ACTIVEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6379\,
            ce => 'H',
            sr => \N__6334\
        );

    \U111_CYCLE_SM.UM_LATCHED_2_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__6589\,
            in1 => \N__6674\,
            in2 => \N__6712\,
            in3 => \N__7139\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6376\,
            ce => 'H',
            sr => \N__6338\
        );

    \U111_CYCLE_SM.UM_LATCHED_0_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7138\,
            in1 => \N__8555\,
            in2 => \N__8540\,
            in3 => \N__6588\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6376\,
            ce => 'H',
            sr => \N__6338\
        );

    \U111_CYCLE_SM.WRITE_CYCLE_ACTIVE_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000101110"
        )
    port map (
            in0 => \N__5783\,
            in1 => \N__6642\,
            in2 => \N__7087\,
            in3 => \N__5801\,
            lcout => \U111_CYCLE_SM.WRITE_CYCLE_ACTIVEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6376\,
            ce => 'H',
            sr => \N__6338\
        );

    \U111_CYCLE_SM.CYCLE_EN_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__7318\,
            in1 => \N__6641\,
            in2 => \_gnd_net_\,
            in3 => \N__6457\,
            lcout => \U111_CYCLE_SM.CYCLE_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6376\,
            ce => 'H',
            sr => \N__6338\
        );

    \U111_CYCLE_SM.UM_LATCHED_6_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__6590\,
            in1 => \N__8477\,
            in2 => \N__8465\,
            in3 => \N__7140\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6376\,
            ce => 'H',
            sr => \N__6338\
        );

    \U111_CYCLE_SM.UU_LATCHED_1_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__6254\,
            in1 => \N__6604\,
            in2 => \N__6306\,
            in3 => \N__7171\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6374\,
            ce => 'H',
            sr => \N__6339\
        );

    \U111_CYCLE_SM.UU_LATCHED_0_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7170\,
            in1 => \N__6215\,
            in2 => \N__6200\,
            in3 => \N__6605\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6374\,
            ce => 'H',
            sr => \N__6339\
        );

    \U111_CYCLE_SM.UM_LATCHED_5_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__7646\,
            in1 => \N__6603\,
            in2 => \N__7694\,
            in3 => \N__7169\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6374\,
            ce => 'H',
            sr => \N__6339\
        );

    \U111_CYCLE_SM.LW_TRANS_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010111001100"
        )
    port map (
            in0 => \N__6533\,
            in1 => \N__6409\,
            in2 => \N__6497\,
            in3 => \N__6462\,
            lcout => \U111_CYCLE_SM.LW_TRANSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6374\,
            ce => 'H',
            sr => \N__6339\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNILHKT_1_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8425\,
            in1 => \N__6292\,
            in2 => \_gnd_net_\,
            in3 => \N__6258\,
            lcout => \N_130\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_RNIJFKT_0_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6219\,
            in1 => \N__6182\,
            in2 => \_gnd_net_\,
            in3 => \N__8424\,
            lcout => \N_131\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_DIS_RNICJKJ_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6138\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7445\,
            lcout => \N_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_RNID9EL_5_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7670\,
            in1 => \N__7653\,
            in2 => \_gnd_net_\,
            in3 => \N__8427\,
            lcout => \un1_D_UM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_RNIB7EL_4_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7611\,
            in1 => \N__7586\,
            in2 => \_gnd_net_\,
            in3 => \N__8426\,
            lcout => \un1_D_UM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIRPPK_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7918\,
            in1 => \N__7527\,
            in2 => \_gnd_net_\,
            in3 => \N__7493\,
            lcout => \un1_D_UU_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LBENn_c_sbtinv_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7408\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \LBENn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIU8T71_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7365\,
            in1 => \N__8544\,
            in2 => \_gnd_net_\,
            in3 => \N__7917\,
            lcout => \un2_D_LL_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_EN_RNI26B3_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7319\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7301\,
            lcout => \CPUBGn_c\,
            ltout => \CPUBGn_c_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.READ_CYCLE_ACTIVE_RNI8QUM_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111010"
        )
    port map (
            in0 => \N__7168\,
            in1 => \_gnd_net_\,
            in2 => \N__7092\,
            in3 => \N__7068\,
            lcout => \N_62_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_RNI73EL_2_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8396\,
            in1 => \N__6713\,
            in2 => \_gnd_net_\,
            in3 => \N__6675\,
            lcout => \un1_D_UM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_RNI3VDL_0_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8556\,
            in1 => \N__8519\,
            in2 => \_gnd_net_\,
            in3 => \N__8364\,
            lcout => \un1_D_UM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_RNIFBEL_6_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8478\,
            in1 => \N__8452\,
            in2 => \_gnd_net_\,
            in3 => \N__8365\,
            lcout => \N_125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNICUN01_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7850\,
            in1 => \N__8279\,
            in2 => \_gnd_net_\,
            in3 => \N__8238\,
            lcout => \un1_D_UM_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8205\,
            lcout => \GB_BUFFER_CLK80_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNINLPK_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7922\,
            in1 => \N__8160\,
            in2 => \_gnd_net_\,
            in3 => \N__8132\,
            lcout => \un1_D_UU_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNIVTPK_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7923\,
            in1 => \N__8073\,
            in2 => \_gnd_net_\,
            in3 => \N__8048\,
            lcout => \un1_D_UU_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.FLIP_WORD_RNII4O01_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7976\,
            in1 => \N__7941\,
            in2 => \_gnd_net_\,
            in3 => \N__7921\,
            lcout => \un1_D_UM_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

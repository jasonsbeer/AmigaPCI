// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     May 8 2025 19:39:32

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    CMA,
    DRA,
    DA,
    A,
    DBRn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    TCIn,
    TBIn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    output [10:0] CMA;
    input [9:0] DRA;
    output [2:0] DA;
    input [20:0] A;
    input DBRn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    output TCIn;
    output TBIn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__12710;
    wire N__12709;
    wire N__12708;
    wire N__12701;
    wire N__12700;
    wire N__12699;
    wire N__12692;
    wire N__12691;
    wire N__12690;
    wire N__12683;
    wire N__12682;
    wire N__12681;
    wire N__12674;
    wire N__12673;
    wire N__12672;
    wire N__12665;
    wire N__12664;
    wire N__12663;
    wire N__12656;
    wire N__12655;
    wire N__12654;
    wire N__12647;
    wire N__12646;
    wire N__12645;
    wire N__12638;
    wire N__12637;
    wire N__12636;
    wire N__12629;
    wire N__12628;
    wire N__12627;
    wire N__12620;
    wire N__12619;
    wire N__12618;
    wire N__12611;
    wire N__12610;
    wire N__12609;
    wire N__12602;
    wire N__12601;
    wire N__12600;
    wire N__12593;
    wire N__12592;
    wire N__12591;
    wire N__12584;
    wire N__12583;
    wire N__12582;
    wire N__12575;
    wire N__12574;
    wire N__12573;
    wire N__12566;
    wire N__12565;
    wire N__12564;
    wire N__12557;
    wire N__12556;
    wire N__12555;
    wire N__12548;
    wire N__12547;
    wire N__12546;
    wire N__12539;
    wire N__12538;
    wire N__12537;
    wire N__12530;
    wire N__12529;
    wire N__12528;
    wire N__12521;
    wire N__12520;
    wire N__12519;
    wire N__12512;
    wire N__12511;
    wire N__12510;
    wire N__12503;
    wire N__12502;
    wire N__12501;
    wire N__12494;
    wire N__12493;
    wire N__12492;
    wire N__12485;
    wire N__12484;
    wire N__12483;
    wire N__12476;
    wire N__12475;
    wire N__12474;
    wire N__12467;
    wire N__12466;
    wire N__12465;
    wire N__12458;
    wire N__12457;
    wire N__12456;
    wire N__12449;
    wire N__12448;
    wire N__12447;
    wire N__12440;
    wire N__12439;
    wire N__12438;
    wire N__12431;
    wire N__12430;
    wire N__12429;
    wire N__12422;
    wire N__12421;
    wire N__12420;
    wire N__12413;
    wire N__12412;
    wire N__12411;
    wire N__12404;
    wire N__12403;
    wire N__12402;
    wire N__12395;
    wire N__12394;
    wire N__12393;
    wire N__12386;
    wire N__12385;
    wire N__12384;
    wire N__12377;
    wire N__12376;
    wire N__12375;
    wire N__12368;
    wire N__12367;
    wire N__12366;
    wire N__12359;
    wire N__12358;
    wire N__12357;
    wire N__12350;
    wire N__12349;
    wire N__12348;
    wire N__12341;
    wire N__12340;
    wire N__12339;
    wire N__12332;
    wire N__12331;
    wire N__12330;
    wire N__12323;
    wire N__12322;
    wire N__12321;
    wire N__12314;
    wire N__12313;
    wire N__12312;
    wire N__12305;
    wire N__12304;
    wire N__12303;
    wire N__12296;
    wire N__12295;
    wire N__12294;
    wire N__12287;
    wire N__12286;
    wire N__12285;
    wire N__12278;
    wire N__12277;
    wire N__12276;
    wire N__12269;
    wire N__12268;
    wire N__12267;
    wire N__12260;
    wire N__12259;
    wire N__12258;
    wire N__12251;
    wire N__12250;
    wire N__12249;
    wire N__12242;
    wire N__12241;
    wire N__12240;
    wire N__12233;
    wire N__12232;
    wire N__12231;
    wire N__12224;
    wire N__12223;
    wire N__12222;
    wire N__12215;
    wire N__12214;
    wire N__12213;
    wire N__12206;
    wire N__12205;
    wire N__12204;
    wire N__12197;
    wire N__12196;
    wire N__12195;
    wire N__12188;
    wire N__12187;
    wire N__12186;
    wire N__12179;
    wire N__12178;
    wire N__12177;
    wire N__12170;
    wire N__12169;
    wire N__12168;
    wire N__12161;
    wire N__12160;
    wire N__12159;
    wire N__12152;
    wire N__12151;
    wire N__12150;
    wire N__12143;
    wire N__12142;
    wire N__12141;
    wire N__12134;
    wire N__12133;
    wire N__12132;
    wire N__12125;
    wire N__12124;
    wire N__12123;
    wire N__12116;
    wire N__12115;
    wire N__12114;
    wire N__12107;
    wire N__12106;
    wire N__12105;
    wire N__12098;
    wire N__12097;
    wire N__12096;
    wire N__12089;
    wire N__12088;
    wire N__12087;
    wire N__12080;
    wire N__12079;
    wire N__12078;
    wire N__12071;
    wire N__12070;
    wire N__12069;
    wire N__12062;
    wire N__12061;
    wire N__12060;
    wire N__12053;
    wire N__12052;
    wire N__12051;
    wire N__12044;
    wire N__12043;
    wire N__12042;
    wire N__12035;
    wire N__12034;
    wire N__12033;
    wire N__12026;
    wire N__12025;
    wire N__12024;
    wire N__12017;
    wire N__12016;
    wire N__12015;
    wire N__12008;
    wire N__12007;
    wire N__12006;
    wire N__11999;
    wire N__11998;
    wire N__11997;
    wire N__11990;
    wire N__11989;
    wire N__11988;
    wire N__11981;
    wire N__11980;
    wire N__11979;
    wire N__11972;
    wire N__11971;
    wire N__11970;
    wire N__11963;
    wire N__11962;
    wire N__11961;
    wire N__11954;
    wire N__11953;
    wire N__11952;
    wire N__11945;
    wire N__11944;
    wire N__11943;
    wire N__11936;
    wire N__11935;
    wire N__11934;
    wire N__11927;
    wire N__11926;
    wire N__11925;
    wire N__11918;
    wire N__11917;
    wire N__11916;
    wire N__11909;
    wire N__11908;
    wire N__11907;
    wire N__11900;
    wire N__11899;
    wire N__11898;
    wire N__11891;
    wire N__11890;
    wire N__11889;
    wire N__11882;
    wire N__11881;
    wire N__11880;
    wire N__11873;
    wire N__11872;
    wire N__11871;
    wire N__11864;
    wire N__11863;
    wire N__11862;
    wire N__11845;
    wire N__11842;
    wire N__11841;
    wire N__11840;
    wire N__11837;
    wire N__11836;
    wire N__11835;
    wire N__11832;
    wire N__11831;
    wire N__11828;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11813;
    wire N__11810;
    wire N__11805;
    wire N__11800;
    wire N__11797;
    wire N__11794;
    wire N__11791;
    wire N__11788;
    wire N__11785;
    wire N__11782;
    wire N__11779;
    wire N__11774;
    wire N__11771;
    wire N__11764;
    wire N__11761;
    wire N__11758;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11739;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11703;
    wire N__11700;
    wire N__11697;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11680;
    wire N__11677;
    wire N__11676;
    wire N__11675;
    wire N__11672;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11662;
    wire N__11661;
    wire N__11660;
    wire N__11659;
    wire N__11658;
    wire N__11657;
    wire N__11656;
    wire N__11655;
    wire N__11654;
    wire N__11653;
    wire N__11650;
    wire N__11649;
    wire N__11648;
    wire N__11647;
    wire N__11646;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11630;
    wire N__11625;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11611;
    wire N__11610;
    wire N__11607;
    wire N__11606;
    wire N__11601;
    wire N__11598;
    wire N__11587;
    wire N__11584;
    wire N__11581;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11573;
    wire N__11572;
    wire N__11569;
    wire N__11568;
    wire N__11565;
    wire N__11562;
    wire N__11553;
    wire N__11550;
    wire N__11547;
    wire N__11542;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11524;
    wire N__11509;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11448;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11437;
    wire N__11436;
    wire N__11435;
    wire N__11434;
    wire N__11431;
    wire N__11430;
    wire N__11427;
    wire N__11424;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11406;
    wire N__11403;
    wire N__11400;
    wire N__11397;
    wire N__11394;
    wire N__11387;
    wire N__11382;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11368;
    wire N__11367;
    wire N__11366;
    wire N__11365;
    wire N__11364;
    wire N__11363;
    wire N__11362;
    wire N__11353;
    wire N__11350;
    wire N__11349;
    wire N__11346;
    wire N__11343;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11332;
    wire N__11329;
    wire N__11326;
    wire N__11323;
    wire N__11318;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11298;
    wire N__11295;
    wire N__11290;
    wire N__11287;
    wire N__11282;
    wire N__11279;
    wire N__11274;
    wire N__11269;
    wire N__11266;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11255;
    wire N__11254;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11238;
    wire N__11229;
    wire N__11226;
    wire N__11223;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11208;
    wire N__11207;
    wire N__11202;
    wire N__11199;
    wire N__11196;
    wire N__11193;
    wire N__11190;
    wire N__11185;
    wire N__11180;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11154;
    wire N__11149;
    wire N__11148;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11140;
    wire N__11139;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11110;
    wire N__11101;
    wire N__11100;
    wire N__11097;
    wire N__11096;
    wire N__11093;
    wire N__11088;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11073;
    wire N__11070;
    wire N__11067;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11053;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11034;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11020;
    wire N__11017;
    wire N__11014;
    wire N__11011;
    wire N__11010;
    wire N__11007;
    wire N__11006;
    wire N__11003;
    wire N__11000;
    wire N__10997;
    wire N__10996;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10962;
    wire N__10957;
    wire N__10956;
    wire N__10951;
    wire N__10950;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10924;
    wire N__10921;
    wire N__10918;
    wire N__10915;
    wire N__10912;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10904;
    wire N__10899;
    wire N__10896;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10878;
    wire N__10873;
    wire N__10870;
    wire N__10867;
    wire N__10864;
    wire N__10863;
    wire N__10862;
    wire N__10861;
    wire N__10858;
    wire N__10857;
    wire N__10854;
    wire N__10853;
    wire N__10852;
    wire N__10851;
    wire N__10850;
    wire N__10849;
    wire N__10848;
    wire N__10847;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10839;
    wire N__10838;
    wire N__10837;
    wire N__10834;
    wire N__10825;
    wire N__10822;
    wire N__10817;
    wire N__10814;
    wire N__10809;
    wire N__10804;
    wire N__10801;
    wire N__10796;
    wire N__10795;
    wire N__10792;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10774;
    wire N__10773;
    wire N__10772;
    wire N__10771;
    wire N__10768;
    wire N__10765;
    wire N__10760;
    wire N__10755;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10738;
    wire N__10733;
    wire N__10728;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10700;
    wire N__10697;
    wire N__10690;
    wire N__10689;
    wire N__10688;
    wire N__10687;
    wire N__10684;
    wire N__10681;
    wire N__10678;
    wire N__10675;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10656;
    wire N__10653;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10639;
    wire N__10636;
    wire N__10633;
    wire N__10632;
    wire N__10631;
    wire N__10630;
    wire N__10629;
    wire N__10628;
    wire N__10615;
    wire N__10612;
    wire N__10609;
    wire N__10608;
    wire N__10607;
    wire N__10606;
    wire N__10605;
    wire N__10604;
    wire N__10603;
    wire N__10602;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10598;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10566;
    wire N__10565;
    wire N__10564;
    wire N__10563;
    wire N__10562;
    wire N__10559;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10541;
    wire N__10540;
    wire N__10539;
    wire N__10536;
    wire N__10535;
    wire N__10532;
    wire N__10531;
    wire N__10530;
    wire N__10529;
    wire N__10528;
    wire N__10525;
    wire N__10524;
    wire N__10523;
    wire N__10522;
    wire N__10519;
    wire N__10518;
    wire N__10517;
    wire N__10516;
    wire N__10515;
    wire N__10514;
    wire N__10513;
    wire N__10512;
    wire N__10511;
    wire N__10510;
    wire N__10509;
    wire N__10508;
    wire N__10507;
    wire N__10506;
    wire N__10505;
    wire N__10504;
    wire N__10503;
    wire N__10502;
    wire N__10501;
    wire N__10500;
    wire N__10499;
    wire N__10498;
    wire N__10497;
    wire N__10496;
    wire N__10495;
    wire N__10494;
    wire N__10493;
    wire N__10490;
    wire N__10489;
    wire N__10488;
    wire N__10487;
    wire N__10396;
    wire N__10393;
    wire N__10390;
    wire N__10389;
    wire N__10386;
    wire N__10385;
    wire N__10384;
    wire N__10381;
    wire N__10380;
    wire N__10377;
    wire N__10374;
    wire N__10371;
    wire N__10368;
    wire N__10365;
    wire N__10362;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10348;
    wire N__10345;
    wire N__10342;
    wire N__10339;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10318;
    wire N__10315;
    wire N__10314;
    wire N__10313;
    wire N__10310;
    wire N__10305;
    wire N__10300;
    wire N__10299;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10284;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10257;
    wire N__10252;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10230;
    wire N__10227;
    wire N__10224;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10207;
    wire N__10206;
    wire N__10203;
    wire N__10202;
    wire N__10201;
    wire N__10200;
    wire N__10199;
    wire N__10198;
    wire N__10197;
    wire N__10194;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10183;
    wire N__10178;
    wire N__10175;
    wire N__10174;
    wire N__10173;
    wire N__10172;
    wire N__10171;
    wire N__10170;
    wire N__10167;
    wire N__10166;
    wire N__10165;
    wire N__10164;
    wire N__10163;
    wire N__10162;
    wire N__10161;
    wire N__10160;
    wire N__10159;
    wire N__10154;
    wire N__10153;
    wire N__10152;
    wire N__10145;
    wire N__10142;
    wire N__10141;
    wire N__10136;
    wire N__10131;
    wire N__10128;
    wire N__10121;
    wire N__10118;
    wire N__10113;
    wire N__10104;
    wire N__10103;
    wire N__10102;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10088;
    wire N__10083;
    wire N__10080;
    wire N__10071;
    wire N__10064;
    wire N__10057;
    wire N__10056;
    wire N__10055;
    wire N__10052;
    wire N__10045;
    wire N__10042;
    wire N__10037;
    wire N__10032;
    wire N__10029;
    wire N__10024;
    wire N__10019;
    wire N__10014;
    wire N__10009;
    wire N__10006;
    wire N__9999;
    wire N__9996;
    wire N__9993;
    wire N__9988;
    wire N__9985;
    wire N__9982;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9969;
    wire N__9968;
    wire N__9967;
    wire N__9966;
    wire N__9965;
    wire N__9964;
    wire N__9963;
    wire N__9962;
    wire N__9961;
    wire N__9960;
    wire N__9959;
    wire N__9958;
    wire N__9957;
    wire N__9956;
    wire N__9955;
    wire N__9954;
    wire N__9953;
    wire N__9952;
    wire N__9951;
    wire N__9950;
    wire N__9949;
    wire N__9948;
    wire N__9947;
    wire N__9946;
    wire N__9945;
    wire N__9944;
    wire N__9943;
    wire N__9942;
    wire N__9941;
    wire N__9940;
    wire N__9939;
    wire N__9938;
    wire N__9937;
    wire N__9936;
    wire N__9935;
    wire N__9934;
    wire N__9931;
    wire N__9930;
    wire N__9929;
    wire N__9928;
    wire N__9927;
    wire N__9926;
    wire N__9925;
    wire N__9924;
    wire N__9923;
    wire N__9832;
    wire N__9829;
    wire N__9828;
    wire N__9823;
    wire N__9822;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9788;
    wire N__9785;
    wire N__9780;
    wire N__9775;
    wire N__9774;
    wire N__9771;
    wire N__9768;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9742;
    wire N__9739;
    wire N__9736;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9714;
    wire N__9711;
    wire N__9708;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9697;
    wire N__9690;
    wire N__9687;
    wire N__9684;
    wire N__9681;
    wire N__9678;
    wire N__9673;
    wire N__9670;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9646;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9638;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9615;
    wire N__9610;
    wire N__9607;
    wire N__9604;
    wire N__9601;
    wire N__9598;
    wire N__9595;
    wire N__9592;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9580;
    wire N__9579;
    wire N__9576;
    wire N__9573;
    wire N__9572;
    wire N__9567;
    wire N__9566;
    wire N__9565;
    wire N__9562;
    wire N__9559;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9541;
    wire N__9538;
    wire N__9535;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9514;
    wire N__9511;
    wire N__9508;
    wire N__9505;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9490;
    wire N__9487;
    wire N__9484;
    wire N__9481;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9469;
    wire N__9466;
    wire N__9463;
    wire N__9460;
    wire N__9459;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9451;
    wire N__9448;
    wire N__9445;
    wire N__9444;
    wire N__9441;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9429;
    wire N__9424;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9412;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9333;
    wire N__9332;
    wire N__9331;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9312;
    wire N__9309;
    wire N__9306;
    wire N__9303;
    wire N__9300;
    wire N__9295;
    wire N__9292;
    wire N__9289;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9270;
    wire N__9265;
    wire N__9262;
    wire N__9259;
    wire N__9256;
    wire N__9255;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9210;
    wire N__9209;
    wire N__9208;
    wire N__9205;
    wire N__9202;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9190;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9170;
    wire N__9167;
    wire N__9164;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9147;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9094;
    wire N__9091;
    wire N__9088;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9037;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9021;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9009;
    wire N__9004;
    wire N__9001;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8986;
    wire N__8983;
    wire N__8980;
    wire N__8977;
    wire N__8974;
    wire N__8971;
    wire N__8970;
    wire N__8967;
    wire N__8966;
    wire N__8965;
    wire N__8964;
    wire N__8963;
    wire N__8962;
    wire N__8961;
    wire N__8960;
    wire N__8959;
    wire N__8958;
    wire N__8953;
    wire N__8952;
    wire N__8951;
    wire N__8950;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8942;
    wire N__8939;
    wire N__8938;
    wire N__8933;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8902;
    wire N__8897;
    wire N__8892;
    wire N__8891;
    wire N__8890;
    wire N__8889;
    wire N__8888;
    wire N__8885;
    wire N__8880;
    wire N__8875;
    wire N__8870;
    wire N__8867;
    wire N__8860;
    wire N__8859;
    wire N__8858;
    wire N__8857;
    wire N__8856;
    wire N__8853;
    wire N__8848;
    wire N__8839;
    wire N__8830;
    wire N__8821;
    wire N__8820;
    wire N__8819;
    wire N__8818;
    wire N__8817;
    wire N__8816;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8802;
    wire N__8797;
    wire N__8788;
    wire N__8785;
    wire N__8784;
    wire N__8783;
    wire N__8782;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8772;
    wire N__8771;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8761;
    wire N__8756;
    wire N__8753;
    wire N__8752;
    wire N__8751;
    wire N__8748;
    wire N__8743;
    wire N__8738;
    wire N__8737;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8704;
    wire N__8701;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8680;
    wire N__8679;
    wire N__8674;
    wire N__8673;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8640;
    wire N__8637;
    wire N__8634;
    wire N__8631;
    wire N__8626;
    wire N__8625;
    wire N__8624;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8610;
    wire N__8609;
    wire N__8606;
    wire N__8605;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8580;
    wire N__8575;
    wire N__8574;
    wire N__8573;
    wire N__8572;
    wire N__8569;
    wire N__8562;
    wire N__8557;
    wire N__8554;
    wire N__8553;
    wire N__8552;
    wire N__8551;
    wire N__8548;
    wire N__8543;
    wire N__8540;
    wire N__8535;
    wire N__8530;
    wire N__8527;
    wire N__8524;
    wire N__8523;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8500;
    wire N__8497;
    wire N__8496;
    wire N__8495;
    wire N__8494;
    wire N__8493;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8476;
    wire N__8467;
    wire N__8464;
    wire N__8463;
    wire N__8460;
    wire N__8457;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8431;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8233;
    wire N__8230;
    wire N__8227;
    wire N__8224;
    wire N__8221;
    wire N__8220;
    wire N__8217;
    wire N__8214;
    wire N__8211;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8185;
    wire N__8182;
    wire N__8179;
    wire N__8178;
    wire N__8177;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8163;
    wire N__8160;
    wire N__8159;
    wire N__8158;
    wire N__8153;
    wire N__8148;
    wire N__8143;
    wire N__8140;
    wire N__8139;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8131;
    wire N__8130;
    wire N__8127;
    wire N__8122;
    wire N__8117;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8098;
    wire N__8095;
    wire N__8092;
    wire N__8089;
    wire N__8086;
    wire N__8083;
    wire N__8080;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8037;
    wire N__8036;
    wire N__8035;
    wire N__8034;
    wire N__8031;
    wire N__8030;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8013;
    wire N__8010;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7990;
    wire N__7989;
    wire N__7986;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7969;
    wire N__7966;
    wire N__7963;
    wire N__7960;
    wire N__7959;
    wire N__7958;
    wire N__7957;
    wire N__7956;
    wire N__7955;
    wire N__7952;
    wire N__7951;
    wire N__7948;
    wire N__7945;
    wire N__7944;
    wire N__7943;
    wire N__7942;
    wire N__7941;
    wire N__7940;
    wire N__7937;
    wire N__7936;
    wire N__7935;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7918;
    wire N__7909;
    wire N__7906;
    wire N__7903;
    wire N__7896;
    wire N__7879;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7867;
    wire N__7864;
    wire N__7861;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7849;
    wire N__7846;
    wire N__7843;
    wire N__7840;
    wire N__7837;
    wire N__7834;
    wire N__7833;
    wire N__7830;
    wire N__7827;
    wire N__7824;
    wire N__7821;
    wire N__7818;
    wire N__7815;
    wire N__7810;
    wire N__7807;
    wire N__7804;
    wire N__7801;
    wire N__7798;
    wire N__7795;
    wire N__7792;
    wire N__7789;
    wire N__7786;
    wire N__7783;
    wire N__7780;
    wire N__7777;
    wire N__7774;
    wire N__7771;
    wire N__7768;
    wire N__7765;
    wire N__7762;
    wire N__7759;
    wire N__7758;
    wire N__7753;
    wire N__7750;
    wire N__7749;
    wire N__7746;
    wire N__7743;
    wire N__7742;
    wire N__7739;
    wire N__7736;
    wire N__7733;
    wire N__7730;
    wire N__7727;
    wire N__7724;
    wire N__7721;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7696;
    wire N__7689;
    wire N__7686;
    wire N__7681;
    wire N__7680;
    wire N__7677;
    wire N__7674;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7654;
    wire N__7651;
    wire N__7648;
    wire N__7645;
    wire N__7642;
    wire N__7641;
    wire N__7640;
    wire N__7637;
    wire N__7636;
    wire N__7633;
    wire N__7632;
    wire N__7629;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7596;
    wire N__7595;
    wire N__7594;
    wire N__7591;
    wire N__7588;
    wire N__7583;
    wire N__7576;
    wire N__7573;
    wire N__7570;
    wire N__7569;
    wire N__7568;
    wire N__7567;
    wire N__7566;
    wire N__7563;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7543;
    wire N__7542;
    wire N__7539;
    wire N__7538;
    wire N__7537;
    wire N__7536;
    wire N__7535;
    wire N__7534;
    wire N__7533;
    wire N__7528;
    wire N__7527;
    wire N__7526;
    wire N__7523;
    wire N__7522;
    wire N__7519;
    wire N__7516;
    wire N__7513;
    wire N__7510;
    wire N__7507;
    wire N__7506;
    wire N__7503;
    wire N__7498;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7477;
    wire N__7462;
    wire N__7459;
    wire N__7456;
    wire N__7455;
    wire N__7452;
    wire N__7449;
    wire N__7446;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7434;
    wire N__7431;
    wire N__7428;
    wire N__7423;
    wire N__7422;
    wire N__7419;
    wire N__7416;
    wire N__7411;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7399;
    wire N__7396;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7386;
    wire N__7385;
    wire N__7384;
    wire N__7381;
    wire N__7376;
    wire N__7373;
    wire N__7366;
    wire N__7363;
    wire N__7360;
    wire N__7357;
    wire N__7356;
    wire N__7353;
    wire N__7350;
    wire N__7345;
    wire N__7344;
    wire N__7341;
    wire N__7340;
    wire N__7337;
    wire N__7336;
    wire N__7335;
    wire N__7332;
    wire N__7329;
    wire N__7326;
    wire N__7325;
    wire N__7322;
    wire N__7319;
    wire N__7316;
    wire N__7313;
    wire N__7310;
    wire N__7309;
    wire N__7308;
    wire N__7307;
    wire N__7306;
    wire N__7305;
    wire N__7304;
    wire N__7303;
    wire N__7302;
    wire N__7299;
    wire N__7294;
    wire N__7291;
    wire N__7286;
    wire N__7281;
    wire N__7278;
    wire N__7273;
    wire N__7266;
    wire N__7249;
    wire N__7246;
    wire N__7245;
    wire N__7244;
    wire N__7243;
    wire N__7240;
    wire N__7237;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7222;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7206;
    wire N__7195;
    wire N__7194;
    wire N__7191;
    wire N__7190;
    wire N__7189;
    wire N__7188;
    wire N__7187;
    wire N__7186;
    wire N__7185;
    wire N__7182;
    wire N__7179;
    wire N__7176;
    wire N__7173;
    wire N__7172;
    wire N__7171;
    wire N__7170;
    wire N__7169;
    wire N__7168;
    wire N__7167;
    wire N__7166;
    wire N__7163;
    wire N__7162;
    wire N__7161;
    wire N__7160;
    wire N__7159;
    wire N__7156;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7129;
    wire N__7128;
    wire N__7127;
    wire N__7126;
    wire N__7125;
    wire N__7124;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7110;
    wire N__7107;
    wire N__7102;
    wire N__7099;
    wire N__7096;
    wire N__7091;
    wire N__7082;
    wire N__7075;
    wire N__7062;
    wire N__7051;
    wire N__7048;
    wire N__7033;
    wire N__7032;
    wire N__7031;
    wire N__7030;
    wire N__7027;
    wire N__7026;
    wire N__7025;
    wire N__7024;
    wire N__7023;
    wire N__7022;
    wire N__7021;
    wire N__7020;
    wire N__7019;
    wire N__7018;
    wire N__7017;
    wire N__7016;
    wire N__7013;
    wire N__7008;
    wire N__7005;
    wire N__7004;
    wire N__7003;
    wire N__7002;
    wire N__7001;
    wire N__7000;
    wire N__6999;
    wire N__6990;
    wire N__6987;
    wire N__6986;
    wire N__6985;
    wire N__6984;
    wire N__6983;
    wire N__6982;
    wire N__6979;
    wire N__6978;
    wire N__6977;
    wire N__6972;
    wire N__6969;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6955;
    wire N__6948;
    wire N__6945;
    wire N__6940;
    wire N__6937;
    wire N__6926;
    wire N__6917;
    wire N__6892;
    wire N__6891;
    wire N__6890;
    wire N__6887;
    wire N__6886;
    wire N__6885;
    wire N__6882;
    wire N__6877;
    wire N__6874;
    wire N__6873;
    wire N__6870;
    wire N__6867;
    wire N__6866;
    wire N__6865;
    wire N__6864;
    wire N__6863;
    wire N__6860;
    wire N__6859;
    wire N__6858;
    wire N__6857;
    wire N__6856;
    wire N__6855;
    wire N__6852;
    wire N__6849;
    wire N__6846;
    wire N__6843;
    wire N__6840;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6822;
    wire N__6819;
    wire N__6816;
    wire N__6793;
    wire N__6792;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6784;
    wire N__6779;
    wire N__6778;
    wire N__6777;
    wire N__6774;
    wire N__6773;
    wire N__6772;
    wire N__6771;
    wire N__6768;
    wire N__6765;
    wire N__6764;
    wire N__6761;
    wire N__6760;
    wire N__6759;
    wire N__6758;
    wire N__6755;
    wire N__6754;
    wire N__6753;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6741;
    wire N__6736;
    wire N__6731;
    wire N__6726;
    wire N__6723;
    wire N__6720;
    wire N__6715;
    wire N__6712;
    wire N__6691;
    wire N__6688;
    wire N__6685;
    wire N__6682;
    wire N__6679;
    wire N__6676;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6664;
    wire N__6661;
    wire N__6658;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6646;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6616;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6603;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6501;
    wire N__6498;
    wire N__6495;
    wire N__6492;
    wire N__6487;
    wire N__6484;
    wire N__6481;
    wire N__6478;
    wire N__6475;
    wire N__6472;
    wire N__6469;
    wire N__6466;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6408;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6373;
    wire N__6370;
    wire N__6369;
    wire N__6366;
    wire N__6363;
    wire N__6360;
    wire N__6355;
    wire N__6352;
    wire N__6349;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6283;
    wire N__6280;
    wire N__6277;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6267;
    wire N__6264;
    wire N__6259;
    wire N__6256;
    wire N__6255;
    wire N__6252;
    wire N__6249;
    wire N__6244;
    wire N__6243;
    wire N__6240;
    wire N__6237;
    wire N__6232;
    wire N__6231;
    wire N__6230;
    wire N__6227;
    wire N__6224;
    wire N__6221;
    wire N__6218;
    wire N__6211;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6199;
    wire N__6196;
    wire N__6193;
    wire N__6190;
    wire N__6187;
    wire N__6186;
    wire N__6183;
    wire N__6180;
    wire N__6177;
    wire N__6172;
    wire N__6169;
    wire N__6168;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6141;
    wire N__6140;
    wire N__6137;
    wire N__6132;
    wire N__6127;
    wire N__6124;
    wire N__6123;
    wire N__6120;
    wire N__6117;
    wire N__6114;
    wire N__6113;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6082;
    wire N__6075;
    wire N__6072;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6042;
    wire N__6039;
    wire N__6036;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5995;
    wire N__5992;
    wire N__5989;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5961;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5944;
    wire N__5941;
    wire N__5940;
    wire N__5939;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5907;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5889;
    wire N__5886;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5874;
    wire N__5871;
    wire N__5868;
    wire N__5865;
    wire N__5862;
    wire N__5859;
    wire N__5854;
    wire N__5853;
    wire N__5848;
    wire N__5845;
    wire N__5842;
    wire N__5839;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5809;
    wire N__5806;
    wire N__5803;
    wire N__5802;
    wire N__5801;
    wire N__5800;
    wire N__5797;
    wire N__5792;
    wire N__5789;
    wire N__5782;
    wire N__5781;
    wire N__5776;
    wire N__5773;
    wire N__5772;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5733;
    wire N__5732;
    wire N__5731;
    wire N__5728;
    wire N__5727;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5707;
    wire N__5706;
    wire N__5703;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5691;
    wire N__5688;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5652;
    wire N__5651;
    wire N__5648;
    wire N__5645;
    wire N__5642;
    wire N__5635;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5596;
    wire N__5595;
    wire N__5590;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5577;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5551;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5532;
    wire N__5529;
    wire N__5526;
    wire N__5523;
    wire N__5518;
    wire N__5515;
    wire N__5514;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5475;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5463;
    wire N__5460;
    wire N__5457;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5434;
    wire N__5431;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5423;
    wire N__5422;
    wire N__5421;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5407;
    wire N__5404;
    wire N__5395;
    wire N__5394;
    wire N__5393;
    wire N__5386;
    wire N__5385;
    wire N__5384;
    wire N__5383;
    wire N__5382;
    wire N__5379;
    wire N__5376;
    wire N__5369;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5331;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5319;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5218;
    wire N__5215;
    wire N__5214;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5188;
    wire N__5187;
    wire N__5184;
    wire N__5183;
    wire N__5182;
    wire N__5179;
    wire N__5172;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5146;
    wire N__5143;
    wire N__5140;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5101;
    wire N__5100;
    wire N__5097;
    wire N__5094;
    wire N__5089;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5040;
    wire N__5039;
    wire N__5034;
    wire N__5033;
    wire N__5032;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5020;
    wire N__5011;
    wire N__5008;
    wire N__5007;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4984;
    wire N__4981;
    wire N__4978;
    wire N__4975;
    wire N__4974;
    wire N__4973;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4954;
    wire N__4951;
    wire N__4942;
    wire N__4939;
    wire N__4936;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4912;
    wire N__4909;
    wire N__4906;
    wire N__4903;
    wire N__4900;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4892;
    wire N__4887;
    wire N__4884;
    wire N__4879;
    wire N__4876;
    wire N__4873;
    wire N__4872;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4855;
    wire N__4854;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4837;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4816;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4804;
    wire N__4801;
    wire N__4798;
    wire N__4797;
    wire N__4796;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4777;
    wire N__4774;
    wire N__4771;
    wire N__4768;
    wire N__4765;
    wire N__4762;
    wire N__4761;
    wire N__4756;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4734;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4695;
    wire N__4692;
    wire N__4689;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4645;
    wire N__4642;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4603;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4591;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4579;
    wire N__4578;
    wire N__4575;
    wire N__4572;
    wire N__4567;
    wire N__4564;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4552;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4540;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4525;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4459;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4429;
    wire N__4426;
    wire N__4423;
    wire N__4420;
    wire N__4417;
    wire N__4414;
    wire N__4411;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4384;
    wire N__4381;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4371;
    wire N__4370;
    wire N__4369;
    wire N__4368;
    wire N__4367;
    wire N__4366;
    wire N__4365;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4324;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4309;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire DBRn_c_i_0;
    wire CLK80_PLL_i_i;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_6_6_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire A_c_2;
    wire A_c_4;
    wire A_c_7;
    wire A_c_8;
    wire REGSPACEn_c;
    wire \U712_CHIP_RAM.m93_i_a2_4_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH5lto7_0_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH5lt7 ;
    wire \U712_CHIP_RAM.N_430_cascade_ ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_4 ;
    wire \U712_CHIP_RAM.N_428 ;
    wire \U712_CHIP_RAM.N_307_cascade_ ;
    wire \U712_CHIP_RAM.N_467_cascade_ ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_3 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0 ;
    wire DBRn_c;
    wire TSn_c;
    wire RAMSPACEn_c;
    wire \U712_CHIP_RAM.N_419 ;
    wire VBENn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDs_0_4 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_ ;
    wire \U712_CHIP_RAM.N_396_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_0_2 ;
    wire \U712_CHIP_RAM.N_397 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_1_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMDs_0_1 ;
    wire \U712_CHIP_RAM.N_194_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_1 ;
    wire \U712_CHIP_RAM.N_305_cascade_ ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ;
    wire \U712_CHIP_RAM.N_325 ;
    wire \U712_CHIP_RAM.N_325_cascade_ ;
    wire \U712_CHIP_RAM.m101_i_0_cascade_ ;
    wire \U712_CHIP_RAM.m101_i_1 ;
    wire \U712_CHIP_RAM.N_376 ;
    wire \U712_CHIP_RAM.m101_i_2_cascade_ ;
    wire \U712_CHIP_RAM.N_436 ;
    wire bfn_8_8_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.N_378 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.N_551_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a3_0_a2_0 ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0 ;
    wire DBDIR_c;
    wire \U712_REG_SM.N_412 ;
    wire \U712_REG_SM.N_402 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_0 ;
    wire REGENn_c;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.REGENn_e_1 ;
    wire A_c_16;
    wire A_c_17;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ;
    wire A_c_18;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.N_555 ;
    wire \U712_CHIP_RAM.N_555_cascade_ ;
    wire \U712_CHIP_RAM.N_194 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_2_2_cascade_ ;
    wire \U712_CHIP_RAM.N_449 ;
    wire \U712_CHIP_RAM.N_476 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.N_304_cascade_ ;
    wire \U712_CHIP_RAM.N_312_cascade_ ;
    wire \U712_CHIP_RAM.N_326_cascade_ ;
    wire \U712_CHIP_RAM.N_467 ;
    wire \U712_CHIP_RAM.N_39 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire \U712_CHIP_RAM.N_440 ;
    wire \U712_CHIP_RAM.N_39_cascade_ ;
    wire \U712_CHIP_RAM.N_326 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.DBENn_7_0_0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_344_cascade_ ;
    wire \U712_CHIP_RAM.N_551 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER41_2_0_cascade_ ;
    wire \U712_CHIP_RAM.LATCH_CLK_6 ;
    wire LATCH_CLK_c;
    wire AWEn_c;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ;
    wire A_c_20;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ;
    wire \U712_CHIP_RAM.N_435 ;
    wire DBR_SYNCZ0Z_0;
    wire \U712_REG_SM.N_413_cascade_ ;
    wire DBENn_c;
    wire DMA_CYCLEm;
    wire \U712_REG_SM.N_308 ;
    wire \U712_REG_SM.N_308_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_STATEZ1Z_2 ;
    wire \U712_REG_SM.N_410_cascade_ ;
    wire \U712_REG_SM.N_331 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire TACK_OUTn;
    wire \U712_REG_SM.N_404 ;
    wire LDSn_c;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.N_459 ;
    wire UDSn_c;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_0 ;
    wire bfn_10_5_0_;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_1 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_2 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_4 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_3 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_5 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_4 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_6 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_5 ;
    wire \U712_CHIP_RAM.un3_DBR_COUNT_cry_6 ;
    wire A_c_12;
    wire A_c_10;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_3 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_2 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_1 ;
    wire \U712_CHIP_RAM.DBR_COUNTZ0Z_7 ;
    wire \U712_CHIP_RAM.m93_i_a2_5 ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.N_304 ;
    wire \U712_CHIP_RAM.N_305 ;
    wire \U712_CHIP_RAM.m123_i_2_cascade_ ;
    wire A_c_15;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_2_0 ;
    wire \U712_CHIP_RAM.N_390 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_2_3 ;
    wire A_c_11;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ;
    wire A_c_3;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ;
    wire A_c_5;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ;
    wire A_c_6;
    wire \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ;
    wire REG_CYCLEm;
    wire N_167_i;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_321 ;
    wire \U712_CHIP_RAM.N_321_cascade_ ;
    wire \U712_CHIP_RAM.N_20_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.m77_0_a2_0_2_cascade_ ;
    wire \U712_CHIP_RAM.N_307 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDsr_6 ;
    wire \U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire N_202_i;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire TACK_EN;
    wire \U712_REG_SM.N_328 ;
    wire \U712_REG_SM.N_406 ;
    wire DBR_SYNCZ0Z_1;
    wire \U712_REG_SM.N_330_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_2 ;
    wire \U712_REG_SM.STATE_COUNTc_0_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_373 ;
    wire \U712_REG_SM.WRITE_CYCLEZ0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_373_cascade_ ;
    wire \U712_REG_SM.N_130 ;
    wire \U712_REG_SM.un1_REGENn_0_sqmuxa_0 ;
    wire \U712_CHIP_RAM.N_335 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire ASn_c;
    wire \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0 ;
    wire N_165_i;
    wire CONSTANT_ONE_NET;
    wire RASn_c;
    wire WEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire \U712_CHIP_RAM.N_314_cascade_ ;
    wire A_c_14;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ;
    wire \U712_CHIP_RAM.un1_CMA25_0_i ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ;
    wire \U712_CHIP_RAM.N_190 ;
    wire A_c_13;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ;
    wire \U712_CYCLE_TERM.N_332 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire \U712_CYCLE_TERM.N_455_cascade_ ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire REG_TACK;
    wire CPU_TACKm;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_1 ;
    wire \U712_REG_SM.START_RSTZ0 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.N_361 ;
    wire \U712_CHIP_RAM.N_367 ;
    wire CMA_c_5;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ;
    wire CMA_c_8;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire A_c_9;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_ ;
    wire \U712_CHIP_RAM.N_314 ;
    wire CMA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.m50_i_a2_0_0 ;
    wire N_200_i;
    wire \U712_CHIP_RAM.N_337 ;
    wire CLK40_PLL_i;
    wire CLK40_PLL_i_i;
    wire RESETn_c_i;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire \U712_CHIP_RAM.CMA_5_i_0_9 ;
    wire A_c_19;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.un1_CMA25_0_i_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire RAS1n_c;
    wire RAS0n_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire RESETn_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_2 ;
    wire CLK80_PLL;
    wire DRA_c_1;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire N_334_cascade_;
    wire N_177_i;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ;
    wire N_336_cascade_;
    wire CPU_CYCLEm;
    wire N_175_i;
    wire N_337_i;
    wire N_336_i;
    wire N_335_i;
    wire A_c_1;
    wire A_c_0;
    wire SIZ_c_1;
    wire SIZ_c_0;
    wire N_334_i;
    wire DRA_c_4;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire DRA_c_6;
    wire AGNUS_REV_c;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire RnW_c;
    wire CASLn_c;
    wire CASUn_c;
    wire DMA_WRITE_CYCLE;
    wire N_379;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__4330),
            .RESETB(N__7834),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__12710),
            .DIN(N__12709),
            .DOUT(N__12708),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__12710),
            .PADOUT(N__12709),
            .PADIN(N__12708),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5815),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__12701),
            .DIN(N__12700),
            .DOUT(N__12699),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__12701),
            .PADOUT(N__12700),
            .PADIN(N__12699),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__12692),
            .DIN(N__12691),
            .DOUT(N__12690),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__12692),
            .PADOUT(N__12691),
            .PADIN(N__12690),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8452),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__12683),
            .DIN(N__12682),
            .DOUT(N__12681),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__12683),
            .PADOUT(N__12682),
            .PADIN(N__12681),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11722),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__12674),
            .DIN(N__12673),
            .DOUT(N__12672),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__12674),
            .PADOUT(N__12673),
            .PADIN(N__12672),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__12665),
            .DIN(N__12664),
            .DOUT(N__12663),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__12665),
            .PADOUT(N__12664),
            .PADIN(N__12663),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__12656),
            .DIN(N__12655),
            .DOUT(N__12654),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__12656),
            .PADOUT(N__12655),
            .PADIN(N__12654),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__12647),
            .DIN(N__12646),
            .DOUT(N__12645),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__12647),
            .PADOUT(N__12646),
            .PADIN(N__12645),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__12638),
            .DIN(N__12637),
            .DOUT(N__12636),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__12638),
            .PADOUT(N__12637),
            .PADIN(N__12636),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__12629),
            .DIN(N__12628),
            .DOUT(N__12627),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__12629),
            .PADOUT(N__12628),
            .PADIN(N__12627),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__12620),
            .DIN(N__12619),
            .DOUT(N__12618),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__12620),
            .PADOUT(N__12619),
            .PADIN(N__12618),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__12611),
            .DIN(N__12610),
            .DOUT(N__12609),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__12611),
            .PADOUT(N__12610),
            .PADIN(N__12609),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9046),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__12602),
            .DIN(N__12601),
            .DOUT(N__12600),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__12602),
            .PADOUT(N__12601),
            .PADIN(N__12600),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11473),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__12593),
            .DIN(N__12592),
            .DOUT(N__12591),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__12593),
            .PADOUT(N__12592),
            .PADIN(N__12591),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__12584),
            .DIN(N__12583),
            .DOUT(N__12582),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__12584),
            .PADOUT(N__12583),
            .PADIN(N__12582),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__12575),
            .DIN(N__12574),
            .DOUT(N__12573),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__12575),
            .PADOUT(N__12574),
            .PADIN(N__12573),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__12566),
            .DIN(N__12565),
            .DOUT(N__12564),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__12566),
            .PADOUT(N__12565),
            .PADIN(N__12564),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4627),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__12557),
            .DIN(N__12556),
            .DOUT(N__12555),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__12557),
            .PADOUT(N__12556),
            .PADIN(N__12555),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__12548),
            .DIN(N__12547),
            .DOUT(N__12546),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__12548),
            .PADOUT(N__12547),
            .PADIN(N__12546),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__12539),
            .DIN(N__12538),
            .DOUT(N__12537),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__12539),
            .PADOUT(N__12538),
            .PADIN(N__12537),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9070),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__12530),
            .DIN(N__12529),
            .DOUT(N__12528),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__12530),
            .PADOUT(N__12529),
            .PADIN(N__12528),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__12521),
            .DIN(N__12520),
            .DOUT(N__12519),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__12521),
            .PADOUT(N__12520),
            .PADIN(N__12519),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9541),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__12512),
            .DIN(N__12511),
            .DOUT(N__12510),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__12512),
            .PADOUT(N__12511),
            .PADIN(N__12510),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__12503),
            .DIN(N__12502),
            .DOUT(N__12501),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__12503),
            .PADOUT(N__12502),
            .PADIN(N__12501),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11461),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__12494),
            .DIN(N__12493),
            .DOUT(N__12492),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__12494),
            .PADOUT(N__12493),
            .PADIN(N__12492),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7749),
            .DIN0(),
            .DOUT0(N__6113),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__12485),
            .DIN(N__12484),
            .DOUT(N__12483),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__12485),
            .PADOUT(N__12484),
            .PADIN(N__12483),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__12476),
            .DIN(N__12475),
            .DOUT(N__12474),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__12476),
            .PADOUT(N__12475),
            .PADIN(N__12474),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__12467),
            .DIN(N__12466),
            .DOUT(N__12465),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__12467),
            .PADOUT(N__12466),
            .PADIN(N__12465),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__12458),
            .DIN(N__12457),
            .DOUT(N__12456),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__12458),
            .PADOUT(N__12457),
            .PADIN(N__12456),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__12449),
            .DIN(N__12448),
            .DOUT(N__12447),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__12449),
            .PADOUT(N__12448),
            .PADIN(N__12447),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__12440),
            .DIN(N__12439),
            .DOUT(N__12438),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__12440),
            .PADOUT(N__12439),
            .PADIN(N__12438),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7852),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__12431),
            .DIN(N__12430),
            .DOUT(N__12429),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__12431),
            .PADOUT(N__12430),
            .PADIN(N__12429),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__12422),
            .DIN(N__12421),
            .DOUT(N__12420),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__12422),
            .PADOUT(N__12421),
            .PADIN(N__12420),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__12413),
            .DIN(N__12412),
            .DOUT(N__12411),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__12413),
            .PADOUT(N__12412),
            .PADIN(N__12411),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__12404),
            .DIN(N__12403),
            .DOUT(N__12402),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__12404),
            .PADOUT(N__12403),
            .PADIN(N__12402),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__12395),
            .DIN(N__12394),
            .DOUT(N__12393),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__12395),
            .PADOUT(N__12394),
            .PADIN(N__12393),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__12386),
            .DIN(N__12385),
            .DOUT(N__12384),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__12386),
            .PADOUT(N__12385),
            .PADIN(N__12384),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7810),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__12377),
            .DIN(N__12376),
            .DOUT(N__12375),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__12377),
            .PADOUT(N__12376),
            .PADIN(N__12375),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__12368),
            .DIN(N__12367),
            .DOUT(N__12366),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__12368),
            .PADOUT(N__12367),
            .PADIN(N__12366),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__12359),
            .DIN(N__12358),
            .DOUT(N__12357),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__12359),
            .PADOUT(N__12358),
            .PADIN(N__12357),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7879),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_0_iopad (
            .OE(N__12350),
            .DIN(N__12349),
            .DOUT(N__12348),
            .PACKAGEPIN(DA[0]));
    defparam DA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_0_preio (
            .PADOEN(N__12350),
            .PADOUT(N__12349),
            .PADIN(N__12348),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9025),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__12341),
            .DIN(N__12340),
            .DOUT(N__12339),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__12341),
            .PADOUT(N__12340),
            .PADIN(N__12339),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__12332),
            .DIN(N__12331),
            .DOUT(N__12330),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__12332),
            .PADOUT(N__12331),
            .PADIN(N__12330),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8404),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__12323),
            .DIN(N__12322),
            .DOUT(N__12321),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__12323),
            .PADOUT(N__12322),
            .PADIN(N__12321),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8329),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__12314),
            .DIN(N__12313),
            .DOUT(N__12312),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__12314),
            .PADOUT(N__12313),
            .PADIN(N__12312),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5227),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__12305),
            .DIN(N__12304),
            .DOUT(N__12303),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__12305),
            .PADOUT(N__12304),
            .PADIN(N__12303),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__12296),
            .DIN(N__12295),
            .DOUT(N__12294),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__12296),
            .PADOUT(N__12295),
            .PADIN(N__12294),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__12287),
            .DIN(N__12286),
            .DOUT(N__12285),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__12287),
            .PADOUT(N__12286),
            .PADIN(N__12285),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9238),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__12278),
            .DIN(N__12277),
            .DOUT(N__12276),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__12278),
            .PADOUT(N__12277),
            .PADIN(N__12276),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7750),
            .DIN0(),
            .DOUT0(N__6127),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__12269),
            .DIN(N__12268),
            .DOUT(N__12267),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__12269),
            .PADOUT(N__12268),
            .PADIN(N__12267),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7789),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__12260),
            .DIN(N__12259),
            .DOUT(N__12258),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__12260),
            .PADOUT(N__12259),
            .PADIN(N__12258),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5077),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__12251),
            .DIN(N__12250),
            .DOUT(N__12249),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__12251),
            .PADOUT(N__12250),
            .PADIN(N__12249),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9736),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__12242),
            .DIN(N__12241),
            .DOUT(N__12240),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__12242),
            .PADOUT(N__12241),
            .PADIN(N__12240),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__12233),
            .DIN(N__12232),
            .DOUT(N__12231),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__12233),
            .PADOUT(N__12232),
            .PADIN(N__12231),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_2_iopad (
            .OE(N__12224),
            .DIN(N__12223),
            .DOUT(N__12222),
            .PACKAGEPIN(DA[2]));
    defparam DA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_2_preio (
            .PADOEN(N__12224),
            .PADOUT(N__12223),
            .PADIN(N__12222),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6532),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__12215),
            .DIN(N__12214),
            .DOUT(N__12213),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__12215),
            .PADOUT(N__12214),
            .PADIN(N__12213),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__12206),
            .DIN(N__12205),
            .DOUT(N__12204),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__12206),
            .PADOUT(N__12205),
            .PADIN(N__12204),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__12197),
            .DIN(N__12196),
            .DOUT(N__12195),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__12197),
            .PADOUT(N__12196),
            .PADIN(N__12195),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8365),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__12188),
            .DIN(N__12187),
            .DOUT(N__12186),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__12188),
            .PADOUT(N__12187),
            .PADIN(N__12186),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11488),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__12179),
            .DIN(N__12178),
            .DOUT(N__12177),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__12179),
            .PADOUT(N__12178),
            .PADIN(N__12177),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__12170),
            .DIN(N__12169),
            .DOUT(N__12168),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__12170),
            .PADOUT(N__12169),
            .PADIN(N__12168),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11509),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__12161),
            .DIN(N__12160),
            .DOUT(N__12159),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__12161),
            .PADOUT(N__12160),
            .PADIN(N__12159),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7742),
            .DIN0(),
            .DOUT0(N__6123),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__12152),
            .DIN(N__12151),
            .DOUT(N__12150),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__12152),
            .PADOUT(N__12151),
            .PADIN(N__12150),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8704),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__12143),
            .DIN(N__12142),
            .DOUT(N__12141),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__12143),
            .PADOUT(N__12142),
            .PADIN(N__12141),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__12134),
            .DIN(N__12133),
            .DOUT(N__12132),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__12134),
            .PADOUT(N__12133),
            .PADIN(N__12132),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__12125),
            .DIN(N__12124),
            .DOUT(N__12123),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__12125),
            .PADOUT(N__12124),
            .PADIN(N__12123),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9094),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__12116),
            .DIN(N__12115),
            .DOUT(N__12114),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__12116),
            .PADOUT(N__12115),
            .PADIN(N__12114),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__12107),
            .DIN(N__12106),
            .DOUT(N__12105),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__12107),
            .PADOUT(N__12106),
            .PADIN(N__12105),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_1_iopad (
            .OE(N__12098),
            .DIN(N__12097),
            .DOUT(N__12096),
            .PACKAGEPIN(DA[1]));
    defparam DA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_1_preio (
            .PADOEN(N__12098),
            .PADOUT(N__12097),
            .PADIN(N__12096),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6292),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__12089),
            .DIN(N__12088),
            .DOUT(N__12087),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__12089),
            .PADOUT(N__12088),
            .PADIN(N__12087),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__12080),
            .DIN(N__12079),
            .DOUT(N__12078),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__12080),
            .PADOUT(N__12079),
            .PADIN(N__12078),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__12071),
            .DIN(N__12070),
            .DOUT(N__12069),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__12071),
            .PADOUT(N__12070),
            .PADIN(N__12069),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8425),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__12062),
            .DIN(N__12061),
            .DOUT(N__12060),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__12062),
            .PADOUT(N__12061),
            .PADIN(N__12060),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5977),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__12053),
            .DIN(N__12052),
            .DOUT(N__12051),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__12053),
            .PADOUT(N__12052),
            .PADIN(N__12051),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11029),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__12044),
            .DIN(N__12043),
            .DOUT(N__12042),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__12044),
            .PADOUT(N__12043),
            .PADIN(N__12042),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5116),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__12035),
            .DIN(N__12034),
            .DOUT(N__12033),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__12035),
            .PADOUT(N__12034),
            .PADIN(N__12033),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__12026),
            .DIN(N__12025),
            .DOUT(N__12024),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__12026),
            .PADOUT(N__12025),
            .PADIN(N__12024),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__12017),
            .DIN(N__12016),
            .DOUT(N__12015),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__12017),
            .PADOUT(N__12016),
            .PADIN(N__12015),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8302),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__12008),
            .DIN(N__12007),
            .DOUT(N__12006),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__12008),
            .PADOUT(N__12007),
            .PADIN(N__12006),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__11999),
            .DIN(N__11998),
            .DOUT(N__11997),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__11999),
            .PADOUT(N__11998),
            .PADIN(N__11997),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__11990),
            .DIN(N__11989),
            .DOUT(N__11988),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__11990),
            .PADOUT(N__11989),
            .PADIN(N__11988),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5626),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__11981),
            .DIN(N__11980),
            .DOUT(N__11979),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__11981),
            .PADOUT(N__11980),
            .PADIN(N__11979),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6058),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11972),
            .DIN(N__11971),
            .DOUT(N__11970),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11972),
            .PADOUT(N__11971),
            .PADIN(N__11970),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9151),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11963),
            .DIN(N__11962),
            .DOUT(N__11961),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11963),
            .PADOUT(N__11962),
            .PADIN(N__11961),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11954),
            .DIN(N__11953),
            .DOUT(N__11952),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11954),
            .PADOUT(N__11953),
            .PADIN(N__11952),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9147),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11945),
            .DIN(N__11944),
            .DOUT(N__11943),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11945),
            .PADOUT(N__11944),
            .PADIN(N__11943),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4420),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11936),
            .DIN(N__11935),
            .DOUT(N__11934),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11936),
            .PADOUT(N__11935),
            .PADIN(N__11934),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8353),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11927),
            .DIN(N__11926),
            .DOUT(N__11925),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11927),
            .PADOUT(N__11926),
            .PADIN(N__11925),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11918),
            .DIN(N__11917),
            .DOUT(N__11916),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11918),
            .PADOUT(N__11917),
            .PADIN(N__11916),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11909),
            .DIN(N__11908),
            .DOUT(N__11907),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11909),
            .PADOUT(N__11908),
            .PADIN(N__11907),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11900),
            .DIN(N__11899),
            .DOUT(N__11898),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11900),
            .PADOUT(N__11899),
            .PADIN(N__11898),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11891),
            .DIN(N__11890),
            .DOUT(N__11889),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11891),
            .PADOUT(N__11890),
            .PADIN(N__11889),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9146),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11882),
            .DIN(N__11881),
            .DOUT(N__11880),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11882),
            .PADOUT(N__11881),
            .PADIN(N__11880),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7411),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11873),
            .DIN(N__11872),
            .DOUT(N__11871),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11873),
            .PADOUT(N__11872),
            .PADIN(N__11871),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6634),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11864),
            .DIN(N__11863),
            .DOUT(N__11862),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11864),
            .PADOUT(N__11863),
            .PADIN(N__11862),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9481),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2884 (
            .O(N__11845),
            .I(N__11842));
    LocalMux I__2883 (
            .O(N__11842),
            .I(N__11837));
    CascadeMux I__2882 (
            .O(N__11841),
            .I(N__11832));
    CascadeMux I__2881 (
            .O(N__11840),
            .I(N__11828));
    Span4Mux_h I__2880 (
            .O(N__11837),
            .I(N__11825));
    InMux I__2879 (
            .O(N__11836),
            .I(N__11822));
    InMux I__2878 (
            .O(N__11835),
            .I(N__11819));
    InMux I__2877 (
            .O(N__11832),
            .I(N__11816));
    InMux I__2876 (
            .O(N__11831),
            .I(N__11813));
    InMux I__2875 (
            .O(N__11828),
            .I(N__11810));
    Sp12to4 I__2874 (
            .O(N__11825),
            .I(N__11805));
    LocalMux I__2873 (
            .O(N__11822),
            .I(N__11805));
    LocalMux I__2872 (
            .O(N__11819),
            .I(N__11800));
    LocalMux I__2871 (
            .O(N__11816),
            .I(N__11800));
    LocalMux I__2870 (
            .O(N__11813),
            .I(N__11797));
    LocalMux I__2869 (
            .O(N__11810),
            .I(N__11794));
    Span12Mux_v I__2868 (
            .O(N__11805),
            .I(N__11791));
    Span12Mux_h I__2867 (
            .O(N__11800),
            .I(N__11788));
    Span12Mux_v I__2866 (
            .O(N__11797),
            .I(N__11785));
    Span4Mux_h I__2865 (
            .O(N__11794),
            .I(N__11782));
    Span12Mux_h I__2864 (
            .O(N__11791),
            .I(N__11779));
    Span12Mux_v I__2863 (
            .O(N__11788),
            .I(N__11774));
    Span12Mux_h I__2862 (
            .O(N__11785),
            .I(N__11774));
    Span4Mux_v I__2861 (
            .O(N__11782),
            .I(N__11771));
    Odrv12 I__2860 (
            .O(N__11779),
            .I(CASUn_c));
    Odrv12 I__2859 (
            .O(N__11774),
            .I(CASUn_c));
    Odrv4 I__2858 (
            .O(N__11771),
            .I(CASUn_c));
    InMux I__2857 (
            .O(N__11764),
            .I(N__11761));
    LocalMux I__2856 (
            .O(N__11761),
            .I(N__11758));
    Span4Mux_v I__2855 (
            .O(N__11758),
            .I(N__11754));
    InMux I__2854 (
            .O(N__11757),
            .I(N__11751));
    Span4Mux_h I__2853 (
            .O(N__11754),
            .I(N__11748));
    LocalMux I__2852 (
            .O(N__11751),
            .I(N__11745));
    Sp12to4 I__2851 (
            .O(N__11748),
            .I(N__11742));
    Span4Mux_v I__2850 (
            .O(N__11745),
            .I(N__11739));
    Span12Mux_h I__2849 (
            .O(N__11742),
            .I(N__11735));
    Span4Mux_v I__2848 (
            .O(N__11739),
            .I(N__11732));
    InMux I__2847 (
            .O(N__11738),
            .I(N__11729));
    Odrv12 I__2846 (
            .O(N__11735),
            .I(DMA_WRITE_CYCLE));
    Odrv4 I__2845 (
            .O(N__11732),
            .I(DMA_WRITE_CYCLE));
    LocalMux I__2844 (
            .O(N__11729),
            .I(DMA_WRITE_CYCLE));
    IoInMux I__2843 (
            .O(N__11722),
            .I(N__11719));
    LocalMux I__2842 (
            .O(N__11719),
            .I(N__11716));
    Span4Mux_s3_h I__2841 (
            .O(N__11716),
            .I(N__11713));
    Span4Mux_v I__2840 (
            .O(N__11713),
            .I(N__11710));
    Odrv4 I__2839 (
            .O(N__11710),
            .I(N_379));
    InMux I__2838 (
            .O(N__11707),
            .I(N__11704));
    LocalMux I__2837 (
            .O(N__11704),
            .I(N__11700));
    InMux I__2836 (
            .O(N__11703),
            .I(N__11697));
    Span4Mux_v I__2835 (
            .O(N__11700),
            .I(N__11694));
    LocalMux I__2834 (
            .O(N__11697),
            .I(N__11691));
    Span4Mux_h I__2833 (
            .O(N__11694),
            .I(N__11688));
    Span4Mux_v I__2832 (
            .O(N__11691),
            .I(N__11685));
    Odrv4 I__2831 (
            .O(N__11688),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ));
    Odrv4 I__2830 (
            .O(N__11685),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ));
    CascadeMux I__2829 (
            .O(N__11680),
            .I(N_336_cascade_));
    CascadeMux I__2828 (
            .O(N__11677),
            .I(N__11672));
    InMux I__2827 (
            .O(N__11676),
            .I(N__11668));
    InMux I__2826 (
            .O(N__11675),
            .I(N__11665));
    InMux I__2825 (
            .O(N__11672),
            .I(N__11662));
    InMux I__2824 (
            .O(N__11671),
            .I(N__11650));
    LocalMux I__2823 (
            .O(N__11668),
            .I(N__11643));
    LocalMux I__2822 (
            .O(N__11665),
            .I(N__11640));
    LocalMux I__2821 (
            .O(N__11662),
            .I(N__11637));
    InMux I__2820 (
            .O(N__11661),
            .I(N__11630));
    InMux I__2819 (
            .O(N__11660),
            .I(N__11630));
    InMux I__2818 (
            .O(N__11659),
            .I(N__11630));
    InMux I__2817 (
            .O(N__11658),
            .I(N__11625));
    InMux I__2816 (
            .O(N__11657),
            .I(N__11625));
    InMux I__2815 (
            .O(N__11656),
            .I(N__11618));
    InMux I__2814 (
            .O(N__11655),
            .I(N__11618));
    InMux I__2813 (
            .O(N__11654),
            .I(N__11618));
    InMux I__2812 (
            .O(N__11653),
            .I(N__11615));
    LocalMux I__2811 (
            .O(N__11650),
            .I(N__11612));
    InMux I__2810 (
            .O(N__11649),
            .I(N__11607));
    InMux I__2809 (
            .O(N__11648),
            .I(N__11601));
    InMux I__2808 (
            .O(N__11647),
            .I(N__11601));
    InMux I__2807 (
            .O(N__11646),
            .I(N__11598));
    Span4Mux_v I__2806 (
            .O(N__11643),
            .I(N__11587));
    Span4Mux_v I__2805 (
            .O(N__11640),
            .I(N__11587));
    Span4Mux_h I__2804 (
            .O(N__11637),
            .I(N__11587));
    LocalMux I__2803 (
            .O(N__11630),
            .I(N__11587));
    LocalMux I__2802 (
            .O(N__11625),
            .I(N__11587));
    LocalMux I__2801 (
            .O(N__11618),
            .I(N__11584));
    LocalMux I__2800 (
            .O(N__11615),
            .I(N__11581));
    Span4Mux_v I__2799 (
            .O(N__11612),
            .I(N__11577));
    InMux I__2798 (
            .O(N__11611),
            .I(N__11574));
    InMux I__2797 (
            .O(N__11610),
            .I(N__11569));
    LocalMux I__2796 (
            .O(N__11607),
            .I(N__11565));
    InMux I__2795 (
            .O(N__11606),
            .I(N__11562));
    LocalMux I__2794 (
            .O(N__11601),
            .I(N__11553));
    LocalMux I__2793 (
            .O(N__11598),
            .I(N__11553));
    Span4Mux_h I__2792 (
            .O(N__11587),
            .I(N__11553));
    Span4Mux_v I__2791 (
            .O(N__11584),
            .I(N__11553));
    Span4Mux_v I__2790 (
            .O(N__11581),
            .I(N__11550));
    InMux I__2789 (
            .O(N__11580),
            .I(N__11547));
    Span4Mux_h I__2788 (
            .O(N__11577),
            .I(N__11542));
    LocalMux I__2787 (
            .O(N__11574),
            .I(N__11542));
    InMux I__2786 (
            .O(N__11573),
            .I(N__11537));
    InMux I__2785 (
            .O(N__11572),
            .I(N__11537));
    LocalMux I__2784 (
            .O(N__11569),
            .I(N__11534));
    InMux I__2783 (
            .O(N__11568),
            .I(N__11531));
    Span4Mux_v I__2782 (
            .O(N__11565),
            .I(N__11524));
    LocalMux I__2781 (
            .O(N__11562),
            .I(N__11524));
    Span4Mux_v I__2780 (
            .O(N__11553),
            .I(N__11524));
    Odrv4 I__2779 (
            .O(N__11550),
            .I(CPU_CYCLEm));
    LocalMux I__2778 (
            .O(N__11547),
            .I(CPU_CYCLEm));
    Odrv4 I__2777 (
            .O(N__11542),
            .I(CPU_CYCLEm));
    LocalMux I__2776 (
            .O(N__11537),
            .I(CPU_CYCLEm));
    Odrv12 I__2775 (
            .O(N__11534),
            .I(CPU_CYCLEm));
    LocalMux I__2774 (
            .O(N__11531),
            .I(CPU_CYCLEm));
    Odrv4 I__2773 (
            .O(N__11524),
            .I(CPU_CYCLEm));
    IoInMux I__2772 (
            .O(N__11509),
            .I(N__11506));
    LocalMux I__2771 (
            .O(N__11506),
            .I(N__11503));
    Span4Mux_s2_h I__2770 (
            .O(N__11503),
            .I(N__11500));
    Span4Mux_v I__2769 (
            .O(N__11500),
            .I(N__11497));
    Sp12to4 I__2768 (
            .O(N__11497),
            .I(N__11494));
    Span12Mux_h I__2767 (
            .O(N__11494),
            .I(N__11491));
    Odrv12 I__2766 (
            .O(N__11491),
            .I(N_175_i));
    IoInMux I__2765 (
            .O(N__11488),
            .I(N__11485));
    LocalMux I__2764 (
            .O(N__11485),
            .I(N__11482));
    IoSpan4Mux I__2763 (
            .O(N__11482),
            .I(N__11479));
    Span4Mux_s3_v I__2762 (
            .O(N__11479),
            .I(N__11476));
    Odrv4 I__2761 (
            .O(N__11476),
            .I(N_337_i));
    IoInMux I__2760 (
            .O(N__11473),
            .I(N__11470));
    LocalMux I__2759 (
            .O(N__11470),
            .I(N__11467));
    Span4Mux_s3_v I__2758 (
            .O(N__11467),
            .I(N__11464));
    Odrv4 I__2757 (
            .O(N__11464),
            .I(N_336_i));
    IoInMux I__2756 (
            .O(N__11461),
            .I(N__11458));
    LocalMux I__2755 (
            .O(N__11458),
            .I(N__11455));
    Span12Mux_s6_v I__2754 (
            .O(N__11455),
            .I(N__11452));
    Odrv12 I__2753 (
            .O(N__11452),
            .I(N_335_i));
    InMux I__2752 (
            .O(N__11449),
            .I(N__11444));
    InMux I__2751 (
            .O(N__11448),
            .I(N__11441));
    InMux I__2750 (
            .O(N__11447),
            .I(N__11438));
    LocalMux I__2749 (
            .O(N__11444),
            .I(N__11431));
    LocalMux I__2748 (
            .O(N__11441),
            .I(N__11427));
    LocalMux I__2747 (
            .O(N__11438),
            .I(N__11424));
    InMux I__2746 (
            .O(N__11437),
            .I(N__11415));
    InMux I__2745 (
            .O(N__11436),
            .I(N__11415));
    InMux I__2744 (
            .O(N__11435),
            .I(N__11415));
    InMux I__2743 (
            .O(N__11434),
            .I(N__11415));
    Span4Mux_v I__2742 (
            .O(N__11431),
            .I(N__11412));
    InMux I__2741 (
            .O(N__11430),
            .I(N__11409));
    Span4Mux_v I__2740 (
            .O(N__11427),
            .I(N__11406));
    Span4Mux_v I__2739 (
            .O(N__11424),
            .I(N__11403));
    LocalMux I__2738 (
            .O(N__11415),
            .I(N__11400));
    Span4Mux_v I__2737 (
            .O(N__11412),
            .I(N__11397));
    LocalMux I__2736 (
            .O(N__11409),
            .I(N__11394));
    Span4Mux_v I__2735 (
            .O(N__11406),
            .I(N__11387));
    Span4Mux_v I__2734 (
            .O(N__11403),
            .I(N__11387));
    Span4Mux_v I__2733 (
            .O(N__11400),
            .I(N__11387));
    Sp12to4 I__2732 (
            .O(N__11397),
            .I(N__11382));
    Span12Mux_v I__2731 (
            .O(N__11394),
            .I(N__11382));
    Sp12to4 I__2730 (
            .O(N__11387),
            .I(N__11379));
    Span12Mux_h I__2729 (
            .O(N__11382),
            .I(N__11376));
    Span12Mux_h I__2728 (
            .O(N__11379),
            .I(N__11373));
    Odrv12 I__2727 (
            .O(N__11376),
            .I(A_c_1));
    Odrv12 I__2726 (
            .O(N__11373),
            .I(A_c_1));
    InMux I__2725 (
            .O(N__11368),
            .I(N__11353));
    InMux I__2724 (
            .O(N__11367),
            .I(N__11353));
    InMux I__2723 (
            .O(N__11366),
            .I(N__11353));
    InMux I__2722 (
            .O(N__11365),
            .I(N__11353));
    InMux I__2721 (
            .O(N__11364),
            .I(N__11350));
    InMux I__2720 (
            .O(N__11363),
            .I(N__11346));
    CascadeMux I__2719 (
            .O(N__11362),
            .I(N__11343));
    LocalMux I__2718 (
            .O(N__11353),
            .I(N__11339));
    LocalMux I__2717 (
            .O(N__11350),
            .I(N__11336));
    InMux I__2716 (
            .O(N__11349),
            .I(N__11333));
    LocalMux I__2715 (
            .O(N__11346),
            .I(N__11329));
    InMux I__2714 (
            .O(N__11343),
            .I(N__11326));
    InMux I__2713 (
            .O(N__11342),
            .I(N__11323));
    Span4Mux_v I__2712 (
            .O(N__11339),
            .I(N__11318));
    Span4Mux_v I__2711 (
            .O(N__11336),
            .I(N__11318));
    LocalMux I__2710 (
            .O(N__11333),
            .I(N__11315));
    InMux I__2709 (
            .O(N__11332),
            .I(N__11312));
    Span4Mux_v I__2708 (
            .O(N__11329),
            .I(N__11309));
    LocalMux I__2707 (
            .O(N__11326),
            .I(N__11306));
    LocalMux I__2706 (
            .O(N__11323),
            .I(N__11303));
    Span4Mux_h I__2705 (
            .O(N__11318),
            .I(N__11298));
    Span4Mux_v I__2704 (
            .O(N__11315),
            .I(N__11298));
    LocalMux I__2703 (
            .O(N__11312),
            .I(N__11295));
    Sp12to4 I__2702 (
            .O(N__11309),
            .I(N__11290));
    Span12Mux_v I__2701 (
            .O(N__11306),
            .I(N__11290));
    Span4Mux_v I__2700 (
            .O(N__11303),
            .I(N__11287));
    Span4Mux_h I__2699 (
            .O(N__11298),
            .I(N__11282));
    Span4Mux_v I__2698 (
            .O(N__11295),
            .I(N__11282));
    Span12Mux_h I__2697 (
            .O(N__11290),
            .I(N__11279));
    Sp12to4 I__2696 (
            .O(N__11287),
            .I(N__11274));
    Sp12to4 I__2695 (
            .O(N__11282),
            .I(N__11274));
    Odrv12 I__2694 (
            .O(N__11279),
            .I(A_c_0));
    Odrv12 I__2693 (
            .O(N__11274),
            .I(A_c_0));
    CascadeMux I__2692 (
            .O(N__11269),
            .I(N__11266));
    InMux I__2691 (
            .O(N__11266),
            .I(N__11259));
    InMux I__2690 (
            .O(N__11265),
            .I(N__11256));
    CascadeMux I__2689 (
            .O(N__11264),
            .I(N__11250));
    CascadeMux I__2688 (
            .O(N__11263),
            .I(N__11247));
    CascadeMux I__2687 (
            .O(N__11262),
            .I(N__11244));
    LocalMux I__2686 (
            .O(N__11259),
            .I(N__11241));
    LocalMux I__2685 (
            .O(N__11256),
            .I(N__11238));
    InMux I__2684 (
            .O(N__11255),
            .I(N__11229));
    InMux I__2683 (
            .O(N__11254),
            .I(N__11229));
    InMux I__2682 (
            .O(N__11253),
            .I(N__11229));
    InMux I__2681 (
            .O(N__11250),
            .I(N__11229));
    InMux I__2680 (
            .O(N__11247),
            .I(N__11226));
    InMux I__2679 (
            .O(N__11244),
            .I(N__11223));
    Span4Mux_v I__2678 (
            .O(N__11241),
            .I(N__11218));
    Span4Mux_v I__2677 (
            .O(N__11238),
            .I(N__11218));
    LocalMux I__2676 (
            .O(N__11229),
            .I(N__11215));
    LocalMux I__2675 (
            .O(N__11226),
            .I(N__11212));
    LocalMux I__2674 (
            .O(N__11223),
            .I(N__11209));
    Span4Mux_v I__2673 (
            .O(N__11218),
            .I(N__11202));
    Span4Mux_h I__2672 (
            .O(N__11215),
            .I(N__11202));
    Span4Mux_v I__2671 (
            .O(N__11212),
            .I(N__11199));
    Span4Mux_v I__2670 (
            .O(N__11209),
            .I(N__11196));
    InMux I__2669 (
            .O(N__11208),
            .I(N__11193));
    InMux I__2668 (
            .O(N__11207),
            .I(N__11190));
    Span4Mux_h I__2667 (
            .O(N__11202),
            .I(N__11185));
    Span4Mux_v I__2666 (
            .O(N__11199),
            .I(N__11185));
    Span4Mux_h I__2665 (
            .O(N__11196),
            .I(N__11180));
    LocalMux I__2664 (
            .O(N__11193),
            .I(N__11180));
    LocalMux I__2663 (
            .O(N__11190),
            .I(N__11177));
    Span4Mux_v I__2662 (
            .O(N__11185),
            .I(N__11174));
    Span4Mux_h I__2661 (
            .O(N__11180),
            .I(N__11171));
    Span12Mux_v I__2660 (
            .O(N__11177),
            .I(N__11168));
    Span4Mux_h I__2659 (
            .O(N__11174),
            .I(N__11165));
    Sp12to4 I__2658 (
            .O(N__11171),
            .I(N__11162));
    Span12Mux_h I__2657 (
            .O(N__11168),
            .I(N__11159));
    Sp12to4 I__2656 (
            .O(N__11165),
            .I(N__11154));
    Span12Mux_v I__2655 (
            .O(N__11162),
            .I(N__11154));
    Odrv12 I__2654 (
            .O(N__11159),
            .I(SIZ_c_1));
    Odrv12 I__2653 (
            .O(N__11154),
            .I(SIZ_c_1));
    CascadeMux I__2652 (
            .O(N__11149),
            .I(N__11144));
    InMux I__2651 (
            .O(N__11148),
            .I(N__11141));
    InMux I__2650 (
            .O(N__11147),
            .I(N__11135));
    InMux I__2649 (
            .O(N__11144),
            .I(N__11132));
    LocalMux I__2648 (
            .O(N__11141),
            .I(N__11129));
    CascadeMux I__2647 (
            .O(N__11140),
            .I(N__11126));
    CascadeMux I__2646 (
            .O(N__11139),
            .I(N__11123));
    CascadeMux I__2645 (
            .O(N__11138),
            .I(N__11120));
    LocalMux I__2644 (
            .O(N__11135),
            .I(N__11116));
    LocalMux I__2643 (
            .O(N__11132),
            .I(N__11113));
    Span4Mux_v I__2642 (
            .O(N__11129),
            .I(N__11110));
    InMux I__2641 (
            .O(N__11126),
            .I(N__11101));
    InMux I__2640 (
            .O(N__11123),
            .I(N__11101));
    InMux I__2639 (
            .O(N__11120),
            .I(N__11101));
    InMux I__2638 (
            .O(N__11119),
            .I(N__11101));
    Span4Mux_v I__2637 (
            .O(N__11116),
            .I(N__11097));
    Span4Mux_v I__2636 (
            .O(N__11113),
            .I(N__11093));
    Span4Mux_v I__2635 (
            .O(N__11110),
            .I(N__11088));
    LocalMux I__2634 (
            .O(N__11101),
            .I(N__11088));
    CascadeMux I__2633 (
            .O(N__11100),
            .I(N__11084));
    Span4Mux_v I__2632 (
            .O(N__11097),
            .I(N__11081));
    InMux I__2631 (
            .O(N__11096),
            .I(N__11078));
    Span4Mux_v I__2630 (
            .O(N__11093),
            .I(N__11073));
    Span4Mux_h I__2629 (
            .O(N__11088),
            .I(N__11073));
    InMux I__2628 (
            .O(N__11087),
            .I(N__11070));
    InMux I__2627 (
            .O(N__11084),
            .I(N__11067));
    Span4Mux_v I__2626 (
            .O(N__11081),
            .I(N__11064));
    LocalMux I__2625 (
            .O(N__11078),
            .I(N__11061));
    Span4Mux_v I__2624 (
            .O(N__11073),
            .I(N__11058));
    LocalMux I__2623 (
            .O(N__11070),
            .I(N__11053));
    LocalMux I__2622 (
            .O(N__11067),
            .I(N__11053));
    Sp12to4 I__2621 (
            .O(N__11064),
            .I(N__11048));
    Span12Mux_v I__2620 (
            .O(N__11061),
            .I(N__11048));
    Span4Mux_h I__2619 (
            .O(N__11058),
            .I(N__11045));
    Sp12to4 I__2618 (
            .O(N__11053),
            .I(N__11042));
    Span12Mux_h I__2617 (
            .O(N__11048),
            .I(N__11039));
    Sp12to4 I__2616 (
            .O(N__11045),
            .I(N__11034));
    Span12Mux_v I__2615 (
            .O(N__11042),
            .I(N__11034));
    Odrv12 I__2614 (
            .O(N__11039),
            .I(SIZ_c_0));
    Odrv12 I__2613 (
            .O(N__11034),
            .I(SIZ_c_0));
    IoInMux I__2612 (
            .O(N__11029),
            .I(N__11026));
    LocalMux I__2611 (
            .O(N__11026),
            .I(N__11023));
    Span4Mux_s2_v I__2610 (
            .O(N__11023),
            .I(N__11020));
    Span4Mux_h I__2609 (
            .O(N__11020),
            .I(N__11017));
    Span4Mux_v I__2608 (
            .O(N__11017),
            .I(N__11014));
    Odrv4 I__2607 (
            .O(N__11014),
            .I(N_334_i));
    InMux I__2606 (
            .O(N__11011),
            .I(N__11007));
    InMux I__2605 (
            .O(N__11010),
            .I(N__11003));
    LocalMux I__2604 (
            .O(N__11007),
            .I(N__11000));
    InMux I__2603 (
            .O(N__11006),
            .I(N__10997));
    LocalMux I__2602 (
            .O(N__11003),
            .I(N__10989));
    Span4Mux_h I__2601 (
            .O(N__11000),
            .I(N__10989));
    LocalMux I__2600 (
            .O(N__10997),
            .I(N__10989));
    InMux I__2599 (
            .O(N__10996),
            .I(N__10986));
    Span4Mux_v I__2598 (
            .O(N__10989),
            .I(N__10983));
    LocalMux I__2597 (
            .O(N__10986),
            .I(N__10980));
    Span4Mux_v I__2596 (
            .O(N__10983),
            .I(N__10977));
    Sp12to4 I__2595 (
            .O(N__10980),
            .I(N__10974));
    Sp12to4 I__2594 (
            .O(N__10977),
            .I(N__10971));
    Span12Mux_v I__2593 (
            .O(N__10974),
            .I(N__10968));
    Span12Mux_h I__2592 (
            .O(N__10971),
            .I(N__10965));
    Span12Mux_h I__2591 (
            .O(N__10968),
            .I(N__10962));
    Odrv12 I__2590 (
            .O(N__10965),
            .I(DRA_c_4));
    Odrv12 I__2589 (
            .O(N__10962),
            .I(DRA_c_4));
    InMux I__2588 (
            .O(N__10957),
            .I(N__10951));
    InMux I__2587 (
            .O(N__10956),
            .I(N__10951));
    LocalMux I__2586 (
            .O(N__10951),
            .I(N__10946));
    InMux I__2585 (
            .O(N__10950),
            .I(N__10943));
    InMux I__2584 (
            .O(N__10949),
            .I(N__10940));
    Span4Mux_h I__2583 (
            .O(N__10946),
            .I(N__10933));
    LocalMux I__2582 (
            .O(N__10943),
            .I(N__10933));
    LocalMux I__2581 (
            .O(N__10940),
            .I(N__10933));
    Span4Mux_h I__2580 (
            .O(N__10933),
            .I(N__10930));
    Sp12to4 I__2579 (
            .O(N__10930),
            .I(N__10927));
    Span12Mux_v I__2578 (
            .O(N__10927),
            .I(N__10924));
    Odrv12 I__2577 (
            .O(N__10924),
            .I(DRA_c_3));
    InMux I__2576 (
            .O(N__10921),
            .I(N__10918));
    LocalMux I__2575 (
            .O(N__10918),
            .I(N__10915));
    Odrv12 I__2574 (
            .O(N__10915),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__2573 (
            .O(N__10912),
            .I(N__10908));
    InMux I__2572 (
            .O(N__10911),
            .I(N__10905));
    LocalMux I__2571 (
            .O(N__10908),
            .I(N__10899));
    LocalMux I__2570 (
            .O(N__10905),
            .I(N__10899));
    InMux I__2569 (
            .O(N__10904),
            .I(N__10896));
    Span4Mux_v I__2568 (
            .O(N__10899),
            .I(N__10892));
    LocalMux I__2567 (
            .O(N__10896),
            .I(N__10889));
    InMux I__2566 (
            .O(N__10895),
            .I(N__10886));
    Span4Mux_v I__2565 (
            .O(N__10892),
            .I(N__10883));
    Sp12to4 I__2564 (
            .O(N__10889),
            .I(N__10878));
    LocalMux I__2563 (
            .O(N__10886),
            .I(N__10878));
    Sp12to4 I__2562 (
            .O(N__10883),
            .I(N__10873));
    Span12Mux_v I__2561 (
            .O(N__10878),
            .I(N__10873));
    Span12Mux_h I__2560 (
            .O(N__10873),
            .I(N__10870));
    Odrv12 I__2559 (
            .O(N__10870),
            .I(DRA_c_6));
    CascadeMux I__2558 (
            .O(N__10867),
            .I(N__10864));
    InMux I__2557 (
            .O(N__10864),
            .I(N__10858));
    CascadeMux I__2556 (
            .O(N__10863),
            .I(N__10854));
    InMux I__2555 (
            .O(N__10862),
            .I(N__10843));
    InMux I__2554 (
            .O(N__10861),
            .I(N__10840));
    LocalMux I__2553 (
            .O(N__10858),
            .I(N__10834));
    InMux I__2552 (
            .O(N__10857),
            .I(N__10825));
    InMux I__2551 (
            .O(N__10854),
            .I(N__10825));
    InMux I__2550 (
            .O(N__10853),
            .I(N__10825));
    InMux I__2549 (
            .O(N__10852),
            .I(N__10825));
    InMux I__2548 (
            .O(N__10851),
            .I(N__10822));
    InMux I__2547 (
            .O(N__10850),
            .I(N__10817));
    InMux I__2546 (
            .O(N__10849),
            .I(N__10817));
    InMux I__2545 (
            .O(N__10848),
            .I(N__10814));
    InMux I__2544 (
            .O(N__10847),
            .I(N__10809));
    InMux I__2543 (
            .O(N__10846),
            .I(N__10809));
    LocalMux I__2542 (
            .O(N__10843),
            .I(N__10804));
    LocalMux I__2541 (
            .O(N__10840),
            .I(N__10804));
    InMux I__2540 (
            .O(N__10839),
            .I(N__10801));
    InMux I__2539 (
            .O(N__10838),
            .I(N__10796));
    InMux I__2538 (
            .O(N__10837),
            .I(N__10796));
    Span4Mux_v I__2537 (
            .O(N__10834),
            .I(N__10792));
    LocalMux I__2536 (
            .O(N__10825),
            .I(N__10781));
    LocalMux I__2535 (
            .O(N__10822),
            .I(N__10781));
    LocalMux I__2534 (
            .O(N__10817),
            .I(N__10781));
    LocalMux I__2533 (
            .O(N__10814),
            .I(N__10781));
    LocalMux I__2532 (
            .O(N__10809),
            .I(N__10781));
    Span4Mux_v I__2531 (
            .O(N__10804),
            .I(N__10778));
    LocalMux I__2530 (
            .O(N__10801),
            .I(N__10775));
    LocalMux I__2529 (
            .O(N__10796),
            .I(N__10768));
    InMux I__2528 (
            .O(N__10795),
            .I(N__10765));
    Span4Mux_h I__2527 (
            .O(N__10792),
            .I(N__10760));
    Span4Mux_v I__2526 (
            .O(N__10781),
            .I(N__10760));
    Span4Mux_h I__2525 (
            .O(N__10778),
            .I(N__10755));
    Span4Mux_v I__2524 (
            .O(N__10775),
            .I(N__10755));
    InMux I__2523 (
            .O(N__10774),
            .I(N__10752));
    InMux I__2522 (
            .O(N__10773),
            .I(N__10749));
    InMux I__2521 (
            .O(N__10772),
            .I(N__10746));
    InMux I__2520 (
            .O(N__10771),
            .I(N__10743));
    Span4Mux_v I__2519 (
            .O(N__10768),
            .I(N__10738));
    LocalMux I__2518 (
            .O(N__10765),
            .I(N__10738));
    Sp12to4 I__2517 (
            .O(N__10760),
            .I(N__10733));
    Sp12to4 I__2516 (
            .O(N__10755),
            .I(N__10733));
    LocalMux I__2515 (
            .O(N__10752),
            .I(N__10728));
    LocalMux I__2514 (
            .O(N__10749),
            .I(N__10728));
    LocalMux I__2513 (
            .O(N__10746),
            .I(N__10723));
    LocalMux I__2512 (
            .O(N__10743),
            .I(N__10723));
    Sp12to4 I__2511 (
            .O(N__10738),
            .I(N__10720));
    Span12Mux_h I__2510 (
            .O(N__10733),
            .I(N__10717));
    Span12Mux_h I__2509 (
            .O(N__10728),
            .I(N__10714));
    Span12Mux_v I__2508 (
            .O(N__10723),
            .I(N__10711));
    Span12Mux_v I__2507 (
            .O(N__10720),
            .I(N__10708));
    Span12Mux_v I__2506 (
            .O(N__10717),
            .I(N__10705));
    Span12Mux_v I__2505 (
            .O(N__10714),
            .I(N__10700));
    Span12Mux_h I__2504 (
            .O(N__10711),
            .I(N__10700));
    Span12Mux_h I__2503 (
            .O(N__10708),
            .I(N__10697));
    Odrv12 I__2502 (
            .O(N__10705),
            .I(AGNUS_REV_c));
    Odrv12 I__2501 (
            .O(N__10700),
            .I(AGNUS_REV_c));
    Odrv12 I__2500 (
            .O(N__10697),
            .I(AGNUS_REV_c));
    InMux I__2499 (
            .O(N__10690),
            .I(N__10684));
    InMux I__2498 (
            .O(N__10689),
            .I(N__10681));
    InMux I__2497 (
            .O(N__10688),
            .I(N__10678));
    InMux I__2496 (
            .O(N__10687),
            .I(N__10675));
    LocalMux I__2495 (
            .O(N__10684),
            .I(N__10668));
    LocalMux I__2494 (
            .O(N__10681),
            .I(N__10668));
    LocalMux I__2493 (
            .O(N__10678),
            .I(N__10668));
    LocalMux I__2492 (
            .O(N__10675),
            .I(N__10665));
    Span4Mux_v I__2491 (
            .O(N__10668),
            .I(N__10662));
    Span4Mux_v I__2490 (
            .O(N__10665),
            .I(N__10659));
    Sp12to4 I__2489 (
            .O(N__10662),
            .I(N__10656));
    Span4Mux_h I__2488 (
            .O(N__10659),
            .I(N__10653));
    Span12Mux_h I__2487 (
            .O(N__10656),
            .I(N__10648));
    Sp12to4 I__2486 (
            .O(N__10653),
            .I(N__10648));
    Odrv12 I__2485 (
            .O(N__10648),
            .I(DRA_c_7));
    InMux I__2484 (
            .O(N__10645),
            .I(N__10642));
    LocalMux I__2483 (
            .O(N__10642),
            .I(N__10639));
    Span4Mux_h I__2482 (
            .O(N__10639),
            .I(N__10636));
    Odrv4 I__2481 (
            .O(N__10636),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    ClkMux I__2480 (
            .O(N__10633),
            .I(N__10615));
    ClkMux I__2479 (
            .O(N__10632),
            .I(N__10615));
    ClkMux I__2478 (
            .O(N__10631),
            .I(N__10615));
    ClkMux I__2477 (
            .O(N__10630),
            .I(N__10615));
    ClkMux I__2476 (
            .O(N__10629),
            .I(N__10615));
    ClkMux I__2475 (
            .O(N__10628),
            .I(N__10615));
    GlobalMux I__2474 (
            .O(N__10615),
            .I(N__10612));
    gio2CtrlBuf I__2473 (
            .O(N__10612),
            .I(C3_c_g));
    CEMux I__2472 (
            .O(N__10609),
            .I(N__10573));
    CEMux I__2471 (
            .O(N__10608),
            .I(N__10573));
    CEMux I__2470 (
            .O(N__10607),
            .I(N__10573));
    CEMux I__2469 (
            .O(N__10606),
            .I(N__10573));
    CEMux I__2468 (
            .O(N__10605),
            .I(N__10573));
    CEMux I__2467 (
            .O(N__10604),
            .I(N__10573));
    CEMux I__2466 (
            .O(N__10603),
            .I(N__10573));
    CEMux I__2465 (
            .O(N__10602),
            .I(N__10573));
    CEMux I__2464 (
            .O(N__10601),
            .I(N__10573));
    CEMux I__2463 (
            .O(N__10600),
            .I(N__10573));
    CEMux I__2462 (
            .O(N__10599),
            .I(N__10573));
    CEMux I__2461 (
            .O(N__10598),
            .I(N__10573));
    GlobalMux I__2460 (
            .O(N__10573),
            .I(N__10570));
    gio2CtrlBuf I__2459 (
            .O(N__10570),
            .I(DBRn_c_i_0_g));
    InMux I__2458 (
            .O(N__10567),
            .I(N__10559));
    InMux I__2457 (
            .O(N__10566),
            .I(N__10556));
    InMux I__2456 (
            .O(N__10565),
            .I(N__10553));
    InMux I__2455 (
            .O(N__10564),
            .I(N__10550));
    InMux I__2454 (
            .O(N__10563),
            .I(N__10547));
    InMux I__2453 (
            .O(N__10562),
            .I(N__10544));
    LocalMux I__2452 (
            .O(N__10559),
            .I(N__10541));
    LocalMux I__2451 (
            .O(N__10556),
            .I(N__10536));
    LocalMux I__2450 (
            .O(N__10553),
            .I(N__10532));
    LocalMux I__2449 (
            .O(N__10550),
            .I(N__10525));
    LocalMux I__2448 (
            .O(N__10547),
            .I(N__10519));
    LocalMux I__2447 (
            .O(N__10544),
            .I(N__10490));
    Glb2LocalMux I__2446 (
            .O(N__10541),
            .I(N__10396));
    SRMux I__2445 (
            .O(N__10540),
            .I(N__10396));
    SRMux I__2444 (
            .O(N__10539),
            .I(N__10396));
    Glb2LocalMux I__2443 (
            .O(N__10536),
            .I(N__10396));
    SRMux I__2442 (
            .O(N__10535),
            .I(N__10396));
    Glb2LocalMux I__2441 (
            .O(N__10532),
            .I(N__10396));
    SRMux I__2440 (
            .O(N__10531),
            .I(N__10396));
    SRMux I__2439 (
            .O(N__10530),
            .I(N__10396));
    SRMux I__2438 (
            .O(N__10529),
            .I(N__10396));
    SRMux I__2437 (
            .O(N__10528),
            .I(N__10396));
    Glb2LocalMux I__2436 (
            .O(N__10525),
            .I(N__10396));
    SRMux I__2435 (
            .O(N__10524),
            .I(N__10396));
    SRMux I__2434 (
            .O(N__10523),
            .I(N__10396));
    SRMux I__2433 (
            .O(N__10522),
            .I(N__10396));
    Glb2LocalMux I__2432 (
            .O(N__10519),
            .I(N__10396));
    SRMux I__2431 (
            .O(N__10518),
            .I(N__10396));
    SRMux I__2430 (
            .O(N__10517),
            .I(N__10396));
    SRMux I__2429 (
            .O(N__10516),
            .I(N__10396));
    SRMux I__2428 (
            .O(N__10515),
            .I(N__10396));
    SRMux I__2427 (
            .O(N__10514),
            .I(N__10396));
    SRMux I__2426 (
            .O(N__10513),
            .I(N__10396));
    SRMux I__2425 (
            .O(N__10512),
            .I(N__10396));
    SRMux I__2424 (
            .O(N__10511),
            .I(N__10396));
    SRMux I__2423 (
            .O(N__10510),
            .I(N__10396));
    SRMux I__2422 (
            .O(N__10509),
            .I(N__10396));
    SRMux I__2421 (
            .O(N__10508),
            .I(N__10396));
    SRMux I__2420 (
            .O(N__10507),
            .I(N__10396));
    SRMux I__2419 (
            .O(N__10506),
            .I(N__10396));
    SRMux I__2418 (
            .O(N__10505),
            .I(N__10396));
    SRMux I__2417 (
            .O(N__10504),
            .I(N__10396));
    SRMux I__2416 (
            .O(N__10503),
            .I(N__10396));
    SRMux I__2415 (
            .O(N__10502),
            .I(N__10396));
    SRMux I__2414 (
            .O(N__10501),
            .I(N__10396));
    SRMux I__2413 (
            .O(N__10500),
            .I(N__10396));
    SRMux I__2412 (
            .O(N__10499),
            .I(N__10396));
    SRMux I__2411 (
            .O(N__10498),
            .I(N__10396));
    SRMux I__2410 (
            .O(N__10497),
            .I(N__10396));
    SRMux I__2409 (
            .O(N__10496),
            .I(N__10396));
    SRMux I__2408 (
            .O(N__10495),
            .I(N__10396));
    SRMux I__2407 (
            .O(N__10494),
            .I(N__10396));
    SRMux I__2406 (
            .O(N__10493),
            .I(N__10396));
    Glb2LocalMux I__2405 (
            .O(N__10490),
            .I(N__10396));
    SRMux I__2404 (
            .O(N__10489),
            .I(N__10396));
    SRMux I__2403 (
            .O(N__10488),
            .I(N__10396));
    SRMux I__2402 (
            .O(N__10487),
            .I(N__10396));
    GlobalMux I__2401 (
            .O(N__10396),
            .I(N__10393));
    gio2CtrlBuf I__2400 (
            .O(N__10393),
            .I(RESETn_c_i_g));
    InMux I__2399 (
            .O(N__10390),
            .I(N__10386));
    InMux I__2398 (
            .O(N__10389),
            .I(N__10381));
    LocalMux I__2397 (
            .O(N__10386),
            .I(N__10377));
    InMux I__2396 (
            .O(N__10385),
            .I(N__10374));
    InMux I__2395 (
            .O(N__10384),
            .I(N__10371));
    LocalMux I__2394 (
            .O(N__10381),
            .I(N__10368));
    InMux I__2393 (
            .O(N__10380),
            .I(N__10365));
    Span4Mux_v I__2392 (
            .O(N__10377),
            .I(N__10362));
    LocalMux I__2391 (
            .O(N__10374),
            .I(N__10357));
    LocalMux I__2390 (
            .O(N__10371),
            .I(N__10357));
    Sp12to4 I__2389 (
            .O(N__10368),
            .I(N__10354));
    LocalMux I__2388 (
            .O(N__10365),
            .I(N__10351));
    Sp12to4 I__2387 (
            .O(N__10362),
            .I(N__10348));
    Span4Mux_v I__2386 (
            .O(N__10357),
            .I(N__10345));
    Span12Mux_h I__2385 (
            .O(N__10354),
            .I(N__10342));
    Span12Mux_h I__2384 (
            .O(N__10351),
            .I(N__10339));
    Span12Mux_h I__2383 (
            .O(N__10348),
            .I(N__10334));
    Sp12to4 I__2382 (
            .O(N__10345),
            .I(N__10334));
    Span12Mux_v I__2381 (
            .O(N__10342),
            .I(N__10331));
    Span12Mux_v I__2380 (
            .O(N__10339),
            .I(N__10328));
    Span12Mux_h I__2379 (
            .O(N__10334),
            .I(N__10325));
    Odrv12 I__2378 (
            .O(N__10331),
            .I(RnW_c));
    Odrv12 I__2377 (
            .O(N__10328),
            .I(RnW_c));
    Odrv12 I__2376 (
            .O(N__10325),
            .I(RnW_c));
    CascadeMux I__2375 (
            .O(N__10318),
            .I(N__10315));
    InMux I__2374 (
            .O(N__10315),
            .I(N__10310));
    InMux I__2373 (
            .O(N__10314),
            .I(N__10305));
    InMux I__2372 (
            .O(N__10313),
            .I(N__10305));
    LocalMux I__2371 (
            .O(N__10310),
            .I(N__10300));
    LocalMux I__2370 (
            .O(N__10305),
            .I(N__10300));
    Span4Mux_v I__2369 (
            .O(N__10300),
            .I(N__10295));
    InMux I__2368 (
            .O(N__10299),
            .I(N__10292));
    InMux I__2367 (
            .O(N__10298),
            .I(N__10289));
    Span4Mux_v I__2366 (
            .O(N__10295),
            .I(N__10284));
    LocalMux I__2365 (
            .O(N__10292),
            .I(N__10284));
    LocalMux I__2364 (
            .O(N__10289),
            .I(N__10281));
    Span4Mux_v I__2363 (
            .O(N__10284),
            .I(N__10278));
    Span4Mux_v I__2362 (
            .O(N__10281),
            .I(N__10275));
    Span4Mux_v I__2361 (
            .O(N__10278),
            .I(N__10271));
    Sp12to4 I__2360 (
            .O(N__10275),
            .I(N__10268));
    InMux I__2359 (
            .O(N__10274),
            .I(N__10265));
    Sp12to4 I__2358 (
            .O(N__10271),
            .I(N__10262));
    Span12Mux_h I__2357 (
            .O(N__10268),
            .I(N__10257));
    LocalMux I__2356 (
            .O(N__10265),
            .I(N__10257));
    Span12Mux_h I__2355 (
            .O(N__10262),
            .I(N__10252));
    Span12Mux_v I__2354 (
            .O(N__10257),
            .I(N__10252));
    Odrv12 I__2353 (
            .O(N__10252),
            .I(CASLn_c));
    InMux I__2352 (
            .O(N__10249),
            .I(N__10246));
    LocalMux I__2351 (
            .O(N__10246),
            .I(N__10243));
    Span12Mux_h I__2350 (
            .O(N__10243),
            .I(N__10240));
    Odrv12 I__2349 (
            .O(N__10240),
            .I(RAS1n_c));
    InMux I__2348 (
            .O(N__10237),
            .I(N__10234));
    LocalMux I__2347 (
            .O(N__10234),
            .I(N__10231));
    Span4Mux_v I__2346 (
            .O(N__10231),
            .I(N__10227));
    InMux I__2345 (
            .O(N__10230),
            .I(N__10224));
    Sp12to4 I__2344 (
            .O(N__10227),
            .I(N__10219));
    LocalMux I__2343 (
            .O(N__10224),
            .I(N__10219));
    Span12Mux_h I__2342 (
            .O(N__10219),
            .I(N__10216));
    Odrv12 I__2341 (
            .O(N__10216),
            .I(RAS0n_c));
    InMux I__2340 (
            .O(N__10213),
            .I(N__10210));
    LocalMux I__2339 (
            .O(N__10210),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2338 (
            .O(N__10207),
            .I(N__10203));
    CascadeMux I__2337 (
            .O(N__10206),
            .I(N__10194));
    LocalMux I__2336 (
            .O(N__10203),
            .I(N__10190));
    InMux I__2335 (
            .O(N__10202),
            .I(N__10187));
    InMux I__2334 (
            .O(N__10201),
            .I(N__10184));
    InMux I__2333 (
            .O(N__10200),
            .I(N__10178));
    InMux I__2332 (
            .O(N__10199),
            .I(N__10178));
    InMux I__2331 (
            .O(N__10198),
            .I(N__10175));
    CascadeMux I__2330 (
            .O(N__10197),
            .I(N__10167));
    InMux I__2329 (
            .O(N__10194),
            .I(N__10154));
    InMux I__2328 (
            .O(N__10193),
            .I(N__10154));
    Span4Mux_v I__2327 (
            .O(N__10190),
            .I(N__10145));
    LocalMux I__2326 (
            .O(N__10187),
            .I(N__10145));
    LocalMux I__2325 (
            .O(N__10184),
            .I(N__10145));
    InMux I__2324 (
            .O(N__10183),
            .I(N__10142));
    LocalMux I__2323 (
            .O(N__10178),
            .I(N__10136));
    LocalMux I__2322 (
            .O(N__10175),
            .I(N__10136));
    InMux I__2321 (
            .O(N__10174),
            .I(N__10131));
    InMux I__2320 (
            .O(N__10173),
            .I(N__10131));
    InMux I__2319 (
            .O(N__10172),
            .I(N__10128));
    InMux I__2318 (
            .O(N__10171),
            .I(N__10121));
    InMux I__2317 (
            .O(N__10170),
            .I(N__10121));
    InMux I__2316 (
            .O(N__10167),
            .I(N__10121));
    InMux I__2315 (
            .O(N__10166),
            .I(N__10118));
    InMux I__2314 (
            .O(N__10165),
            .I(N__10113));
    InMux I__2313 (
            .O(N__10164),
            .I(N__10113));
    InMux I__2312 (
            .O(N__10163),
            .I(N__10104));
    InMux I__2311 (
            .O(N__10162),
            .I(N__10104));
    InMux I__2310 (
            .O(N__10161),
            .I(N__10104));
    InMux I__2309 (
            .O(N__10160),
            .I(N__10104));
    InMux I__2308 (
            .O(N__10159),
            .I(N__10098));
    LocalMux I__2307 (
            .O(N__10154),
            .I(N__10095));
    InMux I__2306 (
            .O(N__10153),
            .I(N__10092));
    InMux I__2305 (
            .O(N__10152),
            .I(N__10089));
    Span4Mux_v I__2304 (
            .O(N__10145),
            .I(N__10083));
    LocalMux I__2303 (
            .O(N__10142),
            .I(N__10083));
    InMux I__2302 (
            .O(N__10141),
            .I(N__10080));
    Span4Mux_h I__2301 (
            .O(N__10136),
            .I(N__10071));
    LocalMux I__2300 (
            .O(N__10131),
            .I(N__10071));
    LocalMux I__2299 (
            .O(N__10128),
            .I(N__10071));
    LocalMux I__2298 (
            .O(N__10121),
            .I(N__10071));
    LocalMux I__2297 (
            .O(N__10118),
            .I(N__10064));
    LocalMux I__2296 (
            .O(N__10113),
            .I(N__10064));
    LocalMux I__2295 (
            .O(N__10104),
            .I(N__10064));
    InMux I__2294 (
            .O(N__10103),
            .I(N__10057));
    InMux I__2293 (
            .O(N__10102),
            .I(N__10057));
    InMux I__2292 (
            .O(N__10101),
            .I(N__10057));
    LocalMux I__2291 (
            .O(N__10098),
            .I(N__10052));
    Span4Mux_h I__2290 (
            .O(N__10095),
            .I(N__10045));
    LocalMux I__2289 (
            .O(N__10092),
            .I(N__10045));
    LocalMux I__2288 (
            .O(N__10089),
            .I(N__10045));
    InMux I__2287 (
            .O(N__10088),
            .I(N__10042));
    Span4Mux_h I__2286 (
            .O(N__10083),
            .I(N__10037));
    LocalMux I__2285 (
            .O(N__10080),
            .I(N__10037));
    Span4Mux_v I__2284 (
            .O(N__10071),
            .I(N__10032));
    Span4Mux_v I__2283 (
            .O(N__10064),
            .I(N__10032));
    LocalMux I__2282 (
            .O(N__10057),
            .I(N__10029));
    InMux I__2281 (
            .O(N__10056),
            .I(N__10024));
    InMux I__2280 (
            .O(N__10055),
            .I(N__10024));
    Span4Mux_v I__2279 (
            .O(N__10052),
            .I(N__10019));
    Span4Mux_v I__2278 (
            .O(N__10045),
            .I(N__10019));
    LocalMux I__2277 (
            .O(N__10042),
            .I(N__10014));
    Sp12to4 I__2276 (
            .O(N__10037),
            .I(N__10014));
    Span4Mux_h I__2275 (
            .O(N__10032),
            .I(N__10009));
    Span4Mux_v I__2274 (
            .O(N__10029),
            .I(N__10009));
    LocalMux I__2273 (
            .O(N__10024),
            .I(N__10006));
    Sp12to4 I__2272 (
            .O(N__10019),
            .I(N__9999));
    Span12Mux_v I__2271 (
            .O(N__10014),
            .I(N__9999));
    Sp12to4 I__2270 (
            .O(N__10009),
            .I(N__9999));
    Span12Mux_h I__2269 (
            .O(N__10006),
            .I(N__9996));
    Span12Mux_h I__2268 (
            .O(N__9999),
            .I(N__9993));
    Odrv12 I__2267 (
            .O(N__9996),
            .I(RESETn_c));
    Odrv12 I__2266 (
            .O(N__9993),
            .I(RESETn_c));
    InMux I__2265 (
            .O(N__9988),
            .I(N__9985));
    LocalMux I__2264 (
            .O(N__9985),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__2263 (
            .O(N__9982),
            .I(N__9979));
    LocalMux I__2262 (
            .O(N__9979),
            .I(N__9976));
    Odrv12 I__2261 (
            .O(N__9976),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ));
    InMux I__2260 (
            .O(N__9973),
            .I(N__9970));
    LocalMux I__2259 (
            .O(N__9970),
            .I(N__9931));
    ClkMux I__2258 (
            .O(N__9969),
            .I(N__9832));
    ClkMux I__2257 (
            .O(N__9968),
            .I(N__9832));
    ClkMux I__2256 (
            .O(N__9967),
            .I(N__9832));
    ClkMux I__2255 (
            .O(N__9966),
            .I(N__9832));
    ClkMux I__2254 (
            .O(N__9965),
            .I(N__9832));
    ClkMux I__2253 (
            .O(N__9964),
            .I(N__9832));
    ClkMux I__2252 (
            .O(N__9963),
            .I(N__9832));
    ClkMux I__2251 (
            .O(N__9962),
            .I(N__9832));
    ClkMux I__2250 (
            .O(N__9961),
            .I(N__9832));
    ClkMux I__2249 (
            .O(N__9960),
            .I(N__9832));
    ClkMux I__2248 (
            .O(N__9959),
            .I(N__9832));
    ClkMux I__2247 (
            .O(N__9958),
            .I(N__9832));
    ClkMux I__2246 (
            .O(N__9957),
            .I(N__9832));
    ClkMux I__2245 (
            .O(N__9956),
            .I(N__9832));
    ClkMux I__2244 (
            .O(N__9955),
            .I(N__9832));
    ClkMux I__2243 (
            .O(N__9954),
            .I(N__9832));
    ClkMux I__2242 (
            .O(N__9953),
            .I(N__9832));
    ClkMux I__2241 (
            .O(N__9952),
            .I(N__9832));
    ClkMux I__2240 (
            .O(N__9951),
            .I(N__9832));
    ClkMux I__2239 (
            .O(N__9950),
            .I(N__9832));
    ClkMux I__2238 (
            .O(N__9949),
            .I(N__9832));
    ClkMux I__2237 (
            .O(N__9948),
            .I(N__9832));
    ClkMux I__2236 (
            .O(N__9947),
            .I(N__9832));
    ClkMux I__2235 (
            .O(N__9946),
            .I(N__9832));
    ClkMux I__2234 (
            .O(N__9945),
            .I(N__9832));
    ClkMux I__2233 (
            .O(N__9944),
            .I(N__9832));
    ClkMux I__2232 (
            .O(N__9943),
            .I(N__9832));
    ClkMux I__2231 (
            .O(N__9942),
            .I(N__9832));
    ClkMux I__2230 (
            .O(N__9941),
            .I(N__9832));
    ClkMux I__2229 (
            .O(N__9940),
            .I(N__9832));
    ClkMux I__2228 (
            .O(N__9939),
            .I(N__9832));
    ClkMux I__2227 (
            .O(N__9938),
            .I(N__9832));
    ClkMux I__2226 (
            .O(N__9937),
            .I(N__9832));
    ClkMux I__2225 (
            .O(N__9936),
            .I(N__9832));
    ClkMux I__2224 (
            .O(N__9935),
            .I(N__9832));
    ClkMux I__2223 (
            .O(N__9934),
            .I(N__9832));
    Glb2LocalMux I__2222 (
            .O(N__9931),
            .I(N__9832));
    ClkMux I__2221 (
            .O(N__9930),
            .I(N__9832));
    ClkMux I__2220 (
            .O(N__9929),
            .I(N__9832));
    ClkMux I__2219 (
            .O(N__9928),
            .I(N__9832));
    ClkMux I__2218 (
            .O(N__9927),
            .I(N__9832));
    ClkMux I__2217 (
            .O(N__9926),
            .I(N__9832));
    ClkMux I__2216 (
            .O(N__9925),
            .I(N__9832));
    ClkMux I__2215 (
            .O(N__9924),
            .I(N__9832));
    ClkMux I__2214 (
            .O(N__9923),
            .I(N__9832));
    GlobalMux I__2213 (
            .O(N__9832),
            .I(CLK80_PLL));
    InMux I__2212 (
            .O(N__9829),
            .I(N__9823));
    InMux I__2211 (
            .O(N__9828),
            .I(N__9823));
    LocalMux I__2210 (
            .O(N__9823),
            .I(N__9818));
    InMux I__2209 (
            .O(N__9822),
            .I(N__9815));
    InMux I__2208 (
            .O(N__9821),
            .I(N__9812));
    Span4Mux_v I__2207 (
            .O(N__9818),
            .I(N__9809));
    LocalMux I__2206 (
            .O(N__9815),
            .I(N__9806));
    LocalMux I__2205 (
            .O(N__9812),
            .I(N__9803));
    Sp12to4 I__2204 (
            .O(N__9809),
            .I(N__9800));
    Sp12to4 I__2203 (
            .O(N__9806),
            .I(N__9797));
    Span12Mux_h I__2202 (
            .O(N__9803),
            .I(N__9794));
    Span12Mux_h I__2201 (
            .O(N__9800),
            .I(N__9791));
    Span12Mux_v I__2200 (
            .O(N__9797),
            .I(N__9788));
    Span12Mux_v I__2199 (
            .O(N__9794),
            .I(N__9785));
    Span12Mux_v I__2198 (
            .O(N__9791),
            .I(N__9780));
    Span12Mux_h I__2197 (
            .O(N__9788),
            .I(N__9780));
    Odrv12 I__2196 (
            .O(N__9785),
            .I(DRA_c_1));
    Odrv12 I__2195 (
            .O(N__9780),
            .I(DRA_c_1));
    InMux I__2194 (
            .O(N__9775),
            .I(N__9771));
    InMux I__2193 (
            .O(N__9774),
            .I(N__9768));
    LocalMux I__2192 (
            .O(N__9771),
            .I(N__9763));
    LocalMux I__2191 (
            .O(N__9768),
            .I(N__9763));
    Span12Mux_h I__2190 (
            .O(N__9763),
            .I(N__9760));
    Span12Mux_v I__2189 (
            .O(N__9760),
            .I(N__9757));
    Odrv12 I__2188 (
            .O(N__9757),
            .I(DRA_c_0));
    InMux I__2187 (
            .O(N__9754),
            .I(N__9751));
    LocalMux I__2186 (
            .O(N__9751),
            .I(N__9748));
    Span4Mux_v I__2185 (
            .O(N__9748),
            .I(N__9745));
    Span4Mux_h I__2184 (
            .O(N__9745),
            .I(N__9742));
    Odrv4 I__2183 (
            .O(N__9742),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    CascadeMux I__2182 (
            .O(N__9739),
            .I(N_334_cascade_));
    IoInMux I__2181 (
            .O(N__9736),
            .I(N__9733));
    LocalMux I__2180 (
            .O(N__9733),
            .I(N__9730));
    Span4Mux_s3_h I__2179 (
            .O(N__9730),
            .I(N__9727));
    Sp12to4 I__2178 (
            .O(N__9727),
            .I(N__9724));
    Span12Mux_s8_v I__2177 (
            .O(N__9724),
            .I(N__9721));
    Span12Mux_h I__2176 (
            .O(N__9721),
            .I(N__9718));
    Odrv12 I__2175 (
            .O(N__9718),
            .I(N_177_i));
    InMux I__2174 (
            .O(N__9715),
            .I(N__9711));
    InMux I__2173 (
            .O(N__9714),
            .I(N__9708));
    LocalMux I__2172 (
            .O(N__9711),
            .I(N__9704));
    LocalMux I__2171 (
            .O(N__9708),
            .I(N__9701));
    InMux I__2170 (
            .O(N__9707),
            .I(N__9698));
    Span4Mux_v I__2169 (
            .O(N__9704),
            .I(N__9690));
    Span4Mux_h I__2168 (
            .O(N__9701),
            .I(N__9690));
    LocalMux I__2167 (
            .O(N__9698),
            .I(N__9690));
    InMux I__2166 (
            .O(N__9697),
            .I(N__9687));
    Span4Mux_v I__2165 (
            .O(N__9690),
            .I(N__9684));
    LocalMux I__2164 (
            .O(N__9687),
            .I(N__9681));
    Span4Mux_v I__2163 (
            .O(N__9684),
            .I(N__9678));
    Span12Mux_v I__2162 (
            .O(N__9681),
            .I(N__9673));
    Sp12to4 I__2161 (
            .O(N__9678),
            .I(N__9673));
    Span12Mux_h I__2160 (
            .O(N__9673),
            .I(N__9670));
    Odrv12 I__2159 (
            .O(N__9670),
            .I(DRA_c_2));
    InMux I__2158 (
            .O(N__9667),
            .I(N__9664));
    LocalMux I__2157 (
            .O(N__9664),
            .I(N__9661));
    Odrv4 I__2156 (
            .O(N__9661),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__2155 (
            .O(N__9658),
            .I(N__9655));
    LocalMux I__2154 (
            .O(N__9655),
            .I(N__9652));
    Odrv4 I__2153 (
            .O(N__9652),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__2152 (
            .O(N__9649),
            .I(N__9646));
    LocalMux I__2151 (
            .O(N__9646),
            .I(N__9642));
    InMux I__2150 (
            .O(N__9645),
            .I(N__9639));
    Span4Mux_v I__2149 (
            .O(N__9642),
            .I(N__9634));
    LocalMux I__2148 (
            .O(N__9639),
            .I(N__9631));
    InMux I__2147 (
            .O(N__9638),
            .I(N__9628));
    InMux I__2146 (
            .O(N__9637),
            .I(N__9625));
    Span4Mux_v I__2145 (
            .O(N__9634),
            .I(N__9622));
    Sp12to4 I__2144 (
            .O(N__9631),
            .I(N__9615));
    LocalMux I__2143 (
            .O(N__9628),
            .I(N__9615));
    LocalMux I__2142 (
            .O(N__9625),
            .I(N__9615));
    Sp12to4 I__2141 (
            .O(N__9622),
            .I(N__9610));
    Span12Mux_v I__2140 (
            .O(N__9615),
            .I(N__9610));
    Span12Mux_h I__2139 (
            .O(N__9610),
            .I(N__9607));
    Odrv12 I__2138 (
            .O(N__9607),
            .I(DRA_c_5));
    InMux I__2137 (
            .O(N__9604),
            .I(N__9601));
    LocalMux I__2136 (
            .O(N__9601),
            .I(N__9598));
    Span12Mux_v I__2135 (
            .O(N__9598),
            .I(N__9595));
    Odrv12 I__2134 (
            .O(N__9595),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    IoInMux I__2133 (
            .O(N__9592),
            .I(N__9589));
    LocalMux I__2132 (
            .O(N__9589),
            .I(N__9586));
    Odrv12 I__2131 (
            .O(N__9586),
            .I(RESETn_c_i));
    InMux I__2130 (
            .O(N__9583),
            .I(N__9580));
    LocalMux I__2129 (
            .O(N__9580),
            .I(N__9576));
    InMux I__2128 (
            .O(N__9579),
            .I(N__9573));
    Span4Mux_h I__2127 (
            .O(N__9576),
            .I(N__9567));
    LocalMux I__2126 (
            .O(N__9573),
            .I(N__9567));
    CascadeMux I__2125 (
            .O(N__9572),
            .I(N__9562));
    Span4Mux_h I__2124 (
            .O(N__9567),
            .I(N__9559));
    InMux I__2123 (
            .O(N__9566),
            .I(N__9556));
    InMux I__2122 (
            .O(N__9565),
            .I(N__9553));
    InMux I__2121 (
            .O(N__9562),
            .I(N__9550));
    Odrv4 I__2120 (
            .O(N__9559),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__2119 (
            .O(N__9556),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__2118 (
            .O(N__9553),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__2117 (
            .O(N__9550),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__2116 (
            .O(N__9541),
            .I(N__9538));
    LocalMux I__2115 (
            .O(N__9538),
            .I(N__9535));
    Span4Mux_s2_v I__2114 (
            .O(N__9535),
            .I(N__9532));
    Span4Mux_v I__2113 (
            .O(N__9532),
            .I(N__9529));
    Span4Mux_v I__2112 (
            .O(N__9529),
            .I(N__9526));
    Span4Mux_h I__2111 (
            .O(N__9526),
            .I(N__9523));
    Odrv4 I__2110 (
            .O(N__9523),
            .I(CRCSn_c));
    InMux I__2109 (
            .O(N__9520),
            .I(N__9517));
    LocalMux I__2108 (
            .O(N__9517),
            .I(N__9514));
    Odrv12 I__2107 (
            .O(N__9514),
            .I(\U712_CHIP_RAM.CMA_5_i_0_9 ));
    InMux I__2106 (
            .O(N__9511),
            .I(N__9508));
    LocalMux I__2105 (
            .O(N__9508),
            .I(N__9505));
    Span4Mux_v I__2104 (
            .O(N__9505),
            .I(N__9502));
    Span4Mux_v I__2103 (
            .O(N__9502),
            .I(N__9499));
    Sp12to4 I__2102 (
            .O(N__9499),
            .I(N__9496));
    Span12Mux_h I__2101 (
            .O(N__9496),
            .I(N__9493));
    Odrv12 I__2100 (
            .O(N__9493),
            .I(A_c_19));
    InMux I__2099 (
            .O(N__9490),
            .I(N__9487));
    LocalMux I__2098 (
            .O(N__9487),
            .I(N__9484));
    Odrv4 I__2097 (
            .O(N__9484),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    IoInMux I__2096 (
            .O(N__9481),
            .I(N__9478));
    LocalMux I__2095 (
            .O(N__9478),
            .I(N__9475));
    Span4Mux_s3_h I__2094 (
            .O(N__9475),
            .I(N__9472));
    Sp12to4 I__2093 (
            .O(N__9472),
            .I(N__9469));
    Span12Mux_s10_v I__2092 (
            .O(N__9469),
            .I(N__9466));
    Span12Mux_h I__2091 (
            .O(N__9466),
            .I(N__9463));
    Odrv12 I__2090 (
            .O(N__9463),
            .I(CMA_c_9));
    CEMux I__2089 (
            .O(N__9460),
            .I(N__9455));
    CEMux I__2088 (
            .O(N__9459),
            .I(N__9452));
    CEMux I__2087 (
            .O(N__9458),
            .I(N__9448));
    LocalMux I__2086 (
            .O(N__9455),
            .I(N__9445));
    LocalMux I__2085 (
            .O(N__9452),
            .I(N__9441));
    CEMux I__2084 (
            .O(N__9451),
            .I(N__9438));
    LocalMux I__2083 (
            .O(N__9448),
            .I(N__9435));
    Span4Mux_v I__2082 (
            .O(N__9445),
            .I(N__9432));
    CEMux I__2081 (
            .O(N__9444),
            .I(N__9429));
    Span4Mux_h I__2080 (
            .O(N__9441),
            .I(N__9424));
    LocalMux I__2079 (
            .O(N__9438),
            .I(N__9424));
    Span4Mux_h I__2078 (
            .O(N__9435),
            .I(N__9421));
    Span4Mux_h I__2077 (
            .O(N__9432),
            .I(N__9418));
    LocalMux I__2076 (
            .O(N__9429),
            .I(N__9415));
    Sp12to4 I__2075 (
            .O(N__9424),
            .I(N__9412));
    Odrv4 I__2074 (
            .O(N__9421),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv4 I__2073 (
            .O(N__9418),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv4 I__2072 (
            .O(N__9415),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv12 I__2071 (
            .O(N__9412),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    CascadeMux I__2070 (
            .O(N__9403),
            .I(N__9400));
    InMux I__2069 (
            .O(N__9400),
            .I(N__9397));
    LocalMux I__2068 (
            .O(N__9397),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2067 (
            .O(N__9394),
            .I(N__9391));
    LocalMux I__2066 (
            .O(N__9391),
            .I(N__9388));
    Span4Mux_h I__2065 (
            .O(N__9388),
            .I(N__9385));
    Odrv4 I__2064 (
            .O(N__9385),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__2063 (
            .O(N__9382),
            .I(N__9379));
    LocalMux I__2062 (
            .O(N__9379),
            .I(N__9376));
    Span4Mux_v I__2061 (
            .O(N__9376),
            .I(N__9373));
    Odrv4 I__2060 (
            .O(N__9373),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2059 (
            .O(N__9370),
            .I(N__9367));
    LocalMux I__2058 (
            .O(N__9367),
            .I(N__9364));
    Span4Mux_h I__2057 (
            .O(N__9364),
            .I(N__9361));
    Odrv4 I__2056 (
            .O(N__9361),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__2055 (
            .O(N__9358),
            .I(N__9355));
    LocalMux I__2054 (
            .O(N__9355),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__2053 (
            .O(N__9352),
            .I(N__9349));
    LocalMux I__2052 (
            .O(N__9349),
            .I(N__9346));
    Odrv4 I__2051 (
            .O(N__9346),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2050 (
            .O(N__9343),
            .I(N__9340));
    LocalMux I__2049 (
            .O(N__9340),
            .I(N__9337));
    Odrv4 I__2048 (
            .O(N__9337),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__2047 (
            .O(N__9334),
            .I(N__9326));
    InMux I__2046 (
            .O(N__9333),
            .I(N__9326));
    InMux I__2045 (
            .O(N__9332),
            .I(N__9323));
    InMux I__2044 (
            .O(N__9331),
            .I(N__9320));
    LocalMux I__2043 (
            .O(N__9326),
            .I(N__9317));
    LocalMux I__2042 (
            .O(N__9323),
            .I(N__9312));
    LocalMux I__2041 (
            .O(N__9320),
            .I(N__9312));
    Span4Mux_v I__2040 (
            .O(N__9317),
            .I(N__9309));
    Span4Mux_h I__2039 (
            .O(N__9312),
            .I(N__9306));
    Span4Mux_h I__2038 (
            .O(N__9309),
            .I(N__9303));
    Span4Mux_h I__2037 (
            .O(N__9306),
            .I(N__9300));
    Sp12to4 I__2036 (
            .O(N__9303),
            .I(N__9295));
    Sp12to4 I__2035 (
            .O(N__9300),
            .I(N__9295));
    Odrv12 I__2034 (
            .O(N__9295),
            .I(DRA_c_8));
    InMux I__2033 (
            .O(N__9292),
            .I(N__9289));
    LocalMux I__2032 (
            .O(N__9289),
            .I(N__9286));
    Span4Mux_h I__2031 (
            .O(N__9286),
            .I(N__9283));
    Odrv4 I__2030 (
            .O(N__9283),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2029 (
            .O(N__9280),
            .I(N__9277));
    LocalMux I__2028 (
            .O(N__9277),
            .I(N__9274));
    Odrv12 I__2027 (
            .O(N__9274),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__2026 (
            .O(N__9271),
            .I(N__9265));
    InMux I__2025 (
            .O(N__9270),
            .I(N__9265));
    LocalMux I__2024 (
            .O(N__9265),
            .I(N__9262));
    Span4Mux_v I__2023 (
            .O(N__9262),
            .I(N__9259));
    Odrv4 I__2022 (
            .O(N__9259),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2021 (
            .O(N__9256),
            .I(N__9252));
    CascadeMux I__2020 (
            .O(N__9255),
            .I(N__9249));
    LocalMux I__2019 (
            .O(N__9252),
            .I(N__9246));
    InMux I__2018 (
            .O(N__9249),
            .I(N__9243));
    Odrv12 I__2017 (
            .O(N__9246),
            .I(\U712_CHIP_RAM.m50_i_a2_0_0 ));
    LocalMux I__2016 (
            .O(N__9243),
            .I(\U712_CHIP_RAM.m50_i_a2_0_0 ));
    IoInMux I__2015 (
            .O(N__9238),
            .I(N__9235));
    LocalMux I__2014 (
            .O(N__9235),
            .I(N__9232));
    Span12Mux_s4_h I__2013 (
            .O(N__9232),
            .I(N__9229));
    Span12Mux_v I__2012 (
            .O(N__9229),
            .I(N__9226));
    Span12Mux_h I__2011 (
            .O(N__9226),
            .I(N__9223));
    Odrv12 I__2010 (
            .O(N__9223),
            .I(N_200_i));
    InMux I__2009 (
            .O(N__9220),
            .I(N__9217));
    LocalMux I__2008 (
            .O(N__9217),
            .I(N__9214));
    Odrv4 I__2007 (
            .O(N__9214),
            .I(\U712_CHIP_RAM.N_337 ));
    CascadeMux I__2006 (
            .O(N__9211),
            .I(N__9205));
    InMux I__2005 (
            .O(N__9210),
            .I(N__9202));
    InMux I__2004 (
            .O(N__9209),
            .I(N__9199));
    InMux I__2003 (
            .O(N__9208),
            .I(N__9196));
    InMux I__2002 (
            .O(N__9205),
            .I(N__9193));
    LocalMux I__2001 (
            .O(N__9202),
            .I(N__9190));
    LocalMux I__2000 (
            .O(N__9199),
            .I(N__9185));
    LocalMux I__1999 (
            .O(N__9196),
            .I(N__9185));
    LocalMux I__1998 (
            .O(N__9193),
            .I(N__9182));
    Span4Mux_v I__1997 (
            .O(N__9190),
            .I(N__9179));
    Span4Mux_v I__1996 (
            .O(N__9185),
            .I(N__9176));
    Span4Mux_v I__1995 (
            .O(N__9182),
            .I(N__9173));
    Span4Mux_h I__1994 (
            .O(N__9179),
            .I(N__9170));
    Sp12to4 I__1993 (
            .O(N__9176),
            .I(N__9167));
    Sp12to4 I__1992 (
            .O(N__9173),
            .I(N__9164));
    Sp12to4 I__1991 (
            .O(N__9170),
            .I(N__9157));
    Span12Mux_h I__1990 (
            .O(N__9167),
            .I(N__9157));
    Span12Mux_h I__1989 (
            .O(N__9164),
            .I(N__9157));
    Span12Mux_v I__1988 (
            .O(N__9157),
            .I(N__9154));
    Odrv12 I__1987 (
            .O(N__9154),
            .I(CLK40_PLL_i));
    IoInMux I__1986 (
            .O(N__9151),
            .I(N__9148));
    LocalMux I__1985 (
            .O(N__9148),
            .I(N__9143));
    IoInMux I__1984 (
            .O(N__9147),
            .I(N__9140));
    IoInMux I__1983 (
            .O(N__9146),
            .I(N__9137));
    IoSpan4Mux I__1982 (
            .O(N__9143),
            .I(N__9132));
    LocalMux I__1981 (
            .O(N__9140),
            .I(N__9132));
    LocalMux I__1980 (
            .O(N__9137),
            .I(N__9129));
    IoSpan4Mux I__1979 (
            .O(N__9132),
            .I(N__9126));
    Span4Mux_s2_h I__1978 (
            .O(N__9129),
            .I(N__9123));
    Span4Mux_s0_v I__1977 (
            .O(N__9126),
            .I(N__9120));
    Span4Mux_v I__1976 (
            .O(N__9123),
            .I(N__9117));
    Sp12to4 I__1975 (
            .O(N__9120),
            .I(N__9114));
    Sp12to4 I__1974 (
            .O(N__9117),
            .I(N__9111));
    Span12Mux_v I__1973 (
            .O(N__9114),
            .I(N__9106));
    Span12Mux_h I__1972 (
            .O(N__9111),
            .I(N__9106));
    Odrv12 I__1971 (
            .O(N__9106),
            .I(CLK40_PLL_i_i));
    InMux I__1970 (
            .O(N__9103),
            .I(N__9100));
    LocalMux I__1969 (
            .O(N__9100),
            .I(N__9097));
    Odrv4 I__1968 (
            .O(N__9097),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ));
    IoInMux I__1967 (
            .O(N__9094),
            .I(N__9091));
    LocalMux I__1966 (
            .O(N__9091),
            .I(N__9088));
    IoSpan4Mux I__1965 (
            .O(N__9088),
            .I(N__9085));
    Span4Mux_s3_h I__1964 (
            .O(N__9085),
            .I(N__9082));
    Span4Mux_v I__1963 (
            .O(N__9082),
            .I(N__9079));
    Span4Mux_h I__1962 (
            .O(N__9079),
            .I(N__9076));
    Sp12to4 I__1961 (
            .O(N__9076),
            .I(N__9073));
    Odrv12 I__1960 (
            .O(N__9073),
            .I(CMA_c_8));
    IoInMux I__1959 (
            .O(N__9070),
            .I(N__9067));
    LocalMux I__1958 (
            .O(N__9067),
            .I(N__9064));
    Span4Mux_s0_v I__1957 (
            .O(N__9064),
            .I(N__9061));
    Sp12to4 I__1956 (
            .O(N__9061),
            .I(N__9058));
    Span12Mux_h I__1955 (
            .O(N__9058),
            .I(N__9055));
    Odrv12 I__1954 (
            .O(N__9055),
            .I(CMA_c_0));
    InMux I__1953 (
            .O(N__9052),
            .I(N__9049));
    LocalMux I__1952 (
            .O(N__9049),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1951 (
            .O(N__9046),
            .I(N__9043));
    LocalMux I__1950 (
            .O(N__9043),
            .I(N__9040));
    IoSpan4Mux I__1949 (
            .O(N__9040),
            .I(N__9037));
    Span4Mux_s2_h I__1948 (
            .O(N__9037),
            .I(N__9034));
    Sp12to4 I__1947 (
            .O(N__9034),
            .I(N__9031));
    Span12Mux_h I__1946 (
            .O(N__9031),
            .I(N__9028));
    Odrv12 I__1945 (
            .O(N__9028),
            .I(CMA_c_7));
    IoInMux I__1944 (
            .O(N__9025),
            .I(N__9022));
    LocalMux I__1943 (
            .O(N__9022),
            .I(N__9018));
    InMux I__1942 (
            .O(N__9021),
            .I(N__9015));
    Span12Mux_s4_v I__1941 (
            .O(N__9018),
            .I(N__9012));
    LocalMux I__1940 (
            .O(N__9015),
            .I(N__9009));
    Span12Mux_v I__1939 (
            .O(N__9012),
            .I(N__9004));
    Span12Mux_v I__1938 (
            .O(N__9009),
            .I(N__9004));
    Span12Mux_h I__1937 (
            .O(N__9004),
            .I(N__9001));
    Odrv12 I__1936 (
            .O(N__9001),
            .I(A_c_9));
    InMux I__1935 (
            .O(N__8998),
            .I(N__8995));
    LocalMux I__1934 (
            .O(N__8995),
            .I(N__8992));
    Odrv12 I__1933 (
            .O(N__8992),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ));
    CascadeMux I__1932 (
            .O(N__8989),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ));
    InMux I__1931 (
            .O(N__8986),
            .I(N__8983));
    LocalMux I__1930 (
            .O(N__8983),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    InMux I__1929 (
            .O(N__8980),
            .I(N__8977));
    LocalMux I__1928 (
            .O(N__8977),
            .I(N__8974));
    Odrv4 I__1927 (
            .O(N__8974),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    CascadeMux I__1926 (
            .O(N__8971),
            .I(N__8967));
    InMux I__1925 (
            .O(N__8970),
            .I(N__8953));
    InMux I__1924 (
            .O(N__8967),
            .I(N__8953));
    CascadeMux I__1923 (
            .O(N__8966),
            .I(N__8946));
    CascadeMux I__1922 (
            .O(N__8965),
            .I(N__8943));
    CascadeMux I__1921 (
            .O(N__8964),
            .I(N__8939));
    InMux I__1920 (
            .O(N__8963),
            .I(N__8933));
    InMux I__1919 (
            .O(N__8962),
            .I(N__8933));
    InMux I__1918 (
            .O(N__8961),
            .I(N__8926));
    InMux I__1917 (
            .O(N__8960),
            .I(N__8926));
    InMux I__1916 (
            .O(N__8959),
            .I(N__8926));
    InMux I__1915 (
            .O(N__8958),
            .I(N__8923));
    LocalMux I__1914 (
            .O(N__8953),
            .I(N__8920));
    InMux I__1913 (
            .O(N__8952),
            .I(N__8913));
    InMux I__1912 (
            .O(N__8951),
            .I(N__8913));
    InMux I__1911 (
            .O(N__8950),
            .I(N__8913));
    InMux I__1910 (
            .O(N__8949),
            .I(N__8910));
    InMux I__1909 (
            .O(N__8946),
            .I(N__8907));
    InMux I__1908 (
            .O(N__8943),
            .I(N__8902));
    InMux I__1907 (
            .O(N__8942),
            .I(N__8902));
    InMux I__1906 (
            .O(N__8939),
            .I(N__8897));
    InMux I__1905 (
            .O(N__8938),
            .I(N__8897));
    LocalMux I__1904 (
            .O(N__8933),
            .I(N__8892));
    LocalMux I__1903 (
            .O(N__8926),
            .I(N__8892));
    LocalMux I__1902 (
            .O(N__8923),
            .I(N__8885));
    Span4Mux_v I__1901 (
            .O(N__8920),
            .I(N__8880));
    LocalMux I__1900 (
            .O(N__8913),
            .I(N__8880));
    LocalMux I__1899 (
            .O(N__8910),
            .I(N__8875));
    LocalMux I__1898 (
            .O(N__8907),
            .I(N__8875));
    LocalMux I__1897 (
            .O(N__8902),
            .I(N__8870));
    LocalMux I__1896 (
            .O(N__8897),
            .I(N__8870));
    Span4Mux_v I__1895 (
            .O(N__8892),
            .I(N__8867));
    InMux I__1894 (
            .O(N__8891),
            .I(N__8860));
    InMux I__1893 (
            .O(N__8890),
            .I(N__8860));
    InMux I__1892 (
            .O(N__8889),
            .I(N__8860));
    InMux I__1891 (
            .O(N__8888),
            .I(N__8853));
    Span4Mux_h I__1890 (
            .O(N__8885),
            .I(N__8848));
    Span4Mux_h I__1889 (
            .O(N__8880),
            .I(N__8848));
    Span4Mux_v I__1888 (
            .O(N__8875),
            .I(N__8839));
    Span4Mux_h I__1887 (
            .O(N__8870),
            .I(N__8839));
    Span4Mux_h I__1886 (
            .O(N__8867),
            .I(N__8839));
    LocalMux I__1885 (
            .O(N__8860),
            .I(N__8839));
    InMux I__1884 (
            .O(N__8859),
            .I(N__8830));
    InMux I__1883 (
            .O(N__8858),
            .I(N__8830));
    InMux I__1882 (
            .O(N__8857),
            .I(N__8830));
    InMux I__1881 (
            .O(N__8856),
            .I(N__8830));
    LocalMux I__1880 (
            .O(N__8853),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1879 (
            .O(N__8848),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1878 (
            .O(N__8839),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1877 (
            .O(N__8830),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    InMux I__1876 (
            .O(N__8821),
            .I(N__8812));
    InMux I__1875 (
            .O(N__8820),
            .I(N__8809));
    InMux I__1874 (
            .O(N__8819),
            .I(N__8802));
    InMux I__1873 (
            .O(N__8818),
            .I(N__8802));
    InMux I__1872 (
            .O(N__8817),
            .I(N__8802));
    InMux I__1871 (
            .O(N__8816),
            .I(N__8797));
    InMux I__1870 (
            .O(N__8815),
            .I(N__8797));
    LocalMux I__1869 (
            .O(N__8812),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ));
    LocalMux I__1868 (
            .O(N__8809),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ));
    LocalMux I__1867 (
            .O(N__8802),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ));
    LocalMux I__1866 (
            .O(N__8797),
            .I(\U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ));
    CascadeMux I__1865 (
            .O(N__8788),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_ ));
    CascadeMux I__1864 (
            .O(N__8785),
            .I(N__8778));
    CascadeMux I__1863 (
            .O(N__8784),
            .I(N__8775));
    CascadeMux I__1862 (
            .O(N__8783),
            .I(N__8772));
    CascadeMux I__1861 (
            .O(N__8782),
            .I(N__8767));
    CascadeMux I__1860 (
            .O(N__8781),
            .I(N__8764));
    InMux I__1859 (
            .O(N__8778),
            .I(N__8761));
    InMux I__1858 (
            .O(N__8775),
            .I(N__8756));
    InMux I__1857 (
            .O(N__8772),
            .I(N__8756));
    CascadeMux I__1856 (
            .O(N__8771),
            .I(N__8753));
    InMux I__1855 (
            .O(N__8770),
            .I(N__8748));
    InMux I__1854 (
            .O(N__8767),
            .I(N__8743));
    InMux I__1853 (
            .O(N__8764),
            .I(N__8743));
    LocalMux I__1852 (
            .O(N__8761),
            .I(N__8738));
    LocalMux I__1851 (
            .O(N__8756),
            .I(N__8738));
    InMux I__1850 (
            .O(N__8753),
            .I(N__8734));
    InMux I__1849 (
            .O(N__8752),
            .I(N__8731));
    InMux I__1848 (
            .O(N__8751),
            .I(N__8728));
    LocalMux I__1847 (
            .O(N__8748),
            .I(N__8723));
    LocalMux I__1846 (
            .O(N__8743),
            .I(N__8723));
    Span4Mux_v I__1845 (
            .O(N__8738),
            .I(N__8720));
    InMux I__1844 (
            .O(N__8737),
            .I(N__8717));
    LocalMux I__1843 (
            .O(N__8734),
            .I(\U712_CHIP_RAM.N_314 ));
    LocalMux I__1842 (
            .O(N__8731),
            .I(\U712_CHIP_RAM.N_314 ));
    LocalMux I__1841 (
            .O(N__8728),
            .I(\U712_CHIP_RAM.N_314 ));
    Odrv4 I__1840 (
            .O(N__8723),
            .I(\U712_CHIP_RAM.N_314 ));
    Odrv4 I__1839 (
            .O(N__8720),
            .I(\U712_CHIP_RAM.N_314 ));
    LocalMux I__1838 (
            .O(N__8717),
            .I(\U712_CHIP_RAM.N_314 ));
    IoInMux I__1837 (
            .O(N__8704),
            .I(N__8701));
    LocalMux I__1836 (
            .O(N__8701),
            .I(N__8698));
    Span12Mux_s0_v I__1835 (
            .O(N__8698),
            .I(N__8695));
    Span12Mux_v I__1834 (
            .O(N__8695),
            .I(N__8692));
    Odrv12 I__1833 (
            .O(N__8692),
            .I(CMA_c_2));
    InMux I__1832 (
            .O(N__8689),
            .I(N__8686));
    LocalMux I__1831 (
            .O(N__8686),
            .I(N__8683));
    Odrv4 I__1830 (
            .O(N__8683),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1829 (
            .O(N__8680),
            .I(N__8674));
    InMux I__1828 (
            .O(N__8679),
            .I(N__8674));
    LocalMux I__1827 (
            .O(N__8674),
            .I(N__8669));
    InMux I__1826 (
            .O(N__8673),
            .I(N__8666));
    InMux I__1825 (
            .O(N__8672),
            .I(N__8663));
    Span4Mux_h I__1824 (
            .O(N__8669),
            .I(N__8658));
    LocalMux I__1823 (
            .O(N__8666),
            .I(N__8658));
    LocalMux I__1822 (
            .O(N__8663),
            .I(N__8655));
    Span4Mux_v I__1821 (
            .O(N__8658),
            .I(N__8652));
    Span4Mux_h I__1820 (
            .O(N__8655),
            .I(N__8649));
    Sp12to4 I__1819 (
            .O(N__8652),
            .I(N__8646));
    Sp12to4 I__1818 (
            .O(N__8649),
            .I(N__8643));
    Span12Mux_h I__1817 (
            .O(N__8646),
            .I(N__8640));
    Span12Mux_v I__1816 (
            .O(N__8643),
            .I(N__8637));
    Span12Mux_v I__1815 (
            .O(N__8640),
            .I(N__8634));
    Span12Mux_h I__1814 (
            .O(N__8637),
            .I(N__8631));
    Odrv12 I__1813 (
            .O(N__8634),
            .I(DRA_c_9));
    Odrv12 I__1812 (
            .O(N__8631),
            .I(DRA_c_9));
    InMux I__1811 (
            .O(N__8626),
            .I(N__8617));
    InMux I__1810 (
            .O(N__8625),
            .I(N__8617));
    InMux I__1809 (
            .O(N__8624),
            .I(N__8617));
    LocalMux I__1808 (
            .O(N__8617),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__1807 (
            .O(N__8614),
            .I(\U712_CYCLE_TERM.N_455_cascade_ ));
    InMux I__1806 (
            .O(N__8611),
            .I(N__8606));
    InMux I__1805 (
            .O(N__8610),
            .I(N__8602));
    CascadeMux I__1804 (
            .O(N__8609),
            .I(N__8599));
    LocalMux I__1803 (
            .O(N__8606),
            .I(N__8596));
    InMux I__1802 (
            .O(N__8605),
            .I(N__8593));
    LocalMux I__1801 (
            .O(N__8602),
            .I(N__8590));
    InMux I__1800 (
            .O(N__8599),
            .I(N__8587));
    Span4Mux_h I__1799 (
            .O(N__8596),
            .I(N__8580));
    LocalMux I__1798 (
            .O(N__8593),
            .I(N__8580));
    Span4Mux_v I__1797 (
            .O(N__8590),
            .I(N__8580));
    LocalMux I__1796 (
            .O(N__8587),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    Odrv4 I__1795 (
            .O(N__8580),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__1794 (
            .O(N__8575),
            .I(N__8569));
    InMux I__1793 (
            .O(N__8574),
            .I(N__8562));
    InMux I__1792 (
            .O(N__8573),
            .I(N__8562));
    InMux I__1791 (
            .O(N__8572),
            .I(N__8562));
    LocalMux I__1790 (
            .O(N__8569),
            .I(REG_TACK));
    LocalMux I__1789 (
            .O(N__8562),
            .I(REG_TACK));
    CascadeMux I__1788 (
            .O(N__8557),
            .I(N__8554));
    InMux I__1787 (
            .O(N__8554),
            .I(N__8548));
    InMux I__1786 (
            .O(N__8553),
            .I(N__8543));
    InMux I__1785 (
            .O(N__8552),
            .I(N__8543));
    InMux I__1784 (
            .O(N__8551),
            .I(N__8540));
    LocalMux I__1783 (
            .O(N__8548),
            .I(N__8535));
    LocalMux I__1782 (
            .O(N__8543),
            .I(N__8535));
    LocalMux I__1781 (
            .O(N__8540),
            .I(CPU_TACKm));
    Odrv12 I__1780 (
            .O(N__8535),
            .I(CPU_TACKm));
    InMux I__1779 (
            .O(N__8530),
            .I(N__8527));
    LocalMux I__1778 (
            .O(N__8527),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__1777 (
            .O(N__8524),
            .I(N__8519));
    InMux I__1776 (
            .O(N__8523),
            .I(N__8516));
    InMux I__1775 (
            .O(N__8522),
            .I(N__8513));
    InMux I__1774 (
            .O(N__8519),
            .I(N__8510));
    LocalMux I__1773 (
            .O(N__8516),
            .I(N__8507));
    LocalMux I__1772 (
            .O(N__8513),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    LocalMux I__1771 (
            .O(N__8510),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    Odrv12 I__1770 (
            .O(N__8507),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    InMux I__1769 (
            .O(N__8500),
            .I(N__8497));
    LocalMux I__1768 (
            .O(N__8497),
            .I(N__8489));
    InMux I__1767 (
            .O(N__8496),
            .I(N__8486));
    InMux I__1766 (
            .O(N__8495),
            .I(N__8483));
    InMux I__1765 (
            .O(N__8494),
            .I(N__8476));
    InMux I__1764 (
            .O(N__8493),
            .I(N__8476));
    InMux I__1763 (
            .O(N__8492),
            .I(N__8476));
    Odrv4 I__1762 (
            .O(N__8489),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__1761 (
            .O(N__8486),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__1760 (
            .O(N__8483),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    LocalMux I__1759 (
            .O(N__8476),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    InMux I__1758 (
            .O(N__8467),
            .I(N__8464));
    LocalMux I__1757 (
            .O(N__8464),
            .I(N__8460));
    InMux I__1756 (
            .O(N__8463),
            .I(N__8457));
    Odrv4 I__1755 (
            .O(N__8460),
            .I(\U712_REG_SM.START_RSTZ0 ));
    LocalMux I__1754 (
            .O(N__8457),
            .I(\U712_REG_SM.START_RSTZ0 ));
    IoInMux I__1753 (
            .O(N__8452),
            .I(N__8449));
    LocalMux I__1752 (
            .O(N__8449),
            .I(N__8446));
    Span12Mux_s9_v I__1751 (
            .O(N__8446),
            .I(N__8443));
    Span12Mux_h I__1750 (
            .O(N__8443),
            .I(N__8440));
    Odrv12 I__1749 (
            .O(N__8440),
            .I(CASn_c));
    InMux I__1748 (
            .O(N__8437),
            .I(N__8434));
    LocalMux I__1747 (
            .O(N__8434),
            .I(\U712_CHIP_RAM.N_361 ));
    InMux I__1746 (
            .O(N__8431),
            .I(N__8428));
    LocalMux I__1745 (
            .O(N__8428),
            .I(\U712_CHIP_RAM.N_367 ));
    IoInMux I__1744 (
            .O(N__8425),
            .I(N__8422));
    LocalMux I__1743 (
            .O(N__8422),
            .I(N__8419));
    IoSpan4Mux I__1742 (
            .O(N__8419),
            .I(N__8416));
    Span4Mux_s2_h I__1741 (
            .O(N__8416),
            .I(N__8413));
    Sp12to4 I__1740 (
            .O(N__8413),
            .I(N__8410));
    Span12Mux_h I__1739 (
            .O(N__8410),
            .I(N__8407));
    Odrv12 I__1738 (
            .O(N__8407),
            .I(CMA_c_5));
    IoInMux I__1737 (
            .O(N__8404),
            .I(N__8401));
    LocalMux I__1736 (
            .O(N__8401),
            .I(N__8398));
    IoSpan4Mux I__1735 (
            .O(N__8398),
            .I(N__8395));
    Span4Mux_s3_v I__1734 (
            .O(N__8395),
            .I(N__8392));
    Span4Mux_v I__1733 (
            .O(N__8392),
            .I(N__8389));
    Span4Mux_h I__1732 (
            .O(N__8389),
            .I(N__8386));
    Odrv4 I__1731 (
            .O(N__8386),
            .I(CMA_c_10));
    InMux I__1730 (
            .O(N__8383),
            .I(N__8380));
    LocalMux I__1729 (
            .O(N__8380),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    InMux I__1728 (
            .O(N__8377),
            .I(N__8374));
    LocalMux I__1727 (
            .O(N__8374),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    InMux I__1726 (
            .O(N__8371),
            .I(N__8368));
    LocalMux I__1725 (
            .O(N__8368),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    IoInMux I__1724 (
            .O(N__8365),
            .I(N__8362));
    LocalMux I__1723 (
            .O(N__8362),
            .I(N__8359));
    Span12Mux_s5_v I__1722 (
            .O(N__8359),
            .I(N__8356));
    Odrv12 I__1721 (
            .O(N__8356),
            .I(CMA_c_1));
    IoInMux I__1720 (
            .O(N__8353),
            .I(N__8350));
    LocalMux I__1719 (
            .O(N__8350),
            .I(N__8347));
    IoSpan4Mux I__1718 (
            .O(N__8347),
            .I(N__8344));
    Span4Mux_s2_h I__1717 (
            .O(N__8344),
            .I(N__8341));
    Sp12to4 I__1716 (
            .O(N__8341),
            .I(N__8338));
    Span12Mux_s9_h I__1715 (
            .O(N__8338),
            .I(N__8335));
    Span12Mux_v I__1714 (
            .O(N__8335),
            .I(N__8332));
    Odrv12 I__1713 (
            .O(N__8332),
            .I(CMA_c_3));
    IoInMux I__1712 (
            .O(N__8329),
            .I(N__8326));
    LocalMux I__1711 (
            .O(N__8326),
            .I(N__8323));
    IoSpan4Mux I__1710 (
            .O(N__8323),
            .I(N__8320));
    Span4Mux_s3_h I__1709 (
            .O(N__8320),
            .I(N__8317));
    Sp12to4 I__1708 (
            .O(N__8317),
            .I(N__8314));
    Span12Mux_h I__1707 (
            .O(N__8314),
            .I(N__8311));
    Odrv12 I__1706 (
            .O(N__8311),
            .I(CMA_c_4));
    InMux I__1705 (
            .O(N__8308),
            .I(N__8305));
    LocalMux I__1704 (
            .O(N__8305),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__1703 (
            .O(N__8302),
            .I(N__8299));
    LocalMux I__1702 (
            .O(N__8299),
            .I(N__8296));
    IoSpan4Mux I__1701 (
            .O(N__8296),
            .I(N__8293));
    Span4Mux_s2_h I__1700 (
            .O(N__8293),
            .I(N__8290));
    Sp12to4 I__1699 (
            .O(N__8290),
            .I(N__8287));
    Span12Mux_s11_h I__1698 (
            .O(N__8287),
            .I(N__8284));
    Span12Mux_v I__1697 (
            .O(N__8284),
            .I(N__8281));
    Odrv12 I__1696 (
            .O(N__8281),
            .I(CMA_c_6));
    CascadeMux I__1695 (
            .O(N__8278),
            .I(N__8275));
    InMux I__1694 (
            .O(N__8275),
            .I(N__8272));
    LocalMux I__1693 (
            .O(N__8272),
            .I(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ));
    InMux I__1692 (
            .O(N__8269),
            .I(N__8266));
    LocalMux I__1691 (
            .O(N__8266),
            .I(\U712_CHIP_RAM.N_190 ));
    InMux I__1690 (
            .O(N__8263),
            .I(N__8260));
    LocalMux I__1689 (
            .O(N__8260),
            .I(N__8257));
    Sp12to4 I__1688 (
            .O(N__8257),
            .I(N__8254));
    Span12Mux_v I__1687 (
            .O(N__8254),
            .I(N__8251));
    Span12Mux_h I__1686 (
            .O(N__8251),
            .I(N__8248));
    Odrv12 I__1685 (
            .O(N__8248),
            .I(A_c_13));
    InMux I__1684 (
            .O(N__8245),
            .I(N__8242));
    LocalMux I__1683 (
            .O(N__8242),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ));
    CascadeMux I__1682 (
            .O(N__8239),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ));
    InMux I__1681 (
            .O(N__8236),
            .I(N__8233));
    LocalMux I__1680 (
            .O(N__8233),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    InMux I__1679 (
            .O(N__8230),
            .I(N__8227));
    LocalMux I__1678 (
            .O(N__8227),
            .I(N__8224));
    Odrv4 I__1677 (
            .O(N__8224),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    CascadeMux I__1676 (
            .O(N__8221),
            .I(N__8217));
    InMux I__1675 (
            .O(N__8220),
            .I(N__8214));
    InMux I__1674 (
            .O(N__8217),
            .I(N__8211));
    LocalMux I__1673 (
            .O(N__8214),
            .I(N__8206));
    LocalMux I__1672 (
            .O(N__8211),
            .I(N__8206));
    Odrv12 I__1671 (
            .O(N__8206),
            .I(DBRn_c_i));
    InMux I__1670 (
            .O(N__8203),
            .I(N__8200));
    LocalMux I__1669 (
            .O(N__8200),
            .I(N__8196));
    InMux I__1668 (
            .O(N__8199),
            .I(N__8193));
    Span4Mux_h I__1667 (
            .O(N__8196),
            .I(N__8190));
    LocalMux I__1666 (
            .O(N__8193),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    Odrv4 I__1665 (
            .O(N__8190),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    InMux I__1664 (
            .O(N__8185),
            .I(N__8182));
    LocalMux I__1663 (
            .O(N__8182),
            .I(\U712_CYCLE_TERM.N_332 ));
    InMux I__1662 (
            .O(N__8179),
            .I(N__8174));
    InMux I__1661 (
            .O(N__8178),
            .I(N__8171));
    CascadeMux I__1660 (
            .O(N__8177),
            .I(N__8168));
    LocalMux I__1659 (
            .O(N__8174),
            .I(N__8163));
    LocalMux I__1658 (
            .O(N__8171),
            .I(N__8163));
    InMux I__1657 (
            .O(N__8168),
            .I(N__8160));
    Span4Mux_v I__1656 (
            .O(N__8163),
            .I(N__8153));
    LocalMux I__1655 (
            .O(N__8160),
            .I(N__8153));
    InMux I__1654 (
            .O(N__8159),
            .I(N__8148));
    InMux I__1653 (
            .O(N__8158),
            .I(N__8148));
    Odrv4 I__1652 (
            .O(N__8153),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__1651 (
            .O(N__8148),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    InMux I__1650 (
            .O(N__8143),
            .I(N__8140));
    LocalMux I__1649 (
            .O(N__8140),
            .I(N__8135));
    InMux I__1648 (
            .O(N__8139),
            .I(N__8132));
    InMux I__1647 (
            .O(N__8138),
            .I(N__8127));
    Span4Mux_v I__1646 (
            .O(N__8135),
            .I(N__8122));
    LocalMux I__1645 (
            .O(N__8132),
            .I(N__8122));
    InMux I__1644 (
            .O(N__8131),
            .I(N__8117));
    InMux I__1643 (
            .O(N__8130),
            .I(N__8117));
    LocalMux I__1642 (
            .O(N__8127),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1641 (
            .O(N__8122),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1640 (
            .O(N__8117),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    CascadeMux I__1639 (
            .O(N__8110),
            .I(\U712_CHIP_RAM.N_314_cascade_ ));
    InMux I__1638 (
            .O(N__8107),
            .I(N__8104));
    LocalMux I__1637 (
            .O(N__8104),
            .I(N__8101));
    Span4Mux_v I__1636 (
            .O(N__8101),
            .I(N__8098));
    Span4Mux_v I__1635 (
            .O(N__8098),
            .I(N__8095));
    Sp12to4 I__1634 (
            .O(N__8095),
            .I(N__8092));
    Span12Mux_h I__1633 (
            .O(N__8092),
            .I(N__8089));
    Odrv12 I__1632 (
            .O(N__8089),
            .I(A_c_14));
    CascadeMux I__1631 (
            .O(N__8086),
            .I(N__8083));
    InMux I__1630 (
            .O(N__8083),
            .I(N__8080));
    LocalMux I__1629 (
            .O(N__8080),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ));
    InMux I__1628 (
            .O(N__8077),
            .I(N__8074));
    LocalMux I__1627 (
            .O(N__8074),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i ));
    InMux I__1626 (
            .O(N__8071),
            .I(N__8068));
    LocalMux I__1625 (
            .O(N__8068),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    InMux I__1624 (
            .O(N__8065),
            .I(N__8062));
    LocalMux I__1623 (
            .O(N__8062),
            .I(N__8059));
    Span12Mux_h I__1622 (
            .O(N__8059),
            .I(N__8056));
    Odrv12 I__1621 (
            .O(N__8056),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ));
    InMux I__1620 (
            .O(N__8053),
            .I(N__8050));
    LocalMux I__1619 (
            .O(N__8050),
            .I(N__8047));
    Odrv4 I__1618 (
            .O(N__8047),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    InMux I__1617 (
            .O(N__8044),
            .I(N__8041));
    LocalMux I__1616 (
            .O(N__8041),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    InMux I__1615 (
            .O(N__8038),
            .I(N__8031));
    InMux I__1614 (
            .O(N__8037),
            .I(N__8025));
    InMux I__1613 (
            .O(N__8036),
            .I(N__8025));
    InMux I__1612 (
            .O(N__8035),
            .I(N__8022));
    InMux I__1611 (
            .O(N__8034),
            .I(N__8019));
    LocalMux I__1610 (
            .O(N__8031),
            .I(N__8016));
    InMux I__1609 (
            .O(N__8030),
            .I(N__8013));
    LocalMux I__1608 (
            .O(N__8025),
            .I(N__8010));
    LocalMux I__1607 (
            .O(N__8022),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1606 (
            .O(N__8019),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv4 I__1605 (
            .O(N__8016),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    LocalMux I__1604 (
            .O(N__8013),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv4 I__1603 (
            .O(N__8010),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    CascadeMux I__1602 (
            .O(N__7999),
            .I(\U712_REG_SM.N_373_cascade_ ));
    InMux I__1601 (
            .O(N__7996),
            .I(N__7993));
    LocalMux I__1600 (
            .O(N__7993),
            .I(\U712_REG_SM.N_130 ));
    InMux I__1599 (
            .O(N__7990),
            .I(N__7986));
    InMux I__1598 (
            .O(N__7989),
            .I(N__7982));
    LocalMux I__1597 (
            .O(N__7986),
            .I(N__7979));
    InMux I__1596 (
            .O(N__7985),
            .I(N__7976));
    LocalMux I__1595 (
            .O(N__7982),
            .I(\U712_REG_SM.un1_REGENn_0_sqmuxa_0 ));
    Odrv4 I__1594 (
            .O(N__7979),
            .I(\U712_REG_SM.un1_REGENn_0_sqmuxa_0 ));
    LocalMux I__1593 (
            .O(N__7976),
            .I(\U712_REG_SM.un1_REGENn_0_sqmuxa_0 ));
    InMux I__1592 (
            .O(N__7969),
            .I(N__7966));
    LocalMux I__1591 (
            .O(N__7966),
            .I(N__7963));
    Odrv4 I__1590 (
            .O(N__7963),
            .I(\U712_CHIP_RAM.N_335 ));
    CascadeMux I__1589 (
            .O(N__7960),
            .I(N__7952));
    InMux I__1588 (
            .O(N__7959),
            .I(N__7948));
    InMux I__1587 (
            .O(N__7958),
            .I(N__7945));
    InMux I__1586 (
            .O(N__7957),
            .I(N__7937));
    CascadeMux I__1585 (
            .O(N__7956),
            .I(N__7932));
    InMux I__1584 (
            .O(N__7955),
            .I(N__7929));
    InMux I__1583 (
            .O(N__7952),
            .I(N__7926));
    InMux I__1582 (
            .O(N__7951),
            .I(N__7923));
    LocalMux I__1581 (
            .O(N__7948),
            .I(N__7918));
    LocalMux I__1580 (
            .O(N__7945),
            .I(N__7918));
    InMux I__1579 (
            .O(N__7944),
            .I(N__7909));
    InMux I__1578 (
            .O(N__7943),
            .I(N__7909));
    InMux I__1577 (
            .O(N__7942),
            .I(N__7909));
    InMux I__1576 (
            .O(N__7941),
            .I(N__7909));
    InMux I__1575 (
            .O(N__7940),
            .I(N__7906));
    LocalMux I__1574 (
            .O(N__7937),
            .I(N__7903));
    InMux I__1573 (
            .O(N__7936),
            .I(N__7896));
    InMux I__1572 (
            .O(N__7935),
            .I(N__7896));
    InMux I__1571 (
            .O(N__7932),
            .I(N__7896));
    LocalMux I__1570 (
            .O(N__7929),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1569 (
            .O(N__7926),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1568 (
            .O(N__7923),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1567 (
            .O(N__7918),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1566 (
            .O(N__7909),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1565 (
            .O(N__7906),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__1564 (
            .O(N__7903),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__1563 (
            .O(N__7896),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    IoInMux I__1562 (
            .O(N__7879),
            .I(N__7876));
    LocalMux I__1561 (
            .O(N__7876),
            .I(N__7873));
    Span12Mux_s11_v I__1560 (
            .O(N__7873),
            .I(N__7870));
    Span12Mux_h I__1559 (
            .O(N__7870),
            .I(N__7867));
    Odrv12 I__1558 (
            .O(N__7867),
            .I(ASn_c));
    CEMux I__1557 (
            .O(N__7864),
            .I(N__7861));
    LocalMux I__1556 (
            .O(N__7861),
            .I(N__7858));
    Span4Mux_h I__1555 (
            .O(N__7858),
            .I(N__7855));
    Odrv4 I__1554 (
            .O(N__7855),
            .I(\U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0 ));
    IoInMux I__1553 (
            .O(N__7852),
            .I(N__7849));
    LocalMux I__1552 (
            .O(N__7849),
            .I(N__7846));
    IoSpan4Mux I__1551 (
            .O(N__7846),
            .I(N__7843));
    Span4Mux_s3_v I__1550 (
            .O(N__7843),
            .I(N__7840));
    Span4Mux_v I__1549 (
            .O(N__7840),
            .I(N__7837));
    Odrv4 I__1548 (
            .O(N__7837),
            .I(N_165_i));
    IoInMux I__1547 (
            .O(N__7834),
            .I(N__7830));
    InMux I__1546 (
            .O(N__7833),
            .I(N__7827));
    LocalMux I__1545 (
            .O(N__7830),
            .I(N__7824));
    LocalMux I__1544 (
            .O(N__7827),
            .I(N__7821));
    Span12Mux_s8_v I__1543 (
            .O(N__7824),
            .I(N__7818));
    Span4Mux_h I__1542 (
            .O(N__7821),
            .I(N__7815));
    Odrv12 I__1541 (
            .O(N__7818),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1540 (
            .O(N__7815),
            .I(CONSTANT_ONE_NET));
    IoInMux I__1539 (
            .O(N__7810),
            .I(N__7807));
    LocalMux I__1538 (
            .O(N__7807),
            .I(N__7804));
    Span4Mux_s2_v I__1537 (
            .O(N__7804),
            .I(N__7801));
    Span4Mux_v I__1536 (
            .O(N__7801),
            .I(N__7798));
    Sp12to4 I__1535 (
            .O(N__7798),
            .I(N__7795));
    Span12Mux_h I__1534 (
            .O(N__7795),
            .I(N__7792));
    Odrv12 I__1533 (
            .O(N__7792),
            .I(RASn_c));
    IoInMux I__1532 (
            .O(N__7789),
            .I(N__7786));
    LocalMux I__1531 (
            .O(N__7786),
            .I(N__7783));
    IoSpan4Mux I__1530 (
            .O(N__7783),
            .I(N__7780));
    IoSpan4Mux I__1529 (
            .O(N__7780),
            .I(N__7777));
    Sp12to4 I__1528 (
            .O(N__7777),
            .I(N__7774));
    Span12Mux_s7_v I__1527 (
            .O(N__7774),
            .I(N__7771));
    Span12Mux_h I__1526 (
            .O(N__7771),
            .I(N__7768));
    Odrv12 I__1525 (
            .O(N__7768),
            .I(WEn_c));
    InMux I__1524 (
            .O(N__7765),
            .I(N__7762));
    LocalMux I__1523 (
            .O(N__7762),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ));
    InMux I__1522 (
            .O(N__7759),
            .I(N__7753));
    InMux I__1521 (
            .O(N__7758),
            .I(N__7753));
    LocalMux I__1520 (
            .O(N__7753),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    IoInMux I__1519 (
            .O(N__7750),
            .I(N__7746));
    IoInMux I__1518 (
            .O(N__7749),
            .I(N__7743));
    LocalMux I__1517 (
            .O(N__7746),
            .I(N__7739));
    LocalMux I__1516 (
            .O(N__7743),
            .I(N__7736));
    IoInMux I__1515 (
            .O(N__7742),
            .I(N__7733));
    Span4Mux_s1_v I__1514 (
            .O(N__7739),
            .I(N__7730));
    IoSpan4Mux I__1513 (
            .O(N__7736),
            .I(N__7727));
    LocalMux I__1512 (
            .O(N__7733),
            .I(N__7724));
    Span4Mux_v I__1511 (
            .O(N__7730),
            .I(N__7721));
    Span4Mux_s2_v I__1510 (
            .O(N__7727),
            .I(N__7718));
    Span4Mux_s2_h I__1509 (
            .O(N__7724),
            .I(N__7715));
    Sp12to4 I__1508 (
            .O(N__7721),
            .I(N__7712));
    Span4Mux_v I__1507 (
            .O(N__7718),
            .I(N__7709));
    Span4Mux_h I__1506 (
            .O(N__7715),
            .I(N__7706));
    Span12Mux_h I__1505 (
            .O(N__7712),
            .I(N__7703));
    Sp12to4 I__1504 (
            .O(N__7709),
            .I(N__7700));
    Sp12to4 I__1503 (
            .O(N__7706),
            .I(N__7697));
    Span12Mux_v I__1502 (
            .O(N__7703),
            .I(N__7689));
    Span12Mux_v I__1501 (
            .O(N__7700),
            .I(N__7689));
    Span12Mux_v I__1500 (
            .O(N__7697),
            .I(N__7689));
    InMux I__1499 (
            .O(N__7696),
            .I(N__7686));
    Odrv12 I__1498 (
            .O(N__7689),
            .I(TACK_EN));
    LocalMux I__1497 (
            .O(N__7686),
            .I(TACK_EN));
    CascadeMux I__1496 (
            .O(N__7681),
            .I(N__7677));
    CascadeMux I__1495 (
            .O(N__7680),
            .I(N__7674));
    InMux I__1494 (
            .O(N__7677),
            .I(N__7670));
    InMux I__1493 (
            .O(N__7674),
            .I(N__7667));
    InMux I__1492 (
            .O(N__7673),
            .I(N__7664));
    LocalMux I__1491 (
            .O(N__7670),
            .I(N__7661));
    LocalMux I__1490 (
            .O(N__7667),
            .I(\U712_REG_SM.N_328 ));
    LocalMux I__1489 (
            .O(N__7664),
            .I(\U712_REG_SM.N_328 ));
    Odrv4 I__1488 (
            .O(N__7661),
            .I(\U712_REG_SM.N_328 ));
    CascadeMux I__1487 (
            .O(N__7654),
            .I(N__7651));
    InMux I__1486 (
            .O(N__7651),
            .I(N__7648));
    LocalMux I__1485 (
            .O(N__7648),
            .I(\U712_REG_SM.N_406 ));
    InMux I__1484 (
            .O(N__7645),
            .I(N__7642));
    LocalMux I__1483 (
            .O(N__7642),
            .I(N__7637));
    InMux I__1482 (
            .O(N__7641),
            .I(N__7633));
    InMux I__1481 (
            .O(N__7640),
            .I(N__7629));
    Span4Mux_h I__1480 (
            .O(N__7637),
            .I(N__7626));
    InMux I__1479 (
            .O(N__7636),
            .I(N__7623));
    LocalMux I__1478 (
            .O(N__7633),
            .I(N__7620));
    InMux I__1477 (
            .O(N__7632),
            .I(N__7617));
    LocalMux I__1476 (
            .O(N__7629),
            .I(N__7614));
    Odrv4 I__1475 (
            .O(N__7626),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1474 (
            .O(N__7623),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1473 (
            .O(N__7620),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__1472 (
            .O(N__7617),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__1471 (
            .O(N__7614),
            .I(DBR_SYNCZ0Z_1));
    CascadeMux I__1470 (
            .O(N__7603),
            .I(\U712_REG_SM.N_330_cascade_ ));
    InMux I__1469 (
            .O(N__7600),
            .I(N__7597));
    LocalMux I__1468 (
            .O(N__7597),
            .I(N__7591));
    InMux I__1467 (
            .O(N__7596),
            .I(N__7588));
    InMux I__1466 (
            .O(N__7595),
            .I(N__7583));
    InMux I__1465 (
            .O(N__7594),
            .I(N__7583));
    Odrv4 I__1464 (
            .O(N__7591),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    LocalMux I__1463 (
            .O(N__7588),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    LocalMux I__1462 (
            .O(N__7583),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    InMux I__1461 (
            .O(N__7576),
            .I(N__7573));
    LocalMux I__1460 (
            .O(N__7573),
            .I(\U712_REG_SM.STATE_COUNTc_0_0 ));
    InMux I__1459 (
            .O(N__7570),
            .I(N__7563));
    InMux I__1458 (
            .O(N__7569),
            .I(N__7558));
    InMux I__1457 (
            .O(N__7568),
            .I(N__7558));
    InMux I__1456 (
            .O(N__7567),
            .I(N__7555));
    InMux I__1455 (
            .O(N__7566),
            .I(N__7552));
    LocalMux I__1454 (
            .O(N__7563),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1453 (
            .O(N__7558),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1452 (
            .O(N__7555),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__1451 (
            .O(N__7552),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    CascadeMux I__1450 (
            .O(N__7543),
            .I(N__7539));
    InMux I__1449 (
            .O(N__7542),
            .I(N__7528));
    InMux I__1448 (
            .O(N__7539),
            .I(N__7528));
    CascadeMux I__1447 (
            .O(N__7538),
            .I(N__7523));
    CascadeMux I__1446 (
            .O(N__7537),
            .I(N__7519));
    InMux I__1445 (
            .O(N__7536),
            .I(N__7516));
    CascadeMux I__1444 (
            .O(N__7535),
            .I(N__7513));
    CascadeMux I__1443 (
            .O(N__7534),
            .I(N__7510));
    CascadeMux I__1442 (
            .O(N__7533),
            .I(N__7507));
    LocalMux I__1441 (
            .O(N__7528),
            .I(N__7503));
    InMux I__1440 (
            .O(N__7527),
            .I(N__7498));
    InMux I__1439 (
            .O(N__7526),
            .I(N__7498));
    InMux I__1438 (
            .O(N__7523),
            .I(N__7493));
    InMux I__1437 (
            .O(N__7522),
            .I(N__7493));
    InMux I__1436 (
            .O(N__7519),
            .I(N__7490));
    LocalMux I__1435 (
            .O(N__7516),
            .I(N__7487));
    InMux I__1434 (
            .O(N__7513),
            .I(N__7484));
    InMux I__1433 (
            .O(N__7510),
            .I(N__7477));
    InMux I__1432 (
            .O(N__7507),
            .I(N__7477));
    InMux I__1431 (
            .O(N__7506),
            .I(N__7477));
    Odrv12 I__1430 (
            .O(N__7503),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1429 (
            .O(N__7498),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1428 (
            .O(N__7493),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1427 (
            .O(N__7490),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1426 (
            .O(N__7487),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1425 (
            .O(N__7484),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1424 (
            .O(N__7477),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__1423 (
            .O(N__7462),
            .I(N__7459));
    LocalMux I__1422 (
            .O(N__7459),
            .I(\U712_REG_SM.N_373 ));
    InMux I__1421 (
            .O(N__7456),
            .I(N__7452));
    InMux I__1420 (
            .O(N__7455),
            .I(N__7449));
    LocalMux I__1419 (
            .O(N__7452),
            .I(N__7446));
    LocalMux I__1418 (
            .O(N__7449),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    Odrv4 I__1417 (
            .O(N__7446),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    InMux I__1416 (
            .O(N__7441),
            .I(N__7438));
    LocalMux I__1415 (
            .O(N__7438),
            .I(N__7435));
    Span4Mux_h I__1414 (
            .O(N__7435),
            .I(N__7431));
    InMux I__1413 (
            .O(N__7434),
            .I(N__7428));
    Span4Mux_v I__1412 (
            .O(N__7431),
            .I(N__7423));
    LocalMux I__1411 (
            .O(N__7428),
            .I(N__7423));
    Span4Mux_v I__1410 (
            .O(N__7423),
            .I(N__7419));
    InMux I__1409 (
            .O(N__7422),
            .I(N__7416));
    Odrv4 I__1408 (
            .O(N__7419),
            .I(REG_CYCLEm));
    LocalMux I__1407 (
            .O(N__7416),
            .I(REG_CYCLEm));
    IoInMux I__1406 (
            .O(N__7411),
            .I(N__7408));
    LocalMux I__1405 (
            .O(N__7408),
            .I(N__7405));
    Span4Mux_s1_v I__1404 (
            .O(N__7405),
            .I(N__7402));
    Span4Mux_v I__1403 (
            .O(N__7402),
            .I(N__7399));
    Sp12to4 I__1402 (
            .O(N__7399),
            .I(N__7396));
    Span12Mux_s10_h I__1401 (
            .O(N__7396),
            .I(N__7393));
    Span12Mux_v I__1400 (
            .O(N__7393),
            .I(N__7390));
    Odrv12 I__1399 (
            .O(N__7390),
            .I(N_167_i));
    InMux I__1398 (
            .O(N__7387),
            .I(N__7381));
    InMux I__1397 (
            .O(N__7386),
            .I(N__7376));
    InMux I__1396 (
            .O(N__7385),
            .I(N__7376));
    InMux I__1395 (
            .O(N__7384),
            .I(N__7373));
    LocalMux I__1394 (
            .O(N__7381),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__1393 (
            .O(N__7376),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__1392 (
            .O(N__7373),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    InMux I__1391 (
            .O(N__7366),
            .I(N__7363));
    LocalMux I__1390 (
            .O(N__7363),
            .I(\U712_CHIP_RAM.N_321 ));
    CascadeMux I__1389 (
            .O(N__7360),
            .I(\U712_CHIP_RAM.N_321_cascade_ ));
    InMux I__1388 (
            .O(N__7357),
            .I(N__7353));
    InMux I__1387 (
            .O(N__7356),
            .I(N__7350));
    LocalMux I__1386 (
            .O(N__7353),
            .I(\U712_CHIP_RAM.N_20_0 ));
    LocalMux I__1385 (
            .O(N__7350),
            .I(\U712_CHIP_RAM.N_20_0 ));
    CascadeMux I__1384 (
            .O(N__7345),
            .I(N__7341));
    CascadeMux I__1383 (
            .O(N__7344),
            .I(N__7337));
    InMux I__1382 (
            .O(N__7341),
            .I(N__7332));
    InMux I__1381 (
            .O(N__7340),
            .I(N__7329));
    InMux I__1380 (
            .O(N__7337),
            .I(N__7326));
    InMux I__1379 (
            .O(N__7336),
            .I(N__7322));
    InMux I__1378 (
            .O(N__7335),
            .I(N__7319));
    LocalMux I__1377 (
            .O(N__7332),
            .I(N__7316));
    LocalMux I__1376 (
            .O(N__7329),
            .I(N__7313));
    LocalMux I__1375 (
            .O(N__7326),
            .I(N__7310));
    InMux I__1374 (
            .O(N__7325),
            .I(N__7299));
    LocalMux I__1373 (
            .O(N__7322),
            .I(N__7294));
    LocalMux I__1372 (
            .O(N__7319),
            .I(N__7294));
    Span4Mux_h I__1371 (
            .O(N__7316),
            .I(N__7291));
    Span4Mux_h I__1370 (
            .O(N__7313),
            .I(N__7286));
    Span4Mux_h I__1369 (
            .O(N__7310),
            .I(N__7286));
    InMux I__1368 (
            .O(N__7309),
            .I(N__7281));
    InMux I__1367 (
            .O(N__7308),
            .I(N__7281));
    InMux I__1366 (
            .O(N__7307),
            .I(N__7278));
    InMux I__1365 (
            .O(N__7306),
            .I(N__7273));
    InMux I__1364 (
            .O(N__7305),
            .I(N__7273));
    InMux I__1363 (
            .O(N__7304),
            .I(N__7266));
    InMux I__1362 (
            .O(N__7303),
            .I(N__7266));
    InMux I__1361 (
            .O(N__7302),
            .I(N__7266));
    LocalMux I__1360 (
            .O(N__7299),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1359 (
            .O(N__7294),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1358 (
            .O(N__7291),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1357 (
            .O(N__7286),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1356 (
            .O(N__7281),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1355 (
            .O(N__7278),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1354 (
            .O(N__7273),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1353 (
            .O(N__7266),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__1352 (
            .O(N__7249),
            .I(\U712_CHIP_RAM.m77_0_a2_0_2_cascade_ ));
    CascadeMux I__1351 (
            .O(N__7246),
            .I(N__7240));
    InMux I__1350 (
            .O(N__7245),
            .I(N__7237));
    InMux I__1349 (
            .O(N__7244),
            .I(N__7232));
    InMux I__1348 (
            .O(N__7243),
            .I(N__7232));
    InMux I__1347 (
            .O(N__7240),
            .I(N__7229));
    LocalMux I__1346 (
            .O(N__7237),
            .I(N__7226));
    LocalMux I__1345 (
            .O(N__7232),
            .I(N__7223));
    LocalMux I__1344 (
            .O(N__7229),
            .I(N__7218));
    Span4Mux_h I__1343 (
            .O(N__7226),
            .I(N__7215));
    Span4Mux_v I__1342 (
            .O(N__7223),
            .I(N__7212));
    InMux I__1341 (
            .O(N__7222),
            .I(N__7209));
    InMux I__1340 (
            .O(N__7221),
            .I(N__7206));
    Odrv4 I__1339 (
            .O(N__7218),
            .I(\U712_CHIP_RAM.N_307 ));
    Odrv4 I__1338 (
            .O(N__7215),
            .I(\U712_CHIP_RAM.N_307 ));
    Odrv4 I__1337 (
            .O(N__7212),
            .I(\U712_CHIP_RAM.N_307 ));
    LocalMux I__1336 (
            .O(N__7209),
            .I(\U712_CHIP_RAM.N_307 ));
    LocalMux I__1335 (
            .O(N__7206),
            .I(\U712_CHIP_RAM.N_307 ));
    CascadeMux I__1334 (
            .O(N__7195),
            .I(N__7191));
    InMux I__1333 (
            .O(N__7194),
            .I(N__7182));
    InMux I__1332 (
            .O(N__7191),
            .I(N__7179));
    CascadeMux I__1331 (
            .O(N__7190),
            .I(N__7176));
    InMux I__1330 (
            .O(N__7189),
            .I(N__7173));
    CascadeMux I__1329 (
            .O(N__7188),
            .I(N__7163));
    InMux I__1328 (
            .O(N__7187),
            .I(N__7156));
    InMux I__1327 (
            .O(N__7186),
            .I(N__7151));
    InMux I__1326 (
            .O(N__7185),
            .I(N__7151));
    LocalMux I__1325 (
            .O(N__7182),
            .I(N__7148));
    LocalMux I__1324 (
            .O(N__7179),
            .I(N__7145));
    InMux I__1323 (
            .O(N__7176),
            .I(N__7142));
    LocalMux I__1322 (
            .O(N__7173),
            .I(N__7139));
    InMux I__1321 (
            .O(N__7172),
            .I(N__7136));
    CascadeMux I__1320 (
            .O(N__7171),
            .I(N__7133));
    CascadeMux I__1319 (
            .O(N__7170),
            .I(N__7130));
    InMux I__1318 (
            .O(N__7169),
            .I(N__7120));
    InMux I__1317 (
            .O(N__7168),
            .I(N__7117));
    InMux I__1316 (
            .O(N__7167),
            .I(N__7110));
    InMux I__1315 (
            .O(N__7166),
            .I(N__7110));
    InMux I__1314 (
            .O(N__7163),
            .I(N__7110));
    InMux I__1313 (
            .O(N__7162),
            .I(N__7107));
    InMux I__1312 (
            .O(N__7161),
            .I(N__7102));
    InMux I__1311 (
            .O(N__7160),
            .I(N__7102));
    InMux I__1310 (
            .O(N__7159),
            .I(N__7099));
    LocalMux I__1309 (
            .O(N__7156),
            .I(N__7096));
    LocalMux I__1308 (
            .O(N__7151),
            .I(N__7091));
    Span4Mux_h I__1307 (
            .O(N__7148),
            .I(N__7091));
    Span4Mux_v I__1306 (
            .O(N__7145),
            .I(N__7082));
    LocalMux I__1305 (
            .O(N__7142),
            .I(N__7082));
    Span4Mux_v I__1304 (
            .O(N__7139),
            .I(N__7082));
    LocalMux I__1303 (
            .O(N__7136),
            .I(N__7082));
    InMux I__1302 (
            .O(N__7133),
            .I(N__7075));
    InMux I__1301 (
            .O(N__7130),
            .I(N__7075));
    InMux I__1300 (
            .O(N__7129),
            .I(N__7075));
    InMux I__1299 (
            .O(N__7128),
            .I(N__7062));
    InMux I__1298 (
            .O(N__7127),
            .I(N__7062));
    InMux I__1297 (
            .O(N__7126),
            .I(N__7062));
    InMux I__1296 (
            .O(N__7125),
            .I(N__7062));
    InMux I__1295 (
            .O(N__7124),
            .I(N__7062));
    InMux I__1294 (
            .O(N__7123),
            .I(N__7062));
    LocalMux I__1293 (
            .O(N__7120),
            .I(N__7051));
    LocalMux I__1292 (
            .O(N__7117),
            .I(N__7051));
    LocalMux I__1291 (
            .O(N__7110),
            .I(N__7051));
    LocalMux I__1290 (
            .O(N__7107),
            .I(N__7051));
    LocalMux I__1289 (
            .O(N__7102),
            .I(N__7051));
    LocalMux I__1288 (
            .O(N__7099),
            .I(N__7048));
    Odrv12 I__1287 (
            .O(N__7096),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1286 (
            .O(N__7091),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1285 (
            .O(N__7082),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1284 (
            .O(N__7075),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1283 (
            .O(N__7062),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1282 (
            .O(N__7051),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1281 (
            .O(N__7048),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1280 (
            .O(N__7033),
            .I(N__7027));
    InMux I__1279 (
            .O(N__7032),
            .I(N__7013));
    InMux I__1278 (
            .O(N__7031),
            .I(N__7008));
    InMux I__1277 (
            .O(N__7030),
            .I(N__7008));
    LocalMux I__1276 (
            .O(N__7027),
            .I(N__7005));
    InMux I__1275 (
            .O(N__7026),
            .I(N__6990));
    InMux I__1274 (
            .O(N__7025),
            .I(N__6990));
    InMux I__1273 (
            .O(N__7024),
            .I(N__6990));
    InMux I__1272 (
            .O(N__7023),
            .I(N__6990));
    CascadeMux I__1271 (
            .O(N__7022),
            .I(N__6987));
    CascadeMux I__1270 (
            .O(N__7021),
            .I(N__6979));
    InMux I__1269 (
            .O(N__7020),
            .I(N__6972));
    InMux I__1268 (
            .O(N__7019),
            .I(N__6972));
    InMux I__1267 (
            .O(N__7018),
            .I(N__6969));
    InMux I__1266 (
            .O(N__7017),
            .I(N__6966));
    InMux I__1265 (
            .O(N__7016),
            .I(N__6963));
    LocalMux I__1264 (
            .O(N__7013),
            .I(N__6960));
    LocalMux I__1263 (
            .O(N__7008),
            .I(N__6955));
    Span4Mux_h I__1262 (
            .O(N__7005),
            .I(N__6955));
    InMux I__1261 (
            .O(N__7004),
            .I(N__6948));
    InMux I__1260 (
            .O(N__7003),
            .I(N__6948));
    InMux I__1259 (
            .O(N__7002),
            .I(N__6948));
    InMux I__1258 (
            .O(N__7001),
            .I(N__6945));
    InMux I__1257 (
            .O(N__7000),
            .I(N__6940));
    InMux I__1256 (
            .O(N__6999),
            .I(N__6940));
    LocalMux I__1255 (
            .O(N__6990),
            .I(N__6937));
    InMux I__1254 (
            .O(N__6987),
            .I(N__6926));
    InMux I__1253 (
            .O(N__6986),
            .I(N__6926));
    InMux I__1252 (
            .O(N__6985),
            .I(N__6926));
    InMux I__1251 (
            .O(N__6984),
            .I(N__6926));
    InMux I__1250 (
            .O(N__6983),
            .I(N__6926));
    InMux I__1249 (
            .O(N__6982),
            .I(N__6917));
    InMux I__1248 (
            .O(N__6979),
            .I(N__6917));
    InMux I__1247 (
            .O(N__6978),
            .I(N__6917));
    InMux I__1246 (
            .O(N__6977),
            .I(N__6917));
    LocalMux I__1245 (
            .O(N__6972),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1244 (
            .O(N__6969),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1243 (
            .O(N__6966),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1242 (
            .O(N__6963),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1241 (
            .O(N__6960),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1240 (
            .O(N__6955),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1239 (
            .O(N__6948),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1238 (
            .O(N__6945),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1237 (
            .O(N__6940),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1236 (
            .O(N__6937),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1235 (
            .O(N__6926),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1234 (
            .O(N__6917),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    CascadeMux I__1233 (
            .O(N__6892),
            .I(N__6887));
    InMux I__1232 (
            .O(N__6891),
            .I(N__6882));
    InMux I__1231 (
            .O(N__6890),
            .I(N__6877));
    InMux I__1230 (
            .O(N__6887),
            .I(N__6877));
    InMux I__1229 (
            .O(N__6886),
            .I(N__6874));
    InMux I__1228 (
            .O(N__6885),
            .I(N__6870));
    LocalMux I__1227 (
            .O(N__6882),
            .I(N__6867));
    LocalMux I__1226 (
            .O(N__6877),
            .I(N__6860));
    LocalMux I__1225 (
            .O(N__6874),
            .I(N__6852));
    InMux I__1224 (
            .O(N__6873),
            .I(N__6849));
    LocalMux I__1223 (
            .O(N__6870),
            .I(N__6846));
    Span4Mux_v I__1222 (
            .O(N__6867),
            .I(N__6843));
    InMux I__1221 (
            .O(N__6866),
            .I(N__6840));
    InMux I__1220 (
            .O(N__6865),
            .I(N__6833));
    InMux I__1219 (
            .O(N__6864),
            .I(N__6833));
    InMux I__1218 (
            .O(N__6863),
            .I(N__6833));
    Span4Mux_h I__1217 (
            .O(N__6860),
            .I(N__6830));
    InMux I__1216 (
            .O(N__6859),
            .I(N__6827));
    InMux I__1215 (
            .O(N__6858),
            .I(N__6822));
    InMux I__1214 (
            .O(N__6857),
            .I(N__6822));
    InMux I__1213 (
            .O(N__6856),
            .I(N__6819));
    InMux I__1212 (
            .O(N__6855),
            .I(N__6816));
    Odrv4 I__1211 (
            .O(N__6852),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1210 (
            .O(N__6849),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1209 (
            .O(N__6846),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1208 (
            .O(N__6843),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1207 (
            .O(N__6840),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1206 (
            .O(N__6833),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1205 (
            .O(N__6830),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1204 (
            .O(N__6827),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1203 (
            .O(N__6822),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1202 (
            .O(N__6819),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1201 (
            .O(N__6816),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    CascadeMux I__1200 (
            .O(N__6793),
            .I(N__6788));
    CascadeMux I__1199 (
            .O(N__6792),
            .I(N__6785));
    InMux I__1198 (
            .O(N__6791),
            .I(N__6779));
    InMux I__1197 (
            .O(N__6788),
            .I(N__6779));
    InMux I__1196 (
            .O(N__6785),
            .I(N__6774));
    InMux I__1195 (
            .O(N__6784),
            .I(N__6768));
    LocalMux I__1194 (
            .O(N__6779),
            .I(N__6765));
    CascadeMux I__1193 (
            .O(N__6778),
            .I(N__6761));
    InMux I__1192 (
            .O(N__6777),
            .I(N__6755));
    LocalMux I__1191 (
            .O(N__6774),
            .I(N__6749));
    InMux I__1190 (
            .O(N__6773),
            .I(N__6746));
    InMux I__1189 (
            .O(N__6772),
            .I(N__6741));
    InMux I__1188 (
            .O(N__6771),
            .I(N__6741));
    LocalMux I__1187 (
            .O(N__6768),
            .I(N__6736));
    Span4Mux_h I__1186 (
            .O(N__6765),
            .I(N__6736));
    InMux I__1185 (
            .O(N__6764),
            .I(N__6731));
    InMux I__1184 (
            .O(N__6761),
            .I(N__6731));
    InMux I__1183 (
            .O(N__6760),
            .I(N__6726));
    InMux I__1182 (
            .O(N__6759),
            .I(N__6726));
    InMux I__1181 (
            .O(N__6758),
            .I(N__6723));
    LocalMux I__1180 (
            .O(N__6755),
            .I(N__6720));
    InMux I__1179 (
            .O(N__6754),
            .I(N__6715));
    InMux I__1178 (
            .O(N__6753),
            .I(N__6715));
    InMux I__1177 (
            .O(N__6752),
            .I(N__6712));
    Odrv4 I__1176 (
            .O(N__6749),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1175 (
            .O(N__6746),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1174 (
            .O(N__6741),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1173 (
            .O(N__6736),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1172 (
            .O(N__6731),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1171 (
            .O(N__6726),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1170 (
            .O(N__6723),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1169 (
            .O(N__6720),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1168 (
            .O(N__6715),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1167 (
            .O(N__6712),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1166 (
            .O(N__6691),
            .I(N__6688));
    LocalMux I__1165 (
            .O(N__6688),
            .I(N__6685));
    Span4Mux_h I__1164 (
            .O(N__6685),
            .I(N__6682));
    Span4Mux_v I__1163 (
            .O(N__6682),
            .I(N__6679));
    Odrv4 I__1162 (
            .O(N__6679),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_6 ));
    SRMux I__1161 (
            .O(N__6676),
            .I(N__6672));
    SRMux I__1160 (
            .O(N__6675),
            .I(N__6669));
    LocalMux I__1159 (
            .O(N__6672),
            .I(N__6664));
    LocalMux I__1158 (
            .O(N__6669),
            .I(N__6664));
    Span4Mux_v I__1157 (
            .O(N__6664),
            .I(N__6661));
    Odrv4 I__1156 (
            .O(N__6661),
            .I(\U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ));
    InMux I__1155 (
            .O(N__6658),
            .I(N__6654));
    InMux I__1154 (
            .O(N__6657),
            .I(N__6651));
    LocalMux I__1153 (
            .O(N__6654),
            .I(N__6646));
    LocalMux I__1152 (
            .O(N__6651),
            .I(N__6646));
    Span4Mux_h I__1151 (
            .O(N__6646),
            .I(N__6642));
    InMux I__1150 (
            .O(N__6645),
            .I(N__6639));
    Odrv4 I__1149 (
            .O(N__6642),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__1148 (
            .O(N__6639),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    IoInMux I__1147 (
            .O(N__6634),
            .I(N__6631));
    LocalMux I__1146 (
            .O(N__6631),
            .I(N__6628));
    IoSpan4Mux I__1145 (
            .O(N__6628),
            .I(N__6625));
    Span4Mux_s2_v I__1144 (
            .O(N__6625),
            .I(N__6622));
    Sp12to4 I__1143 (
            .O(N__6622),
            .I(N__6619));
    Span12Mux_s9_v I__1142 (
            .O(N__6619),
            .I(N__6616));
    Odrv12 I__1141 (
            .O(N__6616),
            .I(N_202_i));
    InMux I__1140 (
            .O(N__6613),
            .I(N__6610));
    LocalMux I__1139 (
            .O(N__6610),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__1138 (
            .O(N__6607),
            .I(N__6604));
    LocalMux I__1137 (
            .O(N__6604),
            .I(N__6599));
    InMux I__1136 (
            .O(N__6603),
            .I(N__6596));
    InMux I__1135 (
            .O(N__6602),
            .I(N__6593));
    Odrv12 I__1134 (
            .O(N__6599),
            .I(\U712_CHIP_RAM.N_305 ));
    LocalMux I__1133 (
            .O(N__6596),
            .I(\U712_CHIP_RAM.N_305 ));
    LocalMux I__1132 (
            .O(N__6593),
            .I(\U712_CHIP_RAM.N_305 ));
    CascadeMux I__1131 (
            .O(N__6586),
            .I(\U712_CHIP_RAM.m123_i_2_cascade_ ));
    InMux I__1130 (
            .O(N__6583),
            .I(N__6580));
    LocalMux I__1129 (
            .O(N__6580),
            .I(N__6577));
    Span4Mux_v I__1128 (
            .O(N__6577),
            .I(N__6574));
    Span4Mux_v I__1127 (
            .O(N__6574),
            .I(N__6571));
    Sp12to4 I__1126 (
            .O(N__6571),
            .I(N__6568));
    Span12Mux_h I__1125 (
            .O(N__6568),
            .I(N__6565));
    Odrv12 I__1124 (
            .O(N__6565),
            .I(A_c_15));
    InMux I__1123 (
            .O(N__6562),
            .I(N__6559));
    LocalMux I__1122 (
            .O(N__6559),
            .I(N__6556));
    Odrv12 I__1121 (
            .O(N__6556),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ));
    CascadeMux I__1120 (
            .O(N__6553),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ));
    InMux I__1119 (
            .O(N__6550),
            .I(N__6547));
    LocalMux I__1118 (
            .O(N__6547),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_2_0 ));
    InMux I__1117 (
            .O(N__6544),
            .I(N__6541));
    LocalMux I__1116 (
            .O(N__6541),
            .I(\U712_CHIP_RAM.N_390 ));
    InMux I__1115 (
            .O(N__6538),
            .I(N__6535));
    LocalMux I__1114 (
            .O(N__6535),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_2_3 ));
    IoInMux I__1113 (
            .O(N__6532),
            .I(N__6529));
    LocalMux I__1112 (
            .O(N__6529),
            .I(N__6526));
    IoSpan4Mux I__1111 (
            .O(N__6526),
            .I(N__6523));
    Span4Mux_s2_v I__1110 (
            .O(N__6523),
            .I(N__6519));
    InMux I__1109 (
            .O(N__6522),
            .I(N__6516));
    Sp12to4 I__1108 (
            .O(N__6519),
            .I(N__6513));
    LocalMux I__1107 (
            .O(N__6516),
            .I(N__6510));
    Span12Mux_s8_v I__1106 (
            .O(N__6513),
            .I(N__6507));
    Span4Mux_v I__1105 (
            .O(N__6510),
            .I(N__6504));
    Span12Mux_h I__1104 (
            .O(N__6507),
            .I(N__6501));
    Sp12to4 I__1103 (
            .O(N__6504),
            .I(N__6498));
    Span12Mux_v I__1102 (
            .O(N__6501),
            .I(N__6495));
    Span12Mux_h I__1101 (
            .O(N__6498),
            .I(N__6492));
    Odrv12 I__1100 (
            .O(N__6495),
            .I(A_c_11));
    Odrv12 I__1099 (
            .O(N__6492),
            .I(A_c_11));
    InMux I__1098 (
            .O(N__6487),
            .I(N__6484));
    LocalMux I__1097 (
            .O(N__6484),
            .I(N__6481));
    Odrv12 I__1096 (
            .O(N__6481),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ));
    InMux I__1095 (
            .O(N__6478),
            .I(N__6475));
    LocalMux I__1094 (
            .O(N__6475),
            .I(N__6472));
    Span12Mux_v I__1093 (
            .O(N__6472),
            .I(N__6469));
    Span12Mux_h I__1092 (
            .O(N__6469),
            .I(N__6466));
    Odrv12 I__1091 (
            .O(N__6466),
            .I(A_c_3));
    InMux I__1090 (
            .O(N__6463),
            .I(N__6460));
    LocalMux I__1089 (
            .O(N__6460),
            .I(N__6457));
    Odrv4 I__1088 (
            .O(N__6457),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ));
    InMux I__1087 (
            .O(N__6454),
            .I(N__6451));
    LocalMux I__1086 (
            .O(N__6451),
            .I(N__6448));
    Span4Mux_v I__1085 (
            .O(N__6448),
            .I(N__6445));
    Span4Mux_v I__1084 (
            .O(N__6445),
            .I(N__6442));
    Sp12to4 I__1083 (
            .O(N__6442),
            .I(N__6439));
    Span12Mux_h I__1082 (
            .O(N__6439),
            .I(N__6436));
    Odrv12 I__1081 (
            .O(N__6436),
            .I(A_c_5));
    InMux I__1080 (
            .O(N__6433),
            .I(N__6430));
    LocalMux I__1079 (
            .O(N__6430),
            .I(N__6427));
    Odrv4 I__1078 (
            .O(N__6427),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ));
    InMux I__1077 (
            .O(N__6424),
            .I(N__6421));
    LocalMux I__1076 (
            .O(N__6421),
            .I(N__6418));
    Span12Mux_v I__1075 (
            .O(N__6418),
            .I(N__6415));
    Span12Mux_h I__1074 (
            .O(N__6415),
            .I(N__6412));
    Odrv12 I__1073 (
            .O(N__6412),
            .I(A_c_6));
    CEMux I__1072 (
            .O(N__6409),
            .I(N__6404));
    CEMux I__1071 (
            .O(N__6408),
            .I(N__6401));
    CEMux I__1070 (
            .O(N__6407),
            .I(N__6398));
    LocalMux I__1069 (
            .O(N__6404),
            .I(N__6395));
    LocalMux I__1068 (
            .O(N__6401),
            .I(N__6392));
    LocalMux I__1067 (
            .O(N__6398),
            .I(N__6389));
    Span4Mux_h I__1066 (
            .O(N__6395),
            .I(N__6386));
    Span4Mux_h I__1065 (
            .O(N__6392),
            .I(N__6383));
    Span4Mux_h I__1064 (
            .O(N__6389),
            .I(N__6380));
    Odrv4 I__1063 (
            .O(N__6386),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    Odrv4 I__1062 (
            .O(N__6383),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    Odrv4 I__1061 (
            .O(N__6380),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ));
    InMux I__1060 (
            .O(N__6373),
            .I(N__6370));
    LocalMux I__1059 (
            .O(N__6370),
            .I(N__6366));
    InMux I__1058 (
            .O(N__6369),
            .I(N__6363));
    Span4Mux_h I__1057 (
            .O(N__6366),
            .I(N__6360));
    LocalMux I__1056 (
            .O(N__6363),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_4 ));
    Odrv4 I__1055 (
            .O(N__6360),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_4 ));
    InMux I__1054 (
            .O(N__6355),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_3 ));
    InMux I__1053 (
            .O(N__6352),
            .I(N__6349));
    LocalMux I__1052 (
            .O(N__6349),
            .I(N__6345));
    InMux I__1051 (
            .O(N__6348),
            .I(N__6342));
    Span4Mux_v I__1050 (
            .O(N__6345),
            .I(N__6339));
    LocalMux I__1049 (
            .O(N__6342),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_5 ));
    Odrv4 I__1048 (
            .O(N__6339),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_5 ));
    InMux I__1047 (
            .O(N__6334),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_4 ));
    InMux I__1046 (
            .O(N__6331),
            .I(N__6328));
    LocalMux I__1045 (
            .O(N__6328),
            .I(N__6324));
    InMux I__1044 (
            .O(N__6327),
            .I(N__6321));
    Span4Mux_v I__1043 (
            .O(N__6324),
            .I(N__6318));
    LocalMux I__1042 (
            .O(N__6321),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_6 ));
    Odrv4 I__1041 (
            .O(N__6318),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_6 ));
    InMux I__1040 (
            .O(N__6313),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_5 ));
    InMux I__1039 (
            .O(N__6310),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_6 ));
    InMux I__1038 (
            .O(N__6307),
            .I(N__6304));
    LocalMux I__1037 (
            .O(N__6304),
            .I(N__6301));
    Span12Mux_v I__1036 (
            .O(N__6301),
            .I(N__6298));
    Span12Mux_h I__1035 (
            .O(N__6298),
            .I(N__6295));
    Odrv12 I__1034 (
            .O(N__6295),
            .I(A_c_12));
    IoInMux I__1033 (
            .O(N__6292),
            .I(N__6289));
    LocalMux I__1032 (
            .O(N__6289),
            .I(N__6286));
    Span4Mux_s0_v I__1031 (
            .O(N__6286),
            .I(N__6283));
    Span4Mux_v I__1030 (
            .O(N__6283),
            .I(N__6280));
    Span4Mux_v I__1029 (
            .O(N__6280),
            .I(N__6277));
    Sp12to4 I__1028 (
            .O(N__6277),
            .I(N__6273));
    InMux I__1027 (
            .O(N__6276),
            .I(N__6270));
    Span12Mux_h I__1026 (
            .O(N__6273),
            .I(N__6267));
    LocalMux I__1025 (
            .O(N__6270),
            .I(N__6264));
    Span12Mux_v I__1024 (
            .O(N__6267),
            .I(N__6259));
    Span12Mux_h I__1023 (
            .O(N__6264),
            .I(N__6259));
    Odrv12 I__1022 (
            .O(N__6259),
            .I(A_c_10));
    InMux I__1021 (
            .O(N__6256),
            .I(N__6252));
    InMux I__1020 (
            .O(N__6255),
            .I(N__6249));
    LocalMux I__1019 (
            .O(N__6252),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_3 ));
    LocalMux I__1018 (
            .O(N__6249),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_3 ));
    InMux I__1017 (
            .O(N__6244),
            .I(N__6240));
    InMux I__1016 (
            .O(N__6243),
            .I(N__6237));
    LocalMux I__1015 (
            .O(N__6240),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_2 ));
    LocalMux I__1014 (
            .O(N__6237),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_2 ));
    CascadeMux I__1013 (
            .O(N__6232),
            .I(N__6227));
    InMux I__1012 (
            .O(N__6231),
            .I(N__6224));
    InMux I__1011 (
            .O(N__6230),
            .I(N__6221));
    InMux I__1010 (
            .O(N__6227),
            .I(N__6218));
    LocalMux I__1009 (
            .O(N__6224),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ));
    LocalMux I__1008 (
            .O(N__6221),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ));
    LocalMux I__1007 (
            .O(N__6218),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ));
    InMux I__1006 (
            .O(N__6211),
            .I(N__6207));
    InMux I__1005 (
            .O(N__6210),
            .I(N__6204));
    LocalMux I__1004 (
            .O(N__6207),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_7 ));
    LocalMux I__1003 (
            .O(N__6204),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_7 ));
    InMux I__1002 (
            .O(N__6199),
            .I(N__6196));
    LocalMux I__1001 (
            .O(N__6196),
            .I(N__6193));
    Odrv4 I__1000 (
            .O(N__6193),
            .I(\U712_CHIP_RAM.m93_i_a2_5 ));
    SRMux I__999 (
            .O(N__6190),
            .I(N__6187));
    LocalMux I__998 (
            .O(N__6187),
            .I(N__6183));
    InMux I__997 (
            .O(N__6186),
            .I(N__6180));
    Span4Mux_v I__996 (
            .O(N__6183),
            .I(N__6177));
    LocalMux I__995 (
            .O(N__6180),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    Odrv4 I__994 (
            .O(N__6177),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__993 (
            .O(N__6172),
            .I(N__6169));
    LocalMux I__992 (
            .O(N__6169),
            .I(N__6164));
    InMux I__991 (
            .O(N__6168),
            .I(N__6161));
    InMux I__990 (
            .O(N__6167),
            .I(N__6158));
    Odrv4 I__989 (
            .O(N__6164),
            .I(\U712_CHIP_RAM.N_304 ));
    LocalMux I__988 (
            .O(N__6161),
            .I(\U712_CHIP_RAM.N_304 ));
    LocalMux I__987 (
            .O(N__6158),
            .I(\U712_CHIP_RAM.N_304 ));
    InMux I__986 (
            .O(N__6151),
            .I(N__6148));
    LocalMux I__985 (
            .O(N__6148),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__984 (
            .O(N__6145),
            .I(N__6142));
    LocalMux I__983 (
            .O(N__6142),
            .I(N__6137));
    InMux I__982 (
            .O(N__6141),
            .I(N__6132));
    InMux I__981 (
            .O(N__6140),
            .I(N__6132));
    Odrv4 I__980 (
            .O(N__6137),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__979 (
            .O(N__6132),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    IoInMux I__978 (
            .O(N__6127),
            .I(N__6124));
    LocalMux I__977 (
            .O(N__6124),
            .I(N__6120));
    IoInMux I__976 (
            .O(N__6123),
            .I(N__6117));
    IoSpan4Mux I__975 (
            .O(N__6120),
            .I(N__6114));
    LocalMux I__974 (
            .O(N__6117),
            .I(N__6110));
    Sp12to4 I__973 (
            .O(N__6114),
            .I(N__6107));
    IoInMux I__972 (
            .O(N__6113),
            .I(N__6104));
    Span4Mux_s1_h I__971 (
            .O(N__6110),
            .I(N__6101));
    Span12Mux_s7_v I__970 (
            .O(N__6107),
            .I(N__6098));
    LocalMux I__969 (
            .O(N__6104),
            .I(N__6095));
    Span4Mux_h I__968 (
            .O(N__6101),
            .I(N__6092));
    Span12Mux_h I__967 (
            .O(N__6098),
            .I(N__6089));
    Span12Mux_s7_v I__966 (
            .O(N__6095),
            .I(N__6086));
    Sp12to4 I__965 (
            .O(N__6092),
            .I(N__6083));
    Span12Mux_v I__964 (
            .O(N__6089),
            .I(N__6075));
    Span12Mux_v I__963 (
            .O(N__6086),
            .I(N__6075));
    Span12Mux_v I__962 (
            .O(N__6083),
            .I(N__6075));
    InMux I__961 (
            .O(N__6082),
            .I(N__6072));
    Odrv12 I__960 (
            .O(N__6075),
            .I(TACK_OUTn));
    LocalMux I__959 (
            .O(N__6072),
            .I(TACK_OUTn));
    InMux I__958 (
            .O(N__6067),
            .I(N__6064));
    LocalMux I__957 (
            .O(N__6064),
            .I(N__6061));
    Odrv4 I__956 (
            .O(N__6061),
            .I(\U712_REG_SM.N_404 ));
    IoInMux I__955 (
            .O(N__6058),
            .I(N__6055));
    LocalMux I__954 (
            .O(N__6055),
            .I(N__6052));
    IoSpan4Mux I__953 (
            .O(N__6052),
            .I(N__6049));
    Span4Mux_s0_v I__952 (
            .O(N__6049),
            .I(N__6046));
    Sp12to4 I__951 (
            .O(N__6046),
            .I(N__6043));
    Span12Mux_v I__950 (
            .O(N__6043),
            .I(N__6039));
    InMux I__949 (
            .O(N__6042),
            .I(N__6036));
    Odrv12 I__948 (
            .O(N__6039),
            .I(LDSn_c));
    LocalMux I__947 (
            .O(N__6036),
            .I(LDSn_c));
    IoInMux I__946 (
            .O(N__6031),
            .I(N__6028));
    LocalMux I__945 (
            .O(N__6028),
            .I(N__6025));
    IoSpan4Mux I__944 (
            .O(N__6025),
            .I(N__6022));
    Span4Mux_s3_h I__943 (
            .O(N__6022),
            .I(N__6019));
    Span4Mux_v I__942 (
            .O(N__6019),
            .I(N__6015));
    InMux I__941 (
            .O(N__6018),
            .I(N__6012));
    Span4Mux_h I__940 (
            .O(N__6015),
            .I(N__6009));
    LocalMux I__939 (
            .O(N__6012),
            .I(N__6006));
    Sp12to4 I__938 (
            .O(N__6009),
            .I(N__6003));
    Span4Mux_v I__937 (
            .O(N__6006),
            .I(N__6000));
    Span12Mux_h I__936 (
            .O(N__6003),
            .I(N__5995));
    Sp12to4 I__935 (
            .O(N__6000),
            .I(N__5995));
    Span12Mux_h I__934 (
            .O(N__5995),
            .I(N__5992));
    Odrv12 I__933 (
            .O(N__5992),
            .I(C3_c));
    InMux I__932 (
            .O(N__5989),
            .I(N__5986));
    LocalMux I__931 (
            .O(N__5986),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__930 (
            .O(N__5983),
            .I(N__5980));
    LocalMux I__929 (
            .O(N__5980),
            .I(\U712_REG_SM.N_459 ));
    IoInMux I__928 (
            .O(N__5977),
            .I(N__5974));
    LocalMux I__927 (
            .O(N__5974),
            .I(N__5971));
    IoSpan4Mux I__926 (
            .O(N__5971),
            .I(N__5968));
    IoSpan4Mux I__925 (
            .O(N__5968),
            .I(N__5965));
    Span4Mux_s3_v I__924 (
            .O(N__5965),
            .I(N__5962));
    Sp12to4 I__923 (
            .O(N__5962),
            .I(N__5958));
    CascadeMux I__922 (
            .O(N__5961),
            .I(N__5955));
    Span12Mux_s11_v I__921 (
            .O(N__5958),
            .I(N__5952));
    InMux I__920 (
            .O(N__5955),
            .I(N__5949));
    Odrv12 I__919 (
            .O(N__5952),
            .I(UDSn_c));
    LocalMux I__918 (
            .O(N__5949),
            .I(UDSn_c));
    InMux I__917 (
            .O(N__5944),
            .I(N__5941));
    LocalMux I__916 (
            .O(N__5941),
            .I(N__5935));
    CascadeMux I__915 (
            .O(N__5940),
            .I(N__5932));
    InMux I__914 (
            .O(N__5939),
            .I(N__5927));
    InMux I__913 (
            .O(N__5938),
            .I(N__5927));
    Span4Mux_h I__912 (
            .O(N__5935),
            .I(N__5924));
    InMux I__911 (
            .O(N__5932),
            .I(N__5921));
    LocalMux I__910 (
            .O(N__5927),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ));
    Odrv4 I__909 (
            .O(N__5924),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ));
    LocalMux I__908 (
            .O(N__5921),
            .I(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ));
    InMux I__907 (
            .O(N__5914),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_1 ));
    InMux I__906 (
            .O(N__5911),
            .I(\U712_CHIP_RAM.un3_DBR_COUNT_cry_2 ));
    InMux I__905 (
            .O(N__5908),
            .I(N__5902));
    InMux I__904 (
            .O(N__5907),
            .I(N__5902));
    LocalMux I__903 (
            .O(N__5902),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    CascadeMux I__902 (
            .O(N__5899),
            .I(\U712_REG_SM.N_410_cascade_ ));
    InMux I__901 (
            .O(N__5896),
            .I(N__5893));
    LocalMux I__900 (
            .O(N__5893),
            .I(\U712_REG_SM.N_331 ));
    InMux I__899 (
            .O(N__5890),
            .I(N__5886));
    IoInMux I__898 (
            .O(N__5889),
            .I(N__5883));
    LocalMux I__897 (
            .O(N__5886),
            .I(N__5880));
    LocalMux I__896 (
            .O(N__5883),
            .I(N__5877));
    Span4Mux_v I__895 (
            .O(N__5880),
            .I(N__5874));
    IoSpan4Mux I__894 (
            .O(N__5877),
            .I(N__5871));
    Sp12to4 I__893 (
            .O(N__5874),
            .I(N__5868));
    IoSpan4Mux I__892 (
            .O(N__5871),
            .I(N__5865));
    Span12Mux_h I__891 (
            .O(N__5868),
            .I(N__5862));
    IoSpan4Mux I__890 (
            .O(N__5865),
            .I(N__5859));
    Odrv12 I__889 (
            .O(N__5862),
            .I(C1_c));
    Odrv4 I__888 (
            .O(N__5859),
            .I(C1_c));
    InMux I__887 (
            .O(N__5854),
            .I(N__5848));
    InMux I__886 (
            .O(N__5853),
            .I(N__5848));
    LocalMux I__885 (
            .O(N__5848),
            .I(N__5845));
    Span4Mux_h I__884 (
            .O(N__5845),
            .I(N__5842));
    Odrv4 I__883 (
            .O(N__5842),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ));
    InMux I__882 (
            .O(N__5839),
            .I(N__5835));
    InMux I__881 (
            .O(N__5838),
            .I(N__5832));
    LocalMux I__880 (
            .O(N__5835),
            .I(\U712_CHIP_RAM.N_435 ));
    LocalMux I__879 (
            .O(N__5832),
            .I(\U712_CHIP_RAM.N_435 ));
    InMux I__878 (
            .O(N__5827),
            .I(N__5824));
    LocalMux I__877 (
            .O(N__5824),
            .I(N__5821));
    Odrv4 I__876 (
            .O(N__5821),
            .I(DBR_SYNCZ0Z_0));
    CascadeMux I__875 (
            .O(N__5818),
            .I(\U712_REG_SM.N_413_cascade_ ));
    IoInMux I__874 (
            .O(N__5815),
            .I(N__5812));
    LocalMux I__873 (
            .O(N__5812),
            .I(N__5809));
    Span4Mux_s3_v I__872 (
            .O(N__5809),
            .I(N__5806));
    Span4Mux_h I__871 (
            .O(N__5806),
            .I(N__5803));
    Sp12to4 I__870 (
            .O(N__5803),
            .I(N__5797));
    InMux I__869 (
            .O(N__5802),
            .I(N__5792));
    InMux I__868 (
            .O(N__5801),
            .I(N__5792));
    InMux I__867 (
            .O(N__5800),
            .I(N__5789));
    Odrv12 I__866 (
            .O(N__5797),
            .I(DBENn_c));
    LocalMux I__865 (
            .O(N__5792),
            .I(DBENn_c));
    LocalMux I__864 (
            .O(N__5789),
            .I(DBENn_c));
    InMux I__863 (
            .O(N__5782),
            .I(N__5776));
    InMux I__862 (
            .O(N__5781),
            .I(N__5776));
    LocalMux I__861 (
            .O(N__5776),
            .I(N__5773));
    Span4Mux_v I__860 (
            .O(N__5773),
            .I(N__5768));
    InMux I__859 (
            .O(N__5772),
            .I(N__5765));
    InMux I__858 (
            .O(N__5771),
            .I(N__5762));
    Odrv4 I__857 (
            .O(N__5768),
            .I(DMA_CYCLEm));
    LocalMux I__856 (
            .O(N__5765),
            .I(DMA_CYCLEm));
    LocalMux I__855 (
            .O(N__5762),
            .I(DMA_CYCLEm));
    InMux I__854 (
            .O(N__5755),
            .I(N__5752));
    LocalMux I__853 (
            .O(N__5752),
            .I(\U712_REG_SM.N_308 ));
    CascadeMux I__852 (
            .O(N__5749),
            .I(\U712_REG_SM.N_308_cascade_ ));
    CascadeMux I__851 (
            .O(N__5746),
            .I(N__5743));
    InMux I__850 (
            .O(N__5743),
            .I(N__5740));
    LocalMux I__849 (
            .O(N__5740),
            .I(\U712_CHIP_RAM.DBENn_7_0_0 ));
    InMux I__848 (
            .O(N__5737),
            .I(N__5734));
    LocalMux I__847 (
            .O(N__5734),
            .I(N__5728));
    InMux I__846 (
            .O(N__5733),
            .I(N__5724));
    CascadeMux I__845 (
            .O(N__5732),
            .I(N__5721));
    CascadeMux I__844 (
            .O(N__5731),
            .I(N__5718));
    Span4Mux_v I__843 (
            .O(N__5728),
            .I(N__5715));
    CascadeMux I__842 (
            .O(N__5727),
            .I(N__5711));
    LocalMux I__841 (
            .O(N__5724),
            .I(N__5708));
    InMux I__840 (
            .O(N__5721),
            .I(N__5703));
    InMux I__839 (
            .O(N__5718),
            .I(N__5699));
    Span4Mux_h I__838 (
            .O(N__5715),
            .I(N__5696));
    InMux I__837 (
            .O(N__5714),
            .I(N__5691));
    InMux I__836 (
            .O(N__5711),
            .I(N__5691));
    Span4Mux_h I__835 (
            .O(N__5708),
            .I(N__5688));
    InMux I__834 (
            .O(N__5707),
            .I(N__5683));
    InMux I__833 (
            .O(N__5706),
            .I(N__5683));
    LocalMux I__832 (
            .O(N__5703),
            .I(N__5680));
    InMux I__831 (
            .O(N__5702),
            .I(N__5677));
    LocalMux I__830 (
            .O(N__5699),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__829 (
            .O(N__5696),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__828 (
            .O(N__5691),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__827 (
            .O(N__5688),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__826 (
            .O(N__5683),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__825 (
            .O(N__5680),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__824 (
            .O(N__5677),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__823 (
            .O(N__5662),
            .I(N__5659));
    LocalMux I__822 (
            .O(N__5659),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1 ));
    CascadeMux I__821 (
            .O(N__5656),
            .I(\U712_CHIP_RAM.N_344_cascade_ ));
    InMux I__820 (
            .O(N__5653),
            .I(N__5648));
    InMux I__819 (
            .O(N__5652),
            .I(N__5645));
    InMux I__818 (
            .O(N__5651),
            .I(N__5642));
    LocalMux I__817 (
            .O(N__5648),
            .I(\U712_CHIP_RAM.N_551 ));
    LocalMux I__816 (
            .O(N__5645),
            .I(\U712_CHIP_RAM.N_551 ));
    LocalMux I__815 (
            .O(N__5642),
            .I(\U712_CHIP_RAM.N_551 ));
    CascadeMux I__814 (
            .O(N__5635),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_2_0_cascade_ ));
    InMux I__813 (
            .O(N__5632),
            .I(N__5629));
    LocalMux I__812 (
            .O(N__5629),
            .I(\U712_CHIP_RAM.LATCH_CLK_6 ));
    IoInMux I__811 (
            .O(N__5626),
            .I(N__5623));
    LocalMux I__810 (
            .O(N__5623),
            .I(N__5620));
    IoSpan4Mux I__809 (
            .O(N__5620),
            .I(N__5617));
    Span4Mux_s3_v I__808 (
            .O(N__5617),
            .I(N__5614));
    Span4Mux_v I__807 (
            .O(N__5614),
            .I(N__5611));
    Sp12to4 I__806 (
            .O(N__5611),
            .I(N__5608));
    Span12Mux_v I__805 (
            .O(N__5608),
            .I(N__5604));
    InMux I__804 (
            .O(N__5607),
            .I(N__5601));
    Odrv12 I__803 (
            .O(N__5604),
            .I(LATCH_CLK_c));
    LocalMux I__802 (
            .O(N__5601),
            .I(LATCH_CLK_c));
    InMux I__801 (
            .O(N__5596),
            .I(N__5590));
    InMux I__800 (
            .O(N__5595),
            .I(N__5590));
    LocalMux I__799 (
            .O(N__5590),
            .I(N__5586));
    InMux I__798 (
            .O(N__5589),
            .I(N__5583));
    Span4Mux_h I__797 (
            .O(N__5586),
            .I(N__5580));
    LocalMux I__796 (
            .O(N__5583),
            .I(N__5577));
    Span4Mux_v I__795 (
            .O(N__5580),
            .I(N__5572));
    Span4Mux_v I__794 (
            .O(N__5577),
            .I(N__5572));
    Span4Mux_h I__793 (
            .O(N__5572),
            .I(N__5569));
    Sp12to4 I__792 (
            .O(N__5569),
            .I(N__5566));
    Odrv12 I__791 (
            .O(N__5566),
            .I(AWEn_c));
    InMux I__790 (
            .O(N__5563),
            .I(N__5559));
    InMux I__789 (
            .O(N__5562),
            .I(N__5556));
    LocalMux I__788 (
            .O(N__5559),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    LocalMux I__787 (
            .O(N__5556),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    InMux I__786 (
            .O(N__5551),
            .I(N__5548));
    LocalMux I__785 (
            .O(N__5548),
            .I(N__5545));
    Sp12to4 I__784 (
            .O(N__5545),
            .I(N__5542));
    Span12Mux_v I__783 (
            .O(N__5542),
            .I(N__5539));
    Span12Mux_h I__782 (
            .O(N__5539),
            .I(N__5536));
    Odrv12 I__781 (
            .O(N__5536),
            .I(A_c_20));
    InMux I__780 (
            .O(N__5533),
            .I(N__5529));
    InMux I__779 (
            .O(N__5532),
            .I(N__5526));
    LocalMux I__778 (
            .O(N__5529),
            .I(N__5523));
    LocalMux I__777 (
            .O(N__5526),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    Odrv12 I__776 (
            .O(N__5523),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    InMux I__775 (
            .O(N__5518),
            .I(N__5515));
    LocalMux I__774 (
            .O(N__5515),
            .I(N__5510));
    InMux I__773 (
            .O(N__5514),
            .I(N__5507));
    InMux I__772 (
            .O(N__5513),
            .I(N__5504));
    Odrv4 I__771 (
            .O(N__5510),
            .I(\U712_CHIP_RAM.N_194 ));
    LocalMux I__770 (
            .O(N__5507),
            .I(\U712_CHIP_RAM.N_194 ));
    LocalMux I__769 (
            .O(N__5504),
            .I(\U712_CHIP_RAM.N_194 ));
    CascadeMux I__768 (
            .O(N__5497),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_2_2_cascade_ ));
    InMux I__767 (
            .O(N__5494),
            .I(N__5491));
    LocalMux I__766 (
            .O(N__5491),
            .I(\U712_CHIP_RAM.N_449 ));
    InMux I__765 (
            .O(N__5488),
            .I(N__5485));
    LocalMux I__764 (
            .O(N__5485),
            .I(N__5481));
    InMux I__763 (
            .O(N__5484),
            .I(N__5478));
    Span4Mux_h I__762 (
            .O(N__5481),
            .I(N__5475));
    LocalMux I__761 (
            .O(N__5478),
            .I(\U712_CHIP_RAM.N_476 ));
    Odrv4 I__760 (
            .O(N__5475),
            .I(\U712_CHIP_RAM.N_476 ));
    InMux I__759 (
            .O(N__5470),
            .I(N__5467));
    LocalMux I__758 (
            .O(N__5467),
            .I(N__5464));
    Span4Mux_v I__757 (
            .O(N__5464),
            .I(N__5460));
    InMux I__756 (
            .O(N__5463),
            .I(N__5457));
    Odrv4 I__755 (
            .O(N__5460),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ));
    LocalMux I__754 (
            .O(N__5457),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ));
    InMux I__753 (
            .O(N__5452),
            .I(N__5449));
    LocalMux I__752 (
            .O(N__5449),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    CascadeMux I__751 (
            .O(N__5446),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_ ));
    CascadeMux I__750 (
            .O(N__5443),
            .I(\U712_CHIP_RAM.N_304_cascade_ ));
    CascadeMux I__749 (
            .O(N__5440),
            .I(\U712_CHIP_RAM.N_312_cascade_ ));
    CascadeMux I__748 (
            .O(N__5437),
            .I(\U712_CHIP_RAM.N_326_cascade_ ));
    InMux I__747 (
            .O(N__5434),
            .I(N__5431));
    LocalMux I__746 (
            .O(N__5431),
            .I(N__5427));
    InMux I__745 (
            .O(N__5430),
            .I(N__5424));
    Span4Mux_v I__744 (
            .O(N__5427),
            .I(N__5417));
    LocalMux I__743 (
            .O(N__5424),
            .I(N__5414));
    InMux I__742 (
            .O(N__5423),
            .I(N__5407));
    InMux I__741 (
            .O(N__5422),
            .I(N__5407));
    InMux I__740 (
            .O(N__5421),
            .I(N__5407));
    InMux I__739 (
            .O(N__5420),
            .I(N__5404));
    Odrv4 I__738 (
            .O(N__5417),
            .I(\U712_CHIP_RAM.N_467 ));
    Odrv4 I__737 (
            .O(N__5414),
            .I(\U712_CHIP_RAM.N_467 ));
    LocalMux I__736 (
            .O(N__5407),
            .I(\U712_CHIP_RAM.N_467 ));
    LocalMux I__735 (
            .O(N__5404),
            .I(\U712_CHIP_RAM.N_467 ));
    InMux I__734 (
            .O(N__5395),
            .I(N__5386));
    InMux I__733 (
            .O(N__5394),
            .I(N__5386));
    InMux I__732 (
            .O(N__5393),
            .I(N__5386));
    LocalMux I__731 (
            .O(N__5386),
            .I(N__5379));
    InMux I__730 (
            .O(N__5385),
            .I(N__5376));
    InMux I__729 (
            .O(N__5384),
            .I(N__5369));
    InMux I__728 (
            .O(N__5383),
            .I(N__5369));
    InMux I__727 (
            .O(N__5382),
            .I(N__5369));
    Odrv4 I__726 (
            .O(N__5379),
            .I(\U712_CHIP_RAM.N_39 ));
    LocalMux I__725 (
            .O(N__5376),
            .I(\U712_CHIP_RAM.N_39 ));
    LocalMux I__724 (
            .O(N__5369),
            .I(\U712_CHIP_RAM.N_39 ));
    InMux I__723 (
            .O(N__5362),
            .I(N__5359));
    LocalMux I__722 (
            .O(N__5359),
            .I(N__5356));
    Odrv4 I__721 (
            .O(N__5356),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    InMux I__720 (
            .O(N__5353),
            .I(N__5350));
    LocalMux I__719 (
            .O(N__5350),
            .I(N__5347));
    Odrv12 I__718 (
            .O(N__5347),
            .I(\U712_CHIP_RAM.N_440 ));
    CascadeMux I__717 (
            .O(N__5344),
            .I(\U712_CHIP_RAM.N_39_cascade_ ));
    InMux I__716 (
            .O(N__5341),
            .I(N__5338));
    LocalMux I__715 (
            .O(N__5338),
            .I(\U712_CHIP_RAM.N_326 ));
    CEMux I__714 (
            .O(N__5335),
            .I(N__5332));
    LocalMux I__713 (
            .O(N__5332),
            .I(N__5328));
    CEMux I__712 (
            .O(N__5331),
            .I(N__5325));
    Span4Mux_h I__711 (
            .O(N__5328),
            .I(N__5322));
    LocalMux I__710 (
            .O(N__5325),
            .I(N__5319));
    Odrv4 I__709 (
            .O(N__5322),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    Odrv12 I__708 (
            .O(N__5319),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__707 (
            .O(N__5314),
            .I(N__5311));
    LocalMux I__706 (
            .O(N__5311),
            .I(N__5308));
    Span4Mux_v I__705 (
            .O(N__5308),
            .I(N__5305));
    Span4Mux_v I__704 (
            .O(N__5305),
            .I(N__5302));
    Sp12to4 I__703 (
            .O(N__5302),
            .I(N__5299));
    Odrv12 I__702 (
            .O(N__5299),
            .I(A_c_17));
    CascadeMux I__701 (
            .O(N__5296),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ));
    InMux I__700 (
            .O(N__5293),
            .I(N__5290));
    LocalMux I__699 (
            .O(N__5290),
            .I(N__5287));
    Sp12to4 I__698 (
            .O(N__5287),
            .I(N__5284));
    Span12Mux_v I__697 (
            .O(N__5284),
            .I(N__5281));
    Span12Mux_h I__696 (
            .O(N__5281),
            .I(N__5278));
    Odrv12 I__695 (
            .O(N__5278),
            .I(A_c_18));
    InMux I__694 (
            .O(N__5275),
            .I(N__5272));
    LocalMux I__693 (
            .O(N__5272),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ));
    CascadeMux I__692 (
            .O(N__5269),
            .I(N__5266));
    InMux I__691 (
            .O(N__5266),
            .I(N__5263));
    LocalMux I__690 (
            .O(N__5263),
            .I(N__5260));
    Odrv4 I__689 (
            .O(N__5260),
            .I(\U712_CHIP_RAM.N_555 ));
    CascadeMux I__688 (
            .O(N__5257),
            .I(\U712_CHIP_RAM.N_555_cascade_ ));
    InMux I__687 (
            .O(N__5254),
            .I(N__5251));
    LocalMux I__686 (
            .O(N__5251),
            .I(\U712_REG_SM.N_412 ));
    InMux I__685 (
            .O(N__5248),
            .I(N__5245));
    LocalMux I__684 (
            .O(N__5245),
            .I(N__5242));
    Odrv12 I__683 (
            .O(N__5242),
            .I(\U712_REG_SM.N_402 ));
    InMux I__682 (
            .O(N__5239),
            .I(N__5235));
    InMux I__681 (
            .O(N__5238),
            .I(N__5232));
    LocalMux I__680 (
            .O(N__5235),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    LocalMux I__679 (
            .O(N__5232),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    IoInMux I__678 (
            .O(N__5227),
            .I(N__5224));
    LocalMux I__677 (
            .O(N__5224),
            .I(N__5221));
    Span4Mux_s3_v I__676 (
            .O(N__5221),
            .I(N__5218));
    Sp12to4 I__675 (
            .O(N__5218),
            .I(N__5215));
    Span12Mux_s9_h I__674 (
            .O(N__5215),
            .I(N__5210));
    CascadeMux I__673 (
            .O(N__5214),
            .I(N__5207));
    InMux I__672 (
            .O(N__5213),
            .I(N__5204));
    Span12Mux_v I__671 (
            .O(N__5210),
            .I(N__5201));
    InMux I__670 (
            .O(N__5207),
            .I(N__5198));
    LocalMux I__669 (
            .O(N__5204),
            .I(N__5195));
    Odrv12 I__668 (
            .O(N__5201),
            .I(REGENn_c));
    LocalMux I__667 (
            .O(N__5198),
            .I(REGENn_c));
    Odrv4 I__666 (
            .O(N__5195),
            .I(REGENn_c));
    CascadeMux I__665 (
            .O(N__5188),
            .I(N__5184));
    InMux I__664 (
            .O(N__5187),
            .I(N__5179));
    InMux I__663 (
            .O(N__5184),
            .I(N__5172));
    InMux I__662 (
            .O(N__5183),
            .I(N__5172));
    InMux I__661 (
            .O(N__5182),
            .I(N__5172));
    LocalMux I__660 (
            .O(N__5179),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__659 (
            .O(N__5172),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__658 (
            .O(N__5167),
            .I(N__5164));
    LocalMux I__657 (
            .O(N__5164),
            .I(N__5161));
    Odrv4 I__656 (
            .O(N__5161),
            .I(\U712_REG_SM.REGENn_e_1 ));
    InMux I__655 (
            .O(N__5158),
            .I(N__5155));
    LocalMux I__654 (
            .O(N__5155),
            .I(N__5152));
    Sp12to4 I__653 (
            .O(N__5152),
            .I(N__5149));
    Span12Mux_v I__652 (
            .O(N__5149),
            .I(N__5146));
    Span12Mux_h I__651 (
            .O(N__5146),
            .I(N__5143));
    Odrv12 I__650 (
            .O(N__5143),
            .I(A_c_16));
    CascadeMux I__649 (
            .O(N__5140),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_cascade_ ));
    InMux I__648 (
            .O(N__5137),
            .I(N__5134));
    LocalMux I__647 (
            .O(N__5134),
            .I(N__5131));
    Odrv12 I__646 (
            .O(N__5131),
            .I(\U712_CHIP_RAM.N_378 ));
    CascadeMux I__645 (
            .O(N__5128),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ));
    CascadeMux I__644 (
            .O(N__5125),
            .I(\U712_CHIP_RAM.N_551_cascade_ ));
    InMux I__643 (
            .O(N__5122),
            .I(N__5119));
    LocalMux I__642 (
            .O(N__5119),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a3_0_a2_0 ));
    IoInMux I__641 (
            .O(N__5116),
            .I(N__5113));
    LocalMux I__640 (
            .O(N__5113),
            .I(N__5110));
    Span4Mux_s0_h I__639 (
            .O(N__5110),
            .I(N__5107));
    Sp12to4 I__638 (
            .O(N__5107),
            .I(N__5104));
    Span12Mux_v I__637 (
            .O(N__5104),
            .I(N__5101));
    Span12Mux_h I__636 (
            .O(N__5101),
            .I(N__5097));
    InMux I__635 (
            .O(N__5100),
            .I(N__5094));
    Odrv12 I__634 (
            .O(N__5097),
            .I(CLK_EN_c));
    LocalMux I__633 (
            .O(N__5094),
            .I(CLK_EN_c));
    InMux I__632 (
            .O(N__5089),
            .I(N__5085));
    InMux I__631 (
            .O(N__5088),
            .I(N__5082));
    LocalMux I__630 (
            .O(N__5085),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0 ));
    LocalMux I__629 (
            .O(N__5082),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0 ));
    IoInMux I__628 (
            .O(N__5077),
            .I(N__5074));
    LocalMux I__627 (
            .O(N__5074),
            .I(N__5071));
    Span4Mux_s3_v I__626 (
            .O(N__5071),
            .I(N__5068));
    Span4Mux_v I__625 (
            .O(N__5068),
            .I(N__5065));
    Span4Mux_v I__624 (
            .O(N__5065),
            .I(N__5062));
    Span4Mux_v I__623 (
            .O(N__5062),
            .I(N__5058));
    InMux I__622 (
            .O(N__5061),
            .I(N__5055));
    Odrv4 I__621 (
            .O(N__5058),
            .I(DBDIR_c));
    LocalMux I__620 (
            .O(N__5055),
            .I(DBDIR_c));
    InMux I__619 (
            .O(N__5050),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__618 (
            .O(N__5047),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__617 (
            .O(N__5044),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__616 (
            .O(N__5041),
            .I(N__5034));
    InMux I__615 (
            .O(N__5040),
            .I(N__5034));
    InMux I__614 (
            .O(N__5039),
            .I(N__5029));
    LocalMux I__613 (
            .O(N__5034),
            .I(N__5026));
    InMux I__612 (
            .O(N__5033),
            .I(N__5023));
    InMux I__611 (
            .O(N__5032),
            .I(N__5020));
    LocalMux I__610 (
            .O(N__5029),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    Odrv4 I__609 (
            .O(N__5026),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__608 (
            .O(N__5023),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__607 (
            .O(N__5020),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__606 (
            .O(N__5011),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__605 (
            .O(N__5008),
            .I(N__5003));
    CascadeMux I__604 (
            .O(N__5007),
            .I(N__5000));
    InMux I__603 (
            .O(N__5006),
            .I(N__4997));
    LocalMux I__602 (
            .O(N__5003),
            .I(N__4994));
    InMux I__601 (
            .O(N__5000),
            .I(N__4991));
    LocalMux I__600 (
            .O(N__4997),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    Odrv4 I__599 (
            .O(N__4994),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__598 (
            .O(N__4991),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__597 (
            .O(N__4984),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    CascadeMux I__596 (
            .O(N__4981),
            .I(N__4978));
    InMux I__595 (
            .O(N__4978),
            .I(N__4975));
    LocalMux I__594 (
            .O(N__4975),
            .I(N__4969));
    InMux I__593 (
            .O(N__4974),
            .I(N__4966));
    InMux I__592 (
            .O(N__4973),
            .I(N__4962));
    InMux I__591 (
            .O(N__4972),
            .I(N__4959));
    Sp12to4 I__590 (
            .O(N__4969),
            .I(N__4954));
    LocalMux I__589 (
            .O(N__4966),
            .I(N__4954));
    InMux I__588 (
            .O(N__4965),
            .I(N__4951));
    LocalMux I__587 (
            .O(N__4962),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__586 (
            .O(N__4959),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    Odrv12 I__585 (
            .O(N__4954),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__584 (
            .O(N__4951),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__583 (
            .O(N__4942),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__582 (
            .O(N__4939),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    InMux I__581 (
            .O(N__4936),
            .I(N__4932));
    InMux I__580 (
            .O(N__4935),
            .I(N__4929));
    LocalMux I__579 (
            .O(N__4932),
            .I(N__4925));
    LocalMux I__578 (
            .O(N__4929),
            .I(N__4922));
    InMux I__577 (
            .O(N__4928),
            .I(N__4919));
    Odrv4 I__576 (
            .O(N__4925),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    Odrv4 I__575 (
            .O(N__4922),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__574 (
            .O(N__4919),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__573 (
            .O(N__4912),
            .I(N__4909));
    LocalMux I__572 (
            .O(N__4909),
            .I(N__4906));
    Odrv4 I__571 (
            .O(N__4906),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_1 ));
    CascadeMux I__570 (
            .O(N__4903),
            .I(\U712_CHIP_RAM.N_305_cascade_ ));
    CascadeMux I__569 (
            .O(N__4900),
            .I(N__4896));
    CascadeMux I__568 (
            .O(N__4899),
            .I(N__4893));
    InMux I__567 (
            .O(N__4896),
            .I(N__4887));
    InMux I__566 (
            .O(N__4893),
            .I(N__4887));
    InMux I__565 (
            .O(N__4892),
            .I(N__4884));
    LocalMux I__564 (
            .O(N__4887),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__563 (
            .O(N__4884),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__562 (
            .O(N__4879),
            .I(N__4876));
    InMux I__561 (
            .O(N__4876),
            .I(N__4873));
    LocalMux I__560 (
            .O(N__4873),
            .I(N__4868));
    InMux I__559 (
            .O(N__4872),
            .I(N__4865));
    InMux I__558 (
            .O(N__4871),
            .I(N__4862));
    Odrv4 I__557 (
            .O(N__4868),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__556 (
            .O(N__4865),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__555 (
            .O(N__4862),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__554 (
            .O(N__4855),
            .I(N__4850));
    InMux I__553 (
            .O(N__4854),
            .I(N__4847));
    InMux I__552 (
            .O(N__4853),
            .I(N__4844));
    LocalMux I__551 (
            .O(N__4850),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    LocalMux I__550 (
            .O(N__4847),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    LocalMux I__549 (
            .O(N__4844),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    InMux I__548 (
            .O(N__4837),
            .I(N__4834));
    LocalMux I__547 (
            .O(N__4834),
            .I(\U712_CHIP_RAM.N_325 ));
    CascadeMux I__546 (
            .O(N__4831),
            .I(\U712_CHIP_RAM.N_325_cascade_ ));
    CascadeMux I__545 (
            .O(N__4828),
            .I(\U712_CHIP_RAM.m101_i_0_cascade_ ));
    InMux I__544 (
            .O(N__4825),
            .I(N__4822));
    LocalMux I__543 (
            .O(N__4822),
            .I(\U712_CHIP_RAM.m101_i_1 ));
    InMux I__542 (
            .O(N__4819),
            .I(N__4816));
    LocalMux I__541 (
            .O(N__4816),
            .I(\U712_CHIP_RAM.N_376 ));
    CascadeMux I__540 (
            .O(N__4813),
            .I(\U712_CHIP_RAM.m101_i_2_cascade_ ));
    InMux I__539 (
            .O(N__4810),
            .I(N__4807));
    LocalMux I__538 (
            .O(N__4807),
            .I(\U712_CHIP_RAM.N_436 ));
    CascadeMux I__537 (
            .O(N__4804),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_ ));
    CascadeMux I__536 (
            .O(N__4801),
            .I(N__4798));
    InMux I__535 (
            .O(N__4798),
            .I(N__4789));
    InMux I__534 (
            .O(N__4797),
            .I(N__4789));
    InMux I__533 (
            .O(N__4796),
            .I(N__4789));
    LocalMux I__532 (
            .O(N__4789),
            .I(\U712_CHIP_RAM.SDRAM_CMDs_0_4 ));
    CascadeMux I__531 (
            .O(N__4786),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_ ));
    CascadeMux I__530 (
            .O(N__4783),
            .I(\U712_CHIP_RAM.N_396_cascade_ ));
    InMux I__529 (
            .O(N__4780),
            .I(N__4777));
    LocalMux I__528 (
            .O(N__4777),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_0_2 ));
    InMux I__527 (
            .O(N__4774),
            .I(N__4771));
    LocalMux I__526 (
            .O(N__4771),
            .I(\U712_CHIP_RAM.N_397 ));
    InMux I__525 (
            .O(N__4768),
            .I(N__4765));
    LocalMux I__524 (
            .O(N__4765),
            .I(\U712_CHIP_RAM.SDRAM_CMDsr_1_3 ));
    InMux I__523 (
            .O(N__4762),
            .I(N__4756));
    InMux I__522 (
            .O(N__4761),
            .I(N__4756));
    LocalMux I__521 (
            .O(N__4756),
            .I(N__4753));
    Odrv4 I__520 (
            .O(N__4753),
            .I(\U712_CHIP_RAM.SDRAM_CMDs_0_1 ));
    CEMux I__519 (
            .O(N__4750),
            .I(N__4747));
    LocalMux I__518 (
            .O(N__4747),
            .I(N__4744));
    Span4Mux_v I__517 (
            .O(N__4744),
            .I(N__4741));
    Span4Mux_h I__516 (
            .O(N__4741),
            .I(N__4738));
    Odrv4 I__515 (
            .O(N__4738),
            .I(\U712_CHIP_RAM.N_194_0 ));
    InMux I__514 (
            .O(N__4735),
            .I(N__4729));
    InMux I__513 (
            .O(N__4734),
            .I(N__4729));
    LocalMux I__512 (
            .O(N__4729),
            .I(N__4726));
    Odrv4 I__511 (
            .O(N__4726),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ));
    CEMux I__510 (
            .O(N__4723),
            .I(N__4720));
    LocalMux I__509 (
            .O(N__4720),
            .I(N__4717));
    Odrv4 I__508 (
            .O(N__4717),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0 ));
    InMux I__507 (
            .O(N__4714),
            .I(N__4710));
    InMux I__506 (
            .O(N__4713),
            .I(N__4707));
    LocalMux I__505 (
            .O(N__4710),
            .I(N__4704));
    LocalMux I__504 (
            .O(N__4707),
            .I(N__4701));
    Span4Mux_v I__503 (
            .O(N__4704),
            .I(N__4698));
    Span4Mux_v I__502 (
            .O(N__4701),
            .I(N__4695));
    Sp12to4 I__501 (
            .O(N__4698),
            .I(N__4692));
    Span4Mux_h I__500 (
            .O(N__4695),
            .I(N__4689));
    Span12Mux_h I__499 (
            .O(N__4692),
            .I(N__4684));
    Sp12to4 I__498 (
            .O(N__4689),
            .I(N__4684));
    Span12Mux_v I__497 (
            .O(N__4684),
            .I(N__4681));
    Odrv12 I__496 (
            .O(N__4681),
            .I(DBRn_c));
    InMux I__495 (
            .O(N__4678),
            .I(N__4675));
    LocalMux I__494 (
            .O(N__4675),
            .I(N__4671));
    InMux I__493 (
            .O(N__4674),
            .I(N__4668));
    Span4Mux_v I__492 (
            .O(N__4671),
            .I(N__4663));
    LocalMux I__491 (
            .O(N__4668),
            .I(N__4663));
    Span4Mux_v I__490 (
            .O(N__4663),
            .I(N__4660));
    Span4Mux_v I__489 (
            .O(N__4660),
            .I(N__4657));
    Span4Mux_h I__488 (
            .O(N__4657),
            .I(N__4654));
    Odrv4 I__487 (
            .O(N__4654),
            .I(TSn_c));
    InMux I__486 (
            .O(N__4651),
            .I(N__4648));
    LocalMux I__485 (
            .O(N__4648),
            .I(N__4645));
    Span12Mux_v I__484 (
            .O(N__4645),
            .I(N__4642));
    Odrv12 I__483 (
            .O(N__4642),
            .I(RAMSPACEn_c));
    InMux I__482 (
            .O(N__4639),
            .I(N__4636));
    LocalMux I__481 (
            .O(N__4636),
            .I(N__4633));
    Span12Mux_v I__480 (
            .O(N__4633),
            .I(N__4630));
    Odrv12 I__479 (
            .O(N__4630),
            .I(\U712_CHIP_RAM.N_419 ));
    IoInMux I__478 (
            .O(N__4627),
            .I(N__4624));
    LocalMux I__477 (
            .O(N__4624),
            .I(N__4621));
    Odrv12 I__476 (
            .O(N__4621),
            .I(VBENn_c));
    InMux I__475 (
            .O(N__4618),
            .I(N__4615));
    LocalMux I__474 (
            .O(N__4615),
            .I(\U712_CHIP_RAM.N_428 ));
    CascadeMux I__473 (
            .O(N__4612),
            .I(\U712_CHIP_RAM.N_307_cascade_ ));
    CascadeMux I__472 (
            .O(N__4609),
            .I(\U712_CHIP_RAM.N_467_cascade_ ));
    CascadeMux I__471 (
            .O(N__4606),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ));
    InMux I__470 (
            .O(N__4603),
            .I(N__4599));
    InMux I__469 (
            .O(N__4602),
            .I(N__4596));
    LocalMux I__468 (
            .O(N__4599),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__467 (
            .O(N__4596),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__466 (
            .O(N__4591),
            .I(N__4587));
    InMux I__465 (
            .O(N__4590),
            .I(N__4584));
    LocalMux I__464 (
            .O(N__4587),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__463 (
            .O(N__4584),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__462 (
            .O(N__4579),
            .I(N__4575));
    InMux I__461 (
            .O(N__4578),
            .I(N__4572));
    LocalMux I__460 (
            .O(N__4575),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__459 (
            .O(N__4572),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    CascadeMux I__458 (
            .O(N__4567),
            .I(\U712_CHIP_RAM.REFRESH5lto7_0_cascade_ ));
    InMux I__457 (
            .O(N__4564),
            .I(N__4560));
    InMux I__456 (
            .O(N__4563),
            .I(N__4557));
    LocalMux I__455 (
            .O(N__4560),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__454 (
            .O(N__4557),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__453 (
            .O(N__4552),
            .I(N__4548));
    InMux I__452 (
            .O(N__4551),
            .I(N__4545));
    LocalMux I__451 (
            .O(N__4548),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__450 (
            .O(N__4545),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    CascadeMux I__449 (
            .O(N__4540),
            .I(N__4536));
    InMux I__448 (
            .O(N__4539),
            .I(N__4533));
    InMux I__447 (
            .O(N__4536),
            .I(N__4530));
    LocalMux I__446 (
            .O(N__4533),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__445 (
            .O(N__4530),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__444 (
            .O(N__4525),
            .I(N__4521));
    InMux I__443 (
            .O(N__4524),
            .I(N__4518));
    LocalMux I__442 (
            .O(N__4521),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__441 (
            .O(N__4518),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__440 (
            .O(N__4513),
            .I(N__4510));
    LocalMux I__439 (
            .O(N__4510),
            .I(\U712_CHIP_RAM.REFRESH5lt7 ));
    CascadeMux I__438 (
            .O(N__4507),
            .I(\U712_CHIP_RAM.N_430_cascade_ ));
    InMux I__437 (
            .O(N__4504),
            .I(N__4501));
    LocalMux I__436 (
            .O(N__4501),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ));
    InMux I__435 (
            .O(N__4498),
            .I(N__4495));
    LocalMux I__434 (
            .O(N__4495),
            .I(N__4492));
    Span4Mux_h I__433 (
            .O(N__4492),
            .I(N__4489));
    Sp12to4 I__432 (
            .O(N__4489),
            .I(N__4486));
    Span12Mux_v I__431 (
            .O(N__4486),
            .I(N__4483));
    Odrv12 I__430 (
            .O(N__4483),
            .I(A_c_2));
    InMux I__429 (
            .O(N__4480),
            .I(N__4477));
    LocalMux I__428 (
            .O(N__4477),
            .I(N__4474));
    Span12Mux_v I__427 (
            .O(N__4474),
            .I(N__4471));
    Odrv12 I__426 (
            .O(N__4471),
            .I(A_c_4));
    InMux I__425 (
            .O(N__4468),
            .I(N__4465));
    LocalMux I__424 (
            .O(N__4465),
            .I(N__4462));
    Span4Mux_v I__423 (
            .O(N__4462),
            .I(N__4459));
    Span4Mux_v I__422 (
            .O(N__4459),
            .I(N__4456));
    Sp12to4 I__421 (
            .O(N__4456),
            .I(N__4453));
    Odrv12 I__420 (
            .O(N__4453),
            .I(A_c_7));
    InMux I__419 (
            .O(N__4450),
            .I(N__4447));
    LocalMux I__418 (
            .O(N__4447),
            .I(N__4444));
    Span12Mux_v I__417 (
            .O(N__4444),
            .I(N__4441));
    Odrv12 I__416 (
            .O(N__4441),
            .I(A_c_8));
    InMux I__415 (
            .O(N__4438),
            .I(N__4435));
    LocalMux I__414 (
            .O(N__4435),
            .I(N__4432));
    Span12Mux_h I__413 (
            .O(N__4432),
            .I(N__4429));
    Span12Mux_v I__412 (
            .O(N__4429),
            .I(N__4426));
    Odrv12 I__411 (
            .O(N__4426),
            .I(REGSPACEn_c));
    CascadeMux I__410 (
            .O(N__4423),
            .I(\U712_CHIP_RAM.m93_i_a2_4_cascade_ ));
    IoInMux I__409 (
            .O(N__4420),
            .I(N__4417));
    LocalMux I__408 (
            .O(N__4417),
            .I(N__4414));
    Span4Mux_s2_v I__407 (
            .O(N__4414),
            .I(N__4411));
    Span4Mux_v I__406 (
            .O(N__4411),
            .I(N__4408));
    Span4Mux_h I__405 (
            .O(N__4408),
            .I(N__4405));
    Odrv4 I__404 (
            .O(N__4405),
            .I(CLK80_PLL_i_i));
    InMux I__403 (
            .O(N__4402),
            .I(N__4399));
    LocalMux I__402 (
            .O(N__4399),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__401 (
            .O(N__4396),
            .I(bfn_6_6_0_));
    InMux I__400 (
            .O(N__4393),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__399 (
            .O(N__4390),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__398 (
            .O(N__4387),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__397 (
            .O(N__4384),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__396 (
            .O(N__4381),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__395 (
            .O(N__4378),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__394 (
            .O(N__4375),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__393 (
            .O(N__4372),
            .I(N__4348));
    ClkMux I__392 (
            .O(N__4371),
            .I(N__4348));
    ClkMux I__391 (
            .O(N__4370),
            .I(N__4348));
    ClkMux I__390 (
            .O(N__4369),
            .I(N__4348));
    ClkMux I__389 (
            .O(N__4368),
            .I(N__4348));
    ClkMux I__388 (
            .O(N__4367),
            .I(N__4348));
    ClkMux I__387 (
            .O(N__4366),
            .I(N__4348));
    ClkMux I__386 (
            .O(N__4365),
            .I(N__4348));
    GlobalMux I__385 (
            .O(N__4348),
            .I(N__4345));
    gio2CtrlBuf I__384 (
            .O(N__4345),
            .I(C1_c_g));
    IoInMux I__383 (
            .O(N__4342),
            .I(N__4339));
    LocalMux I__382 (
            .O(N__4339),
            .I(N__4336));
    Span12Mux_s4_h I__381 (
            .O(N__4336),
            .I(N__4333));
    Odrv12 I__380 (
            .O(N__4333),
            .I(DBRn_c_i_0));
    IoInMux I__379 (
            .O(N__4330),
            .I(N__4327));
    LocalMux I__378 (
            .O(N__4327),
            .I(N__4324));
    Span4Mux_s0_v I__377 (
            .O(N__4324),
            .I(N__4321));
    Span4Mux_v I__376 (
            .O(N__4321),
            .I(N__4318));
    Sp12to4 I__375 (
            .O(N__4318),
            .I(N__4315));
    Span12Mux_h I__374 (
            .O(N__4315),
            .I(N__4312));
    Span12Mux_v I__373 (
            .O(N__4312),
            .I(N__4309));
    Odrv12 I__372 (
            .O(N__4309),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .I(N__4371));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__4365));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__4366));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__4369));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__4368));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .I(N__4367));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__4370));
    defparam IN_MUX_bfv_10_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_5_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__5889),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__9592),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4342),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__6031),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_10_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_1_10_1  (
            .in0(N__8220),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10567),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_5_1_6.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_5_1_6.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_5_1_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_5_1_6 (
            .in0(N__9973),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_6_6_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_6_6_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_6_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__4402),
            .in2(_gnd_net_),
            .in3(N__4396),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__4372),
            .ce(),
            .sr(N__6190));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_6_6_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_6_6_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_6_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__4525),
            .in2(_gnd_net_),
            .in3(N__4393),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__4372),
            .ce(),
            .sr(N__6190));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_6_6_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_6_6_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_6_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__4552),
            .in2(_gnd_net_),
            .in3(N__4390),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__4372),
            .ce(),
            .sr(N__6190));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_6_6_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_6_6_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_6_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__4564),
            .in2(_gnd_net_),
            .in3(N__4387),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__4372),
            .ce(),
            .sr(N__6190));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_6_6_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_6_6_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_6_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__4539),
            .in2(_gnd_net_),
            .in3(N__4384),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__4372),
            .ce(),
            .sr(N__6190));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_6_6_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_6_6_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_6_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_6_6_5  (
            .in0(_gnd_net_),
            .in1(N__4591),
            .in2(_gnd_net_),
            .in3(N__4381),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__4372),
            .ce(),
            .sr(N__6190));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_6_6_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_6_6_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_6_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(N__4603),
            .in2(_gnd_net_),
            .in3(N__4378),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__4372),
            .ce(),
            .sr(N__6190));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_6_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_6_6_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_6_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(N__4578),
            .in2(_gnd_net_),
            .in3(N__4375),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4372),
            .ce(),
            .sr(N__6190));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_6_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_6_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_6_7_0  (
            .in0(N__4498),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9948),
            .ce(N__6407),
            .sr(N__10539));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_6_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_6_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_6_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4480),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9948),
            .ce(N__6407),
            .sr(N__10539));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_6_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_6_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_6_7_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_6_7_3  (
            .in0(N__4468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9948),
            .ce(N__6407),
            .sr(N__10539));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_6_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_6_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4450),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9948),
            .ce(N__6407),
            .sr(N__10539));
    defparam DBRn_ibuf_RNIBAB_LC_6_10_1.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_6_10_1.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_6_10_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_6_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4713),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_4 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_4  (
            .in0(N__4438),
            .in1(N__4678),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.N_402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_7_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_7_5_1 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIOO5O1_3_LC_7_5_1  (
            .in0(N__6885),
            .in1(N__7194),
            .in2(N__7344),
            .in3(N__7033),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDs_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_7_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_7_6_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_7_6_1  (
            .in0(N__4855),
            .in1(N__6352),
            .in2(_gnd_net_),
            .in3(N__6373),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m93_i_a2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_7_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_7_6_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_7_6_2  (
            .in0(N__6331),
            .in1(N__6199),
            .in2(N__4423),
            .in3(N__5944),
            .lcout(\U712_CHIP_RAM.N_428 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_7_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_7_6_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__4602),
            .in2(_gnd_net_),
            .in3(N__4590),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH5lto7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_7_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_7_6_4 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_7_6_4  (
            .in0(N__10207),
            .in1(N__4579),
            .in2(N__4567),
            .in3(N__4513),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9943),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_7_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_7_6_5 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_7_6_5  (
            .in0(N__4563),
            .in1(N__4551),
            .in2(N__4540),
            .in3(N__4524),
            .lcout(\U712_CHIP_RAM.REFRESH5lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ORT_7_LC_7_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ORT_7_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ORT_7_LC_7_6_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6ORT_7_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(N__4935),
            .in2(_gnd_net_),
            .in3(N__5008),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDs_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJNSTA_0_LC_7_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJNSTA_0_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJNSTA_0_LC_7_7_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIJNSTA_0_LC_7_7_0  (
            .in0(N__10566),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5513),
            .lcout(\U712_CHIP_RAM.N_194_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_7_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_7_7_1  (
            .in0(N__6657),
            .in1(N__4734),
            .in2(_gnd_net_),
            .in3(N__4504),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_430_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_7_2 .LUT_INIT=16'b1100000011001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_7_7_2  (
            .in0(N__5707),
            .in1(N__10199),
            .in2(N__4507),
            .in3(N__5772),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9945),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_7_3 .LUT_INIT=16'b1000100011001000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_7_3  (
            .in0(N__4639),
            .in1(N__10193),
            .in2(N__4900),
            .in3(N__11675),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9945),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_7_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_7_7_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_4_LC_7_7_4  (
            .in0(N__4735),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10200),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9945),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_7_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_7_7_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_7_7_5  (
            .in0(N__4872),
            .in1(N__4854),
            .in2(N__4899),
            .in3(N__5706),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_7_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_7_7_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_7_7_6  (
            .in0(N__6658),
            .in1(N__7645),
            .in2(N__10206),
            .in3(N__4618),
            .lcout(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9945),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_7_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_7_7_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3M1M2_1_LC_7_7_7  (
            .in0(N__7159),
            .in1(N__6856),
            .in2(_gnd_net_),
            .in3(N__7221),
            .lcout(\U712_CHIP_RAM.m101_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_7_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_7_8_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_7_8_0  (
            .in0(N__4837),
            .in1(N__10202),
            .in2(N__5727),
            .in3(N__5484),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_7_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_7_8_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_7_8_1  (
            .in0(N__4965),
            .in1(N__5032),
            .in2(N__5007),
            .in3(N__4928),
            .lcout(\U712_CHIP_RAM.N_307 ),
            .ltout(\U712_CHIP_RAM.N_307_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_7_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_7_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_3_LC_7_8_2  (
            .in0(N__6777),
            .in1(N__6859),
            .in2(N__4612),
            .in3(N__7307),
            .lcout(\U712_CHIP_RAM.N_467 ),
            .ltout(\U712_CHIP_RAM.N_467_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_7_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_7_8_3 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__7023),
            .in2(N__4609),
            .in3(N__7129),
            .lcout(\U712_CHIP_RAM.N_476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU7TF5_LC_7_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU7TF5_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU7TF5_LC_7_8_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU7TF5_LC_7_8_4  (
            .in0(N__7024),
            .in1(N__5463),
            .in2(N__7170),
            .in3(N__5421),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKHPV5_LC_7_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKHPV5_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKHPV5_LC_7_8_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKHPV5_LC_7_8_5  (
            .in0(N__10565),
            .in1(_gnd_net_),
            .in2(N__4606),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_8_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_7_8_6  (
            .in0(N__7025),
            .in1(_gnd_net_),
            .in2(N__7171),
            .in3(N__5422),
            .lcout(\U712_CHIP_RAM.N_440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_8_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_8_7  (
            .in0(N__5423),
            .in1(N__7026),
            .in2(N__7195),
            .in3(N__5714),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9949),
            .ce(N__4723),
            .sr(N__10529));
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_7_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_7_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_7_9_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_3_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(N__10201),
            .in2(_gnd_net_),
            .in3(N__9982),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9954),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_9_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(N__10564),
            .in2(_gnd_net_),
            .in3(N__5088),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_0_LC_7_10_4.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_7_10_4.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_7_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_0_LC_7_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4714),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9959),
            .ce(),
            .sr(N__10515));
    defparam \U712_REG_SM.WRITE_CYCLE_LC_7_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_7_13_2 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_REG_SM.WRITE_CYCLE_LC_7_13_2  (
            .in0(N__10380),
            .in1(N__7455),
            .in2(_gnd_net_),
            .in3(N__8522),
            .lcout(\U712_REG_SM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9968),
            .ce(),
            .sr(N__10500));
    defparam \U712_REG_SM.LDSn_RNO_0_LC_7_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_7_14_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_REG_SM.LDSn_RNO_0_LC_7_14_0  (
            .in0(N__11208),
            .in1(N__11332),
            .in2(N__11100),
            .in3(N__10384),
            .lcout(\U712_REG_SM.N_404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_7_16_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_7_16_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_7_16_3  (
            .in0(N__4674),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4651),
            .lcout(\U712_CHIP_RAM.N_419 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_LC_8_4_0  (
            .in0(N__11676),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7441),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_5_0 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_8_5_0  (
            .in0(N__6172),
            .in1(N__7187),
            .in2(N__4801),
            .in3(N__4912),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMDsr_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_5_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_5_1 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_8_5_1  (
            .in0(N__6691),
            .in1(N__5518),
            .in2(N__4804),
            .in3(N__8138),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9936),
            .ce(),
            .sr(N__10540));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_1_LC_8_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_1_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_1_LC_8_5_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_1_LC_8_5_4  (
            .in0(N__4796),
            .in1(N__5041),
            .in2(N__4981),
            .in3(N__5137),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_2_LC_8_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_2_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_2_LC_8_5_6 .LUT_INIT=16'b1111111111011110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_2_2_LC_8_5_6  (
            .in0(N__7032),
            .in1(N__4974),
            .in2(N__6793),
            .in3(N__5040),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMDsr_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_2_LC_8_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_2_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_2_LC_8_5_7 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_2_LC_8_5_7  (
            .in0(N__7335),
            .in1(N__4797),
            .in2(N__4786),
            .in3(N__6791),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_1_LC_8_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_1_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_1_LC_8_6_0 .LUT_INIT=16'b0010001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_1_LC_8_6_0  (
            .in0(N__6886),
            .in1(N__7031),
            .in2(N__4879),
            .in3(N__7186),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_396_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_1_LC_8_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_1_LC_8_6_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_1_LC_8_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_1_LC_8_6_1  (
            .in0(N__4774),
            .in1(N__4761),
            .in2(N__4783),
            .in3(N__4780),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9939),
            .ce(N__4750),
            .sr(N__10535));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_1_LC_8_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_1_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_1_LC_8_6_2 .LUT_INIT=16'b1000100011001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_1_1_LC_8_6_2  (
            .in0(N__7336),
            .in1(N__7185),
            .in2(N__5731),
            .in3(N__7030),
            .lcout(\U712_CHIP_RAM.N_397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_2_LC_8_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_2_LC_8_6_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_2_LC_8_6_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_2_LC_8_6_3  (
            .in0(N__4768),
            .in1(N__5494),
            .in2(N__5269),
            .in3(N__4762),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9939),
            .ce(N__4750),
            .sr(N__10535));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_6_6  (
            .in0(N__6784),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7833),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_8_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_8_7_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_8_7_0  (
            .in0(N__7304),
            .in1(N__4972),
            .in2(_gnd_net_),
            .in3(N__5033),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_7_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_1_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__6855),
            .in2(_gnd_net_),
            .in3(N__6752),
            .lcout(\U712_CHIP_RAM.N_305 ),
            .ltout(\U712_CHIP_RAM.N_305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_8_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_8_7_2 .LUT_INIT=16'b1010010110100001;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI7MCB2_LC_8_7_2  (
            .in0(N__7302),
            .in1(N__5702),
            .in2(N__4903),
            .in3(N__6977),
            .lcout(\U712_CHIP_RAM.N_376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_8_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_8_7_3 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_8_7_3  (
            .in0(N__4892),
            .in1(N__4871),
            .in2(_gnd_net_),
            .in3(N__4853),
            .lcout(\U712_CHIP_RAM.N_325 ),
            .ltout(\U712_CHIP_RAM.N_325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNICN5A2_2_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNICN5A2_2_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNICN5A2_2_LC_8_7_4 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNICN5A2_2_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__6978),
            .in2(N__4831),
            .in3(N__6602),
            .lcout(\U712_CHIP_RAM.N_436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_8_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_8_7_5 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIGB4P1_3_LC_8_7_5  (
            .in0(N__10198),
            .in1(N__7160),
            .in2(N__7021),
            .in3(N__7303),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m101_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7AC23_0_LC_8_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7AC23_0_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7AC23_0_LC_8_7_6 .LUT_INIT=16'b1111000111110101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI7AC23_0_LC_8_7_6  (
            .in0(N__7161),
            .in1(N__6758),
            .in2(N__4828),
            .in3(N__6982),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m101_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITD0EA_0_LC_8_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITD0EA_0_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITD0EA_0_LC_8_7_7 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITD0EA_0_LC_8_7_7  (
            .in0(N__4825),
            .in1(N__4819),
            .in2(N__4813),
            .in3(N__4810),
            .lcout(\U712_CHIP_RAM.N_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_8_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_8_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__6773),
            .in2(_gnd_net_),
            .in3(N__5771),
            .lcout(\U712_CHIP_RAM.LATCH_CLK_6 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_8_1  (
            .in0(N__5393),
            .in1(N__6873),
            .in2(_gnd_net_),
            .in3(N__5050),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__9946),
            .ce(N__5331),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__7018),
            .in2(_gnd_net_),
            .in3(N__5047),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3  (
            .in0(N__5394),
            .in1(N__7325),
            .in2(_gnd_net_),
            .in3(N__5044),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__9946),
            .ce(N__5331),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4  (
            .in0(N__5382),
            .in1(N__5039),
            .in2(_gnd_net_),
            .in3(N__5011),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__9946),
            .ce(N__5331),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5  (
            .in0(N__5395),
            .in1(N__5006),
            .in2(_gnd_net_),
            .in3(N__4984),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__9946),
            .ce(N__5331),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6  (
            .in0(N__5383),
            .in1(N__4973),
            .in2(_gnd_net_),
            .in3(N__4942),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__9946),
            .ce(N__5331),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7  (
            .in0(N__4936),
            .in1(N__5384),
            .in2(_gnd_net_),
            .in3(N__4939),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9946),
            .ce(N__5331),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_9_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_9_0  (
            .in0(N__7126),
            .in1(N__7306),
            .in2(N__6792),
            .in3(N__6986),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_0_a3_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_9_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_9_1  (
            .in0(N__6764),
            .in1(N__5652),
            .in2(N__7022),
            .in3(N__7127),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_2_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_9_2 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_8_9_2  (
            .in0(N__7128),
            .in1(_gnd_net_),
            .in2(N__5140),
            .in3(N__10172),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9950),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_1_LC_8_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_1_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_1_LC_8_9_3 .LUT_INIT=16'b1111000011010011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_3_1_LC_8_9_3  (
            .in0(N__6985),
            .in1(N__6858),
            .in2(N__6778),
            .in3(N__7125),
            .lcout(\U712_CHIP_RAM.N_378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_8_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_8_9_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_8_9_4  (
            .in0(N__7124),
            .in1(N__6984),
            .in2(N__5732),
            .in3(N__5420),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_8_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_8_9_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI41RO8_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5128),
            .in3(N__5838),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_8_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_8_9_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_3_LC_8_9_6  (
            .in0(N__6857),
            .in1(N__7305),
            .in2(_gnd_net_),
            .in3(N__7222),
            .lcout(\U712_CHIP_RAM.N_551 ),
            .ltout(\U712_CHIP_RAM.N_551_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_8_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_8_9_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOBA64_LC_8_9_7  (
            .in0(N__6983),
            .in1(N__7123),
            .in2(N__5125),
            .in3(N__6167),
            .lcout(\U712_CHIP_RAM.N_435 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_8_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_8_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_8_10_0 .LUT_INIT=16'b1111011100000010;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_8_10_0  (
            .in0(N__5122),
            .in1(N__7357),
            .in2(N__7246),
            .in3(N__5100),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9955),
            .ce(),
            .sr(N__10509));
    defparam \U712_CHIP_RAM.DBENn_LC_8_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_8_10_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_8_10_1 .LUT_INIT=16'b0101111111001100;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_8_10_1  (
            .in0(N__5434),
            .in1(N__5800),
            .in2(N__5746),
            .in3(N__5089),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9955),
            .ce(),
            .sr(N__10509));
    defparam \U712_CHIP_RAM.DBDIR_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_8_10_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_8_10_7 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_8_10_7  (
            .in0(N__5589),
            .in1(N__5061),
            .in2(_gnd_net_),
            .in3(N__5562),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9955),
            .ce(),
            .sr(N__10509));
    defparam \U712_REG_SM.REGENn_LC_8_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_8_11_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_8_11_6 .LUT_INIT=16'b1011010010110000;
    LogicCell40 \U712_REG_SM.REGENn_LC_8_11_6  (
            .in0(N__7958),
            .in1(N__5167),
            .in2(N__5214),
            .in3(N__5239),
            .lcout(REGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9960),
            .ce(),
            .sr(N__10504));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_12_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_8_12_0 .LUT_INIT=16'b1100110011001101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_8_12_0  (
            .in0(N__5755),
            .in1(N__5254),
            .in2(N__7680),
            .in3(N__8035),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9963),
            .ce(),
            .sr(N__10501));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_8_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_8_13_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_8_13_2  (
            .in0(N__7570),
            .in1(N__8038),
            .in2(N__7681),
            .in3(N__5183),
            .lcout(\U712_REG_SM.N_412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_13_5 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_8_13_5  (
            .in0(N__10166),
            .in1(N__5248),
            .in2(N__5188),
            .in3(N__8467),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9965),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_8_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_8_13_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_8_13_7  (
            .in0(N__5182),
            .in1(N__5238),
            .in2(N__7535),
            .in3(N__7940),
            .lcout(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_RNO_0_LC_8_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_RNO_0_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REGENn_RNO_0_LC_8_14_1 .LUT_INIT=16'b0000100001011000;
    LogicCell40 \U712_REG_SM.REGENn_RNO_0_LC_8_14_1  (
            .in0(N__5213),
            .in1(N__8495),
            .in2(N__7537),
            .in3(N__5187),
            .lcout(\U712_REG_SM.REGENn_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDSn_RNO_0_LC_8_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_8_15_7 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \U712_REG_SM.UDSn_RNO_0_LC_8_15_7  (
            .in0(N__11342),
            .in1(N__11087),
            .in2(N__11263),
            .in3(N__10385),
            .lcout(\U712_REG_SM.N_459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBR_COUNT_1_LC_9_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_COUNT_1_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_1_LC_9_5_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_1_LC_9_5_1  (
            .in0(N__5939),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6231),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9934),
            .ce(),
            .sr(N__6676));
    defparam \U712_CHIP_RAM.DBR_COUNT_0_LC_9_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_COUNT_0_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_0_LC_9_5_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_0_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5938),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9934),
            .ce(),
            .sr(N__6676));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_1  (
            .in0(N__5158),
            .in1(N__5275),
            .in2(_gnd_net_),
            .in3(N__8857),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_9_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_9_6_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_9_6_2  (
            .in0(N__8858),
            .in1(N__5314),
            .in2(_gnd_net_),
            .in3(N__5533),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_9_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_9_6_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_9_6_3  (
            .in0(N__11610),
            .in1(N__8859),
            .in2(N__5296),
            .in3(N__8203),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_9_6_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_9_6_4  (
            .in0(N__5293),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9937),
            .ce(N__6409),
            .sr(N__10530));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_6_6 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_9_6_6  (
            .in0(N__8131),
            .in1(N__8888),
            .in2(_gnd_net_),
            .in3(N__8159),
            .lcout(\U712_CHIP_RAM.CMA_5_i_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIUI4B1_0_LC_9_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIUI4B1_0_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIUI4B1_0_LC_9_6_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIUI4B1_0_LC_9_6_7  (
            .in0(N__8158),
            .in1(N__8130),
            .in2(N__9572),
            .in3(N__8856),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_9_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_9_7_0 .LUT_INIT=16'b1100110100001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_3_3_LC_9_7_0  (
            .in0(N__6760),
            .in1(N__7308),
            .in2(N__7188),
            .in3(N__7002),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMT791_1_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMT791_1_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMT791_1_LC_9_7_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIMT791_1_LC_9_7_1  (
            .in0(N__7162),
            .in1(N__6863),
            .in2(_gnd_net_),
            .in3(N__6759),
            .lcout(\U712_CHIP_RAM.N_555 ),
            .ltout(\U712_CHIP_RAM.N_555_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_7_2 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_3_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__6603),
            .in2(N__5257),
            .in3(N__7309),
            .lcout(\U712_CHIP_RAM.N_390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_7_3 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_9_7_3  (
            .in0(N__7004),
            .in1(N__7167),
            .in2(_gnd_net_),
            .in3(N__6865),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMDsr_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_7_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_7_4 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_7_4  (
            .in0(N__6538),
            .in1(N__5514),
            .in2(N__5497),
            .in3(N__9566),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9940),
            .ce(),
            .sr(N__10522));
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_2_LC_9_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_2_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_2_LC_9_7_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_ess_RNO_0_2_LC_9_7_7  (
            .in0(N__7003),
            .in1(N__7166),
            .in2(_gnd_net_),
            .in3(N__6864),
            .lcout(\U712_CHIP_RAM.N_449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIB0JV5_LC_9_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIB0JV5_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIB0JV5_LC_9_8_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIB0JV5_LC_9_8_1  (
            .in0(N__5488),
            .in1(N__5470),
            .in2(_gnd_net_),
            .in3(N__5733),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_8_2  (
            .in0(N__10173),
            .in1(N__5452),
            .in2(N__5446),
            .in3(N__5385),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9944),
            .ce(N__5335),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_9_8_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__7384),
            .in2(_gnd_net_),
            .in3(N__6753),
            .lcout(\U712_CHIP_RAM.N_304 ),
            .ltout(\U712_CHIP_RAM.N_304_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_9_8_4 .LUT_INIT=16'b0011000010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNID3LR1_0_LC_9_8_4  (
            .in0(N__6754),
            .in1(N__6999),
            .in2(N__5443),
            .in3(N__7168),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_312_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIBB455_0_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIBB455_0_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIBB455_0_LC_9_8_5 .LUT_INIT=16'b1111001100110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIBB455_0_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__10174),
            .in2(N__5440),
            .in3(N__5651),
            .lcout(\U712_CHIP_RAM.N_326 ),
            .ltout(\U712_CHIP_RAM.N_326_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_9_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_9_8_6 .LUT_INIT=16'b1111101111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIA8V79_LC_9_8_6  (
            .in0(N__7169),
            .in1(N__7000),
            .in2(N__5437),
            .in3(N__5430),
            .lcout(\U712_CHIP_RAM.N_39 ),
            .ltout(\U712_CHIP_RAM.N_39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_7 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_9_8_7  (
            .in0(N__5362),
            .in1(N__5353),
            .in2(N__5344),
            .in3(N__5341),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9944),
            .ce(N__5335),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__7019),
            .in2(_gnd_net_),
            .in3(N__9754),
            .lcout(\U712_CHIP_RAM.DBENn_7_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_9_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_9_1  (
            .in0(N__5737),
            .in1(N__10389),
            .in2(_gnd_net_),
            .in3(N__5596),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_344_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_9_9_2 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_9_9_2  (
            .in0(N__10171),
            .in1(N__5662),
            .in2(N__5656),
            .in3(N__7386),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9947),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_9_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_9_9_3  (
            .in0(N__7020),
            .in1(N__7366),
            .in2(N__7190),
            .in3(N__5653),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER41_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_9_9_4 .LUT_INIT=16'b1010100000001000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_9_9_4  (
            .in0(N__10170),
            .in1(N__5607),
            .in2(N__5635),
            .in3(N__5632),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9947),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_9_9_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIDTSL_LC_9_9_5  (
            .in0(N__7385),
            .in1(N__6866),
            .in2(_gnd_net_),
            .in3(N__11568),
            .lcout(\U712_CHIP_RAM.N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_9_9_6 .LUT_INIT=16'b0101000011000000;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_9_9_6  (
            .in0(N__5595),
            .in1(N__11738),
            .in2(N__10197),
            .in3(N__5563),
            .lcout(DMA_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9947),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_9_10_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_9_10_0  (
            .in0(N__5854),
            .in1(N__5551),
            .in2(N__10867),
            .in3(N__5532),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9951),
            .ce(),
            .sr(N__10505));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_1  (
            .in0(N__11606),
            .in1(N__5853),
            .in2(_gnd_net_),
            .in3(N__5839),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9951),
            .ce(),
            .sr(N__10505));
    defparam DBR_SYNC_1_LC_9_10_3.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_9_10_3.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_9_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_9_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5827),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9951),
            .ce(),
            .sr(N__10505));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_9_11_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_0_LC_9_11_0  (
            .in0(N__5801),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5781),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_11_3 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_11_3  (
            .in0(N__8030),
            .in1(N__7600),
            .in2(N__7543),
            .in3(N__7632),
            .lcout(),
            .ltout(\U712_REG_SM.N_413_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_9_11_4 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_9_11_4  (
            .in0(N__10183),
            .in1(N__7542),
            .in2(N__5818),
            .in3(N__7959),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9956),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFFA4_LC_9_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFFA4_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFFA4_LC_9_11_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFFA4_LC_9_11_6  (
            .in0(N__5802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5782),
            .lcout(\U712_CHIP_RAM.m50_i_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_9_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_9_12_0 .LUT_INIT=16'b1000100011101110;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_9_12_0  (
            .in0(N__7568),
            .in1(N__7536),
            .in2(_gnd_net_),
            .in3(N__7957),
            .lcout(\U712_REG_SM.N_308 ),
            .ltout(\U712_REG_SM.N_308_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_9_12_1 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_9_12_1  (
            .in0(N__10163),
            .in1(N__8034),
            .in2(N__5749),
            .in3(N__7569),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9961),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_12_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_12_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_9_12_3  (
            .in0(N__10160),
            .in1(N__9210),
            .in2(_gnd_net_),
            .in3(N__8611),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9961),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_9_12_4  (
            .in0(N__5908),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10161),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9961),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_9_12_5  (
            .in0(N__10162),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6141),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9961),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_9_12_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_9_12_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__6140),
            .in2(_gnd_net_),
            .in3(N__5907),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_9_13_0 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_9_13_0  (
            .in0(N__10165),
            .in1(N__5896),
            .in2(N__8524),
            .in3(N__8494),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9964),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_9_13_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__7594),
            .in2(_gnd_net_),
            .in3(N__8492),
            .lcout(\U712_REG_SM.N_328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_13_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_13_3  (
            .in0(N__7595),
            .in1(N__7641),
            .in2(N__7534),
            .in3(N__7936),
            .lcout(),
            .ltout(\U712_REG_SM.N_410_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_9_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_13_4 .LUT_INIT=16'b1110110011100100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_9_13_4  (
            .in0(N__10164),
            .in1(N__7422),
            .in2(N__5899),
            .in3(N__7462),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9964),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_9_13_6 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_9_13_6  (
            .in0(N__7566),
            .in1(N__7506),
            .in2(N__7956),
            .in3(N__8493),
            .lcout(\U712_REG_SM.un1_REGENn_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_13_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7533),
            .in3(N__7935),
            .lcout(\U712_REG_SM.N_331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_14_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_14_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_9_14_0  (
            .in0(N__5890),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9966),
            .ce(),
            .sr(N__10493));
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_14_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6151),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9966),
            .ce(),
            .sr(N__10493));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_9_14_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_9_14_3 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_9_14_3 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_9_14_3  (
            .in0(N__6082),
            .in1(N__6145),
            .in2(N__9211),
            .in3(N__8610),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9966),
            .ce(),
            .sr(N__10493));
    defparam \U712_REG_SM.LDSn_LC_9_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_9_14_4 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_9_14_4 .LUT_INIT=16'b1011101110111000;
    LogicCell40 \U712_REG_SM.LDSn_LC_9_14_4  (
            .in0(N__6042),
            .in1(N__7989),
            .in2(N__7960),
            .in3(N__6067),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9966),
            .ce(),
            .sr(N__10493));
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_14_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6018),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9966),
            .ce(),
            .sr(N__10493));
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_14_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_9_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5989),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9966),
            .ce(),
            .sr(N__10493));
    defparam \U712_REG_SM.UDSn_LC_9_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_9_15_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_9_15_0 .LUT_INIT=16'b1111001111100010;
    LogicCell40 \U712_REG_SM.UDSn_LC_9_15_0  (
            .in0(N__5983),
            .in1(N__7990),
            .in2(N__5961),
            .in3(N__7951),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9969),
            .ce(),
            .sr(N__10488));
    defparam \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_10_5_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_10_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U712_CHIP_RAM.un3_DBR_COUNT_cry_1_c_LC_10_5_0  (
            .in0(_gnd_net_),
            .in1(N__6230),
            .in2(N__5940),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_5_0_),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBR_COUNT_2_LC_10_5_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_2_LC_10_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_2_LC_10_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_2_LC_10_5_1  (
            .in0(_gnd_net_),
            .in1(N__6244),
            .in2(_gnd_net_),
            .in3(N__5914),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_1 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_2 ),
            .clk(N__9929),
            .ce(),
            .sr(N__6675));
    defparam \U712_CHIP_RAM.DBR_COUNT_3_LC_10_5_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_3_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_3_LC_10_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_3_LC_10_5_2  (
            .in0(_gnd_net_),
            .in1(N__6256),
            .in2(_gnd_net_),
            .in3(N__5911),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_2 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_3 ),
            .clk(N__9929),
            .ce(),
            .sr(N__6675));
    defparam \U712_CHIP_RAM.DBR_COUNT_4_LC_10_5_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_4_LC_10_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_4_LC_10_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_4_LC_10_5_3  (
            .in0(_gnd_net_),
            .in1(N__6369),
            .in2(_gnd_net_),
            .in3(N__6355),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_3 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_4 ),
            .clk(N__9929),
            .ce(),
            .sr(N__6675));
    defparam \U712_CHIP_RAM.DBR_COUNT_5_LC_10_5_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_5_LC_10_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_5_LC_10_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_5_LC_10_5_4  (
            .in0(_gnd_net_),
            .in1(N__6348),
            .in2(_gnd_net_),
            .in3(N__6334),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_4 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_5 ),
            .clk(N__9929),
            .ce(),
            .sr(N__6675));
    defparam \U712_CHIP_RAM.DBR_COUNT_6_LC_10_5_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.DBR_COUNT_6_LC_10_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_6_LC_10_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_6_LC_10_5_5  (
            .in0(_gnd_net_),
            .in1(N__6327),
            .in2(_gnd_net_),
            .in3(N__6313),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un3_DBR_COUNT_cry_5 ),
            .carryout(\U712_CHIP_RAM.un3_DBR_COUNT_cry_6 ),
            .clk(N__9929),
            .ce(),
            .sr(N__6675));
    defparam \U712_CHIP_RAM.DBR_COUNT_7_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_COUNT_7_LC_10_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DBR_COUNT_7_LC_10_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.DBR_COUNT_7_LC_10_5_6  (
            .in0(_gnd_net_),
            .in1(N__6211),
            .in2(_gnd_net_),
            .in3(N__6310),
            .lcout(\U712_CHIP_RAM.DBR_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9929),
            .ce(),
            .sr(N__6675));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_10_6_0  (
            .in0(N__6307),
            .in1(N__6433),
            .in2(_gnd_net_),
            .in3(N__8890),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_6_2  (
            .in0(N__6276),
            .in1(N__6463),
            .in2(_gnd_net_),
            .in3(N__8891),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_10_6_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_2_LC_10_6_6  (
            .in0(N__6255),
            .in1(N__6243),
            .in2(N__6232),
            .in3(N__6210),
            .lcout(\U712_CHIP_RAM.m93_i_a2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIB72G2_3_LC_10_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIB72G2_3_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIB72G2_3_LC_10_6_7 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIB72G2_3_LC_10_6_7  (
            .in0(N__8889),
            .in1(N__9565),
            .in2(N__8177),
            .in3(N__6186),
            .lcout(\U712_CHIP_RAM.un1_CMA25_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_7_0 .LUT_INIT=16'b1110011110100111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_10_7_0  (
            .in0(N__7017),
            .in1(N__6891),
            .in2(N__7345),
            .in3(N__6168),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m123_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_7_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_7_1  (
            .in0(N__7189),
            .in1(N__6607),
            .in2(N__6586),
            .in3(N__7244),
            .lcout(\U712_CHIP_RAM.N_190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_3  (
            .in0(N__6583),
            .in1(N__6562),
            .in2(_gnd_net_),
            .in3(N__8960),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_4  (
            .in0(N__8961),
            .in1(N__11611),
            .in2(N__6553),
            .in3(N__9292),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_7_6 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_7_6  (
            .in0(N__7243),
            .in1(N__6550),
            .in2(_gnd_net_),
            .in3(N__6544),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_7  (
            .in0(N__6522),
            .in1(N__6487),
            .in2(_gnd_net_),
            .in3(N__8959),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_10_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6478),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9941),
            .ce(N__6408),
            .sr(N__10510));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_10_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_10_8_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_10_8_2  (
            .in0(N__6454),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9941),
            .ce(N__6408),
            .sr(N__10510));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_10_8_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_10_8_5  (
            .in0(N__6424),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9941),
            .ce(N__6408),
            .sr(N__10510));
    defparam \U712_BUFFERS.N_167_i_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_167_i_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_167_i_LC_10_9_0 .LUT_INIT=16'b0000000011101010;
    LogicCell40 \U712_BUFFERS.N_167_i_LC_10_9_0  (
            .in0(N__11573),
            .in1(N__11845),
            .in2(N__10318),
            .in3(N__7434),
            .lcout(N_167_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_10_9_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_0_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__7387),
            .in2(_gnd_net_),
            .in3(N__6772),
            .lcout(\U712_CHIP_RAM.N_321 ),
            .ltout(\U712_CHIP_RAM.N_321_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_9_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_10_9_4  (
            .in0(N__11572),
            .in1(N__7016),
            .in2(N__7360),
            .in3(N__6890),
            .lcout(),
            .ltout(\U712_CHIP_RAM.m77_0_a2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_9_5 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_9_5  (
            .in0(N__7356),
            .in1(N__7340),
            .in2(N__7249),
            .in3(N__7245),
            .lcout(\U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_9_7 .LUT_INIT=16'b0111111101101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_9_7  (
            .in0(N__7172),
            .in1(N__7001),
            .in2(N__6892),
            .in3(N__6771),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDsr_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_10_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_10_10_2 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNIEU0T_1_LC_10_10_2  (
            .in0(N__10152),
            .in1(N__6645),
            .in2(_gnd_net_),
            .in3(N__7636),
            .lcout(\U712_CHIP_RAM.CAS_SYNC_RNIEU0TZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_10_11_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_10_11_0  (
            .in0(N__10056),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6613),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9952),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNIVU9S_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNIVU9S_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNIVU9S_LC_10_11_5 .LUT_INIT=16'b0111011100000111;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNIVU9S_LC_10_11_5  (
            .in0(N__11580),
            .in1(N__7969),
            .in2(N__9255),
            .in3(N__10314),
            .lcout(N_202_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_10_11_7 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_10_11_7  (
            .in0(N__11835),
            .in1(N__10055),
            .in2(_gnd_net_),
            .in3(N__10313),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9952),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_12_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_12_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_12_0 .LUT_INIT=16'b0000111000001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_10_12_0  (
            .in0(N__7765),
            .in1(N__7759),
            .in2(N__8609),
            .in3(N__8530),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9957),
            .ce(),
            .sr(N__10495));
    defparam \U712_CYCLE_TERM.TACK_EN_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_10_12_3 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_LC_10_12_3  (
            .in0(N__7758),
            .in1(N__7696),
            .in2(_gnd_net_),
            .in3(N__8185),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9957),
            .ce(),
            .sr(N__10495));
    defparam \U712_REG_SM.REG_TACK_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_10_12_5 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_10_12_5  (
            .in0(N__8575),
            .in1(N__7673),
            .in2(N__7654),
            .in3(N__7996),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9957),
            .ce(),
            .sr(N__10495));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_10_13_0 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_10_13_0  (
            .in0(N__7942),
            .in1(N__8037),
            .in2(_gnd_net_),
            .in3(N__7526),
            .lcout(\U712_REG_SM.N_406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_13_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__7527),
            .in2(_gnd_net_),
            .in3(N__7640),
            .lcout(),
            .ltout(\U712_REG_SM.N_330_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_10_13_3 .LUT_INIT=16'b0010000000100010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_10_13_3  (
            .in0(N__10159),
            .in1(N__7576),
            .in2(N__7603),
            .in3(N__7944),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9962),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_10_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_10_13_4 .LUT_INIT=16'b0000000011111011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_10_13_4  (
            .in0(N__7943),
            .in1(N__8496),
            .in2(N__7538),
            .in3(N__7596),
            .lcout(\U712_REG_SM.STATE_COUNTc_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_13_5 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_13_5  (
            .in0(N__7567),
            .in1(N__7522),
            .in2(_gnd_net_),
            .in3(N__7941),
            .lcout(\U712_REG_SM.N_373 ),
            .ltout(\U712_REG_SM.N_373_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_6 .LUT_INIT=16'b0100111001001110;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_10_13_6  (
            .in0(N__7456),
            .in1(N__8036),
            .in2(N__7999),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.N_130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_RNO_LC_10_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_10_14_1 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U712_REG_SM.ASn_ess_RNO_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__10562),
            .in2(_gnd_net_),
            .in3(N__7985),
            .lcout(\U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m37_i_o2_LC_10_14_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m37_i_o2_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m37_i_o2_LC_10_14_5 .LUT_INIT=16'b1111101010001111;
    LogicCell40 \U712_CHIP_RAM.m37_i_o2_LC_10_14_5  (
            .in0(N__11447),
            .in1(N__11349),
            .in2(N__11149),
            .in3(N__11207),
            .lcout(\U712_CHIP_RAM.N_335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_LC_10_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_LC_10_15_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_ess_LC_10_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.ASn_ess_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7955),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9967),
            .ce(N__7864),
            .sr(N__10487));
    defparam \U712_BUFFERS.N_165_i_LC_10_19_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_165_i_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_165_i_LC_10_19_1 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \U712_BUFFERS.N_165_i_LC_10_19_1  (
            .in0(N__11831),
            .in1(N__10299),
            .in2(_gnd_net_),
            .in3(N__11757),
            .lcout(N_165_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_11_3_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_3_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_3_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_3_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RASn_LC_11_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_11_4_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_11_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8179),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9925),
            .ce(),
            .sr(N__10531));
    defparam \U712_CHIP_RAM.WEn_LC_11_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_11_4_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_11_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_11_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8143),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9925),
            .ce(),
            .sr(N__10531));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_5_0 .LUT_INIT=16'b0100000000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_5_0  (
            .in0(N__11655),
            .in1(N__9271),
            .in2(N__8966),
            .in3(N__8737),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIE8IL_0_LC_11_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIE8IL_0_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIE8IL_0_LC_11_5_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIE8IL_0_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__8178),
            .in2(_gnd_net_),
            .in3(N__8139),
            .lcout(\U712_CHIP_RAM.N_314 ),
            .ltout(\U712_CHIP_RAM.N_314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_5_4 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_5_4  (
            .in0(N__11654),
            .in1(N__9270),
            .in2(N__8110),
            .in3(N__8949),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_5_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_11_5_7  (
            .in0(N__8107),
            .in1(N__11656),
            .in2(_gnd_net_),
            .in3(N__9604),
            .lcout(\U712_CHIP_RAM.N_361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_6_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_6_0  (
            .in0(N__8942),
            .in1(N__11658),
            .in2(N__8086),
            .in3(N__9394),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI1HUV2_3_LC_11_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI1HUV2_3_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI1HUV2_3_LC_11_6_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI1HUV2_3_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__10563),
            .in2(_gnd_net_),
            .in3(N__8077),
            .lcout(\U712_CHIP_RAM.un1_CMA25_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_6_2 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_6_2  (
            .in0(N__11659),
            .in1(N__8071),
            .in2(N__8965),
            .in3(N__9370),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNII0RI_LC_11_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNII0RI_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNII0RI_LC_11_6_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNII0RI_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(N__11657),
            .in2(_gnd_net_),
            .in3(N__8938),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_RNII0RIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_6_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_6_6  (
            .in0(N__11660),
            .in1(N__8065),
            .in2(_gnd_net_),
            .in3(N__9382),
            .lcout(\U712_CHIP_RAM.N_367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_6_7 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_6_7  (
            .in0(N__8053),
            .in1(N__11661),
            .in2(N__8964),
            .in3(N__8230),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_11_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_11_7_0 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_11_7_0  (
            .in0(N__8817),
            .in1(N__10921),
            .in2(N__8783),
            .in3(N__8044),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9935),
            .ce(N__9451),
            .sr(N__10511));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_7_1 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_11_7_1  (
            .in0(N__9358),
            .in1(N__8818),
            .in2(N__8785),
            .in3(N__8236),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9935),
            .ce(N__9451),
            .sr(N__10511));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_11_7_2 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_11_7_2  (
            .in0(N__8819),
            .in1(N__10645),
            .in2(N__8784),
            .in3(N__8308),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9935),
            .ce(N__9451),
            .sr(N__10511));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_11_8_1 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_11_8_1  (
            .in0(N__8551),
            .in1(N__10153),
            .in2(N__8278),
            .in3(N__8269),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9938),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_8_6  (
            .in0(N__8263),
            .in1(N__8245),
            .in2(_gnd_net_),
            .in3(N__8962),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_8_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_8_7  (
            .in0(N__8963),
            .in1(N__11646),
            .in2(N__8239),
            .in3(N__9658),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_9_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_9_5  (
            .in0(N__8673),
            .in1(N__10862),
            .in2(_gnd_net_),
            .in3(N__9332),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__10598),
            .sr(N__10502));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_10_0 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_11_10_0  (
            .in0(N__10861),
            .in1(N__8672),
            .in2(N__8221),
            .in3(N__8199),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .ce(),
            .sr(N__10497));
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_12_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_12_0 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_11_12_0  (
            .in0(N__8572),
            .in1(N__8553),
            .in2(_gnd_net_),
            .in3(N__8624),
            .lcout(\U712_CYCLE_TERM.N_332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_12_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_12_2 .LUT_INIT=16'b0000000000110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_11_12_2  (
            .in0(N__8574),
            .in1(N__8625),
            .in2(N__8557),
            .in3(N__8605),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_455_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_12_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_11_12_3 .LUT_INIT=16'b0000110000001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_11_12_3  (
            .in0(N__8626),
            .in1(N__10141),
            .in2(N__8614),
            .in3(N__9208),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9953),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_12_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_12_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_11_12_6  (
            .in0(N__8573),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8552),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.START_RST_LC_11_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_11_13_3 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \U712_REG_SM.START_RST_LC_11_13_3  (
            .in0(N__8463),
            .in1(N__8523),
            .in2(_gnd_net_),
            .in3(N__8500),
            .lcout(\U712_REG_SM.START_RSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9958),
            .ce(),
            .sr(N__10489));
    defparam \U712_CHIP_RAM.CASn_LC_12_3_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_12_3_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_12_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8958),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9923),
            .ce(),
            .sr(N__10528));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_12_5_3 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_12_5_3  (
            .in0(N__8752),
            .in1(N__8437),
            .in2(N__8971),
            .in3(N__8431),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9924),
            .ce(N__9460),
            .sr(N__10514));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_12_5_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_12_5_6  (
            .in0(N__8751),
            .in1(N__9579),
            .in2(_gnd_net_),
            .in3(N__8970),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9924),
            .ce(N__9460),
            .sr(N__10514));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_5_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_5_7  (
            .in0(N__8383),
            .in1(N__8377),
            .in2(_gnd_net_),
            .in3(N__8371),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9924),
            .ce(N__9460),
            .sr(N__10514));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_12_6_0 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_12_6_0  (
            .in0(N__8820),
            .in1(N__8689),
            .in2(N__8771),
            .in3(N__9103),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9926),
            .ce(N__9459),
            .sr(N__10508));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_12_6_1 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_12_6_1  (
            .in0(N__8815),
            .in1(N__9280),
            .in2(N__8781),
            .in3(N__8986),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9926),
            .ce(N__9459),
            .sr(N__10508));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_6_3 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_12_6_3  (
            .in0(N__8816),
            .in1(N__9352),
            .in2(N__8782),
            .in3(N__9052),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9926),
            .ce(N__9459),
            .sr(N__10508));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_7_0  (
            .in0(N__9021),
            .in1(N__8998),
            .in2(_gnd_net_),
            .in3(N__8950),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_7_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_7_1  (
            .in0(N__8951),
            .in1(N__11647),
            .in2(N__8989),
            .in3(N__9343),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_4 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_4  (
            .in0(N__11648),
            .in1(N__8980),
            .in2(N__9403),
            .in3(N__8952),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_7_5 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_12_7_5  (
            .in0(N__8821),
            .in1(N__9667),
            .in2(N__8788),
            .in3(N__8770),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9928),
            .ce(N__9458),
            .sr(N__10503));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_8_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_12_8_0  (
            .in0(N__9334),
            .in1(_gnd_net_),
            .in2(N__10863),
            .in3(N__8679),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10633),
            .ce(N__10602),
            .sr(N__10499));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_8_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_12_8_2  (
            .in0(N__10857),
            .in1(N__10230),
            .in2(_gnd_net_),
            .in3(N__8680),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10633),
            .ce(N__10602),
            .sr(N__10499));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_8_3  (
            .in0(N__11010),
            .in1(N__10852),
            .in2(_gnd_net_),
            .in3(N__9649),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10633),
            .ce(N__10602),
            .sr(N__10499));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_12_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_12_8_7  (
            .in0(N__10690),
            .in1(N__9333),
            .in2(_gnd_net_),
            .in3(N__10853),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10633),
            .ce(N__10602),
            .sr(N__10499));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_12_9_3  (
            .in0(N__10848),
            .in1(N__9714),
            .in2(_gnd_net_),
            .in3(N__9821),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10600),
            .sr(N__10496));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_9_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_12_9_6  (
            .in0(N__10851),
            .in1(N__9331),
            .in2(_gnd_net_),
            .in3(N__10689),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10600),
            .sr(N__10496));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_10_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_12_10_2  (
            .in0(N__10846),
            .in1(N__9828),
            .in2(_gnd_net_),
            .in3(N__9775),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10630),
            .ce(N__10599),
            .sr(N__10494));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_10_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_12_10_3  (
            .in0(N__9829),
            .in1(N__10847),
            .in2(_gnd_net_),
            .in3(N__9707),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10630),
            .ce(N__10599),
            .sr(N__10494));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8LI41_LC_12_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8LI41_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNI8LI41_LC_12_11_1 .LUT_INIT=16'b0101000111110011;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNI8LI41_LC_12_11_1  (
            .in0(N__9220),
            .in1(N__9256),
            .in2(N__11841),
            .in3(N__11649),
            .lcout(N_200_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.m34_i_o2_LC_12_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m34_i_o2_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m34_i_o2_LC_12_13_2 .LUT_INIT=16'b1100111000111011;
    LogicCell40 \U712_CHIP_RAM.m34_i_o2_LC_12_13_2  (
            .in0(N__11430),
            .in1(N__11265),
            .in2(N__11362),
            .in3(N__11096),
            .lcout(\U712_CHIP_RAM.N_337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pll_RNI8MQ3_LC_12_14_6.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_12_14_6.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_12_14_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 pll_RNI8MQ3_LC_12_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9209),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_2.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_2.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_18_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_18_2 (
            .in0(N__10088),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CRCSn_LC_13_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_5_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_13_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_13_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9583),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9927),
            .ce(),
            .sr(N__10523));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_6_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_13_6_3  (
            .in0(N__9520),
            .in1(N__9511),
            .in2(N__11677),
            .in3(N__9490),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9930),
            .ce(N__9444),
            .sr(N__10516));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_7_0  (
            .in0(N__10838),
            .in1(N__11011),
            .in2(_gnd_net_),
            .in3(N__10957),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__10605),
            .sr(N__10512));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_7_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_7_3  (
            .in0(N__10956),
            .in1(N__10837),
            .in2(_gnd_net_),
            .in3(N__9715),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__10605),
            .sr(N__10512));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_3  (
            .in0(N__10904),
            .in1(N__10850),
            .in2(_gnd_net_),
            .in3(N__10688),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__10603),
            .sr(N__10506));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_7  (
            .in0(N__9645),
            .in1(N__10849),
            .in2(_gnd_net_),
            .in3(N__11006),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__10603),
            .sr(N__10506));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_13_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_13_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_13_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__10102),
            .in2(_gnd_net_),
            .in3(N__10213),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9942),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_13_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_13_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_13_9_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_13_9_3  (
            .in0(N__10101),
            .in1(N__10249),
            .in2(_gnd_net_),
            .in3(N__10237),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9942),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_13_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_13_9_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_2_LC_13_9_5  (
            .in0(N__10103),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9988),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9942),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_0  (
            .in0(N__9822),
            .in1(N__9774),
            .in2(_gnd_net_),
            .in3(N__10795),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10601),
            .sr(N__10498));
    defparam \U712_CHIP_RAM.m40_i_o2_LC_13_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m40_i_o2_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m40_i_o2_LC_13_13_1 .LUT_INIT=16'b1111010001011111;
    LogicCell40 \U712_CHIP_RAM.m40_i_o2_LC_13_13_1  (
            .in0(N__11449),
            .in1(N__11363),
            .in2(N__11269),
            .in3(N__11147),
            .lcout(),
            .ltout(N_334_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_177_i_LC_13_13_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_177_i_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_177_i_LC_13_13_2 .LUT_INIT=16'b0101111100010011;
    LogicCell40 \U712_BYTE_ENABLE.N_177_i_LC_13_13_2  (
            .in0(N__11653),
            .in1(N__11703),
            .in2(N__9739),
            .in3(N__10298),
            .lcout(N_177_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_0  (
            .in0(N__10950),
            .in1(N__10774),
            .in2(_gnd_net_),
            .in3(N__9697),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10632),
            .ce(N__10607),
            .sr(N__10517));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_8_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_14_8_2  (
            .in0(N__10912),
            .in1(N__10772),
            .in2(_gnd_net_),
            .in3(N__9638),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net ),
            .ce(N__10606),
            .sr(N__10513));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_9_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_9_7  (
            .in0(N__10895),
            .in1(N__10771),
            .in2(_gnd_net_),
            .in3(N__9637),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10628),
            .ce(N__10604),
            .sr(N__10507));
    defparam \U712_CHIP_RAM.m58_i_o2_LC_14_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.m58_i_o2_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.m58_i_o2_LC_14_13_6 .LUT_INIT=16'b1111000100011111;
    LogicCell40 \U712_CHIP_RAM.m58_i_o2_LC_14_13_6  (
            .in0(N__11448),
            .in1(N__11364),
            .in2(N__11262),
            .in3(N__11148),
            .lcout(),
            .ltout(N_336_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_175_i_LC_14_13_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_175_i_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_175_i_LC_14_13_7 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \U712_BYTE_ENABLE.N_175_i_LC_14_13_7  (
            .in0(N__11836),
            .in1(N__11707),
            .in2(N__11680),
            .in3(N__11671),
            .lcout(N_175_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.N_337_i_LC_14_20_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.N_337_i_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.N_337_i_LC_14_20_2 .LUT_INIT=16'b0000101110110000;
    LogicCell40 \U712_CHIP_RAM.N_337_i_LC_14_20_2  (
            .in0(N__11368),
            .in1(N__11437),
            .in2(N__11140),
            .in3(N__11255),
            .lcout(N_337_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.N_336_i_LC_14_20_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.N_336_i_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.N_336_i_LC_14_20_4 .LUT_INIT=16'b0000111011100000;
    LogicCell40 \U712_CHIP_RAM.N_336_i_LC_14_20_4  (
            .in0(N__11367),
            .in1(N__11436),
            .in2(N__11139),
            .in3(N__11254),
            .lcout(N_336_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.N_335_i_LC_14_20_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.N_335_i_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.N_335_i_LC_14_20_6 .LUT_INIT=16'b0000001101110000;
    LogicCell40 \U712_CHIP_RAM.N_335_i_LC_14_20_6  (
            .in0(N__11366),
            .in1(N__11435),
            .in2(N__11138),
            .in3(N__11253),
            .lcout(N_335_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.N_334_i_LC_14_20_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.N_334_i_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.N_334_i_LC_14_20_7 .LUT_INIT=16'b0000101110100000;
    LogicCell40 \U712_CHIP_RAM.N_334_i_LC_14_20_7  (
            .in0(N__11434),
            .in1(N__11365),
            .in2(N__11264),
            .in3(N__11119),
            .lcout(N_334_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_7_3  (
            .in0(N__10773),
            .in1(N__10996),
            .in2(_gnd_net_),
            .in3(N__10949),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10631),
            .ce(N__10609),
            .sr(N__10524));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_8_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_15_8_6  (
            .in0(N__10911),
            .in1(N__10839),
            .in2(_gnd_net_),
            .in3(N__10687),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10629),
            .ce(N__10608),
            .sr(N__10518));
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_1 .LUT_INIT=16'b0100000001111111;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_1  (
            .in0(N__10390),
            .in1(N__10274),
            .in2(N__11840),
            .in3(N__11764),
            .lcout(N_379),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 30 2025 11:26:14

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4230\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \N_812_i\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \U712_REG_SM.N_266_cascade_\ : std_logic;
signal \U712_REG_SM.N_269_cascade_\ : std_logic;
signal \U712_REG_SM.N_233\ : std_logic;
signal \U712_REG_SM.N_191_cascade_\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.N_85\ : std_logic;
signal \U712_REG_SM.N_263\ : std_logic;
signal \U712_REG_SM.N_209\ : std_logic;
signal \U712_REG_SM.STATE_COUNTc_1_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_272_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_srsts_i_0_a5_0_0_0\ : std_logic;
signal \U712_REG_SM.N_207\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_191\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_0\ : std_logic;
signal \U712_REG_SM.DS_EN_RNOZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a5_0_0_0\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_i_i_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_i_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_23\ : std_logic;
signal \U712_REG_SM.N_219\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_261\ : std_logic;
signal \U712_BYTE_ENABLE.N_215_cascade_\ : std_logic;
signal \N_167_i\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_219_0_0\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \N_165_i\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_CHIP_RAM.N_279_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_187_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_316_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_316\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a5_1\ : std_logic;
signal \U712_CHIP_RAM.N_283_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_258\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_\ : std_logic;
signal \N_235\ : std_logic;
signal \RnW_c\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_222\ : std_logic;
signal \U712_BYTE_ENABLE.N_217\ : std_logic;
signal \DMA_LATCH_EN_c\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_10\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.N_340\ : std_logic;
signal \U712_CHIP_RAM.N_340_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_97\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.N_312\ : std_logic;
signal \U712_CHIP_RAM.N_206_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_329\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_323_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_374\ : std_logic;
signal \U712_CHIP_RAM.N_378\ : std_logic;
signal \U712_CHIP_RAM.N_184\ : std_logic;
signal \U712_CHIP_RAM.N_335_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_280\ : std_logic;
signal \U712_CHIP_RAM.N_284\ : std_logic;
signal \U712_CHIP_RAM.N_284_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_218\ : std_logic;
signal \U712_CHIP_RAM.N_218_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_259\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a2_0_a5_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_i_a5_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_257_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_i_0\ : std_logic;
signal \U712_CHIP_RAM.N_338_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_284_2\ : std_logic;
signal \U712_CHIP_RAM.N_253\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.N_284_2_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_254\ : std_logic;
signal \U712_CHIP_RAM.N_322\ : std_logic;
signal \U712_CHIP_RAM.N_206\ : std_logic;
signal \U712_CHIP_RAM.N_338\ : std_logic;
signal \U712_CHIP_RAM.N_256\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.N_211_i_0_en_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_211_i_0_en_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_339_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_335\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_296\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_181\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.N_289_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_288\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a5_0\ : std_logic;
signal \U712_CHIP_RAM.N_186\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0\ : std_logic;
signal \U712_CHIP_RAM.N_341\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_331\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.N_331_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_337\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.un3_DMA_CYCLE_START\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \A_c_7\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \U712_CHIP_RAM.N_327\ : std_logic;
signal \U712_CHIP_RAM.N_339\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \WRITE_CYCLEm\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\ : std_logic;
signal \N_118_i\ : std_logic;
signal \N_119_i\ : std_logic;
signal \U712_CHIP_RAM.N_323\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_a5_0_1_0\ : std_logic;
signal \U712_CHIP_RAM.N_287\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_a5_0Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.UUBE\ : std_logic;
signal \U712_BYTE_ENABLE.N_216\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \N_163\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_146\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_6_0_a5_2\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \DS_ENm\ : std_logic;
signal \U712_BYTE_ENABLE_un1_UDSn_i\ : std_logic;
signal \WEn_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_BYTE_ENABLE_UUBE_i\ : std_logic;
signal \N_215_i\ : std_logic;
signal \N_217_i\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \N_216_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \RASn_c\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__3939\,
            RESETB => \N__6459\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11659\,
            DIN => \N__11658\,
            DOUT => \N__11657\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11659\,
            PADOUT => \N__11658\,
            PADIN => \N__11657\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7002\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11650\,
            DIN => \N__11649\,
            DOUT => \N__11648\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11650\,
            PADOUT => \N__11649\,
            PADIN => \N__11648\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11641\,
            DIN => \N__11640\,
            DOUT => \N__11639\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11641\,
            PADOUT => \N__11640\,
            PADIN => \N__11639\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8514\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11632\,
            DIN => \N__11631\,
            DOUT => \N__11630\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11632\,
            PADOUT => \N__11631\,
            PADIN => \N__11630\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5034\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11623\,
            DIN => \N__11622\,
            DOUT => \N__11621\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11623\,
            PADOUT => \N__11622\,
            PADIN => \N__11621\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11614\,
            DIN => \N__11613\,
            DOUT => \N__11612\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11614\,
            PADOUT => \N__11613\,
            PADIN => \N__11612\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11605\,
            DIN => \N__11604\,
            DOUT => \N__11603\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11605\,
            PADOUT => \N__11604\,
            PADIN => \N__11603\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11596\,
            DIN => \N__11595\,
            DOUT => \N__11594\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11596\,
            PADOUT => \N__11595\,
            PADIN => \N__11594\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11587\,
            DIN => \N__11586\,
            DOUT => \N__11585\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11587\,
            PADOUT => \N__11586\,
            PADIN => \N__11585\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11578\,
            DIN => \N__11577\,
            DOUT => \N__11576\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11578\,
            PADOUT => \N__11577\,
            PADIN => \N__11576\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11569\,
            DIN => \N__11568\,
            DOUT => \N__11567\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11569\,
            PADOUT => \N__11568\,
            PADIN => \N__11567\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7914\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11560\,
            DIN => \N__11559\,
            DOUT => \N__11558\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11560\,
            PADOUT => \N__11559\,
            PADIN => \N__11558\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8895\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11551\,
            DIN => \N__11550\,
            DOUT => \N__11549\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11551\,
            PADOUT => \N__11550\,
            PADIN => \N__11549\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11542\,
            DIN => \N__11541\,
            DOUT => \N__11540\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11542\,
            PADOUT => \N__11541\,
            PADIN => \N__11540\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11533\,
            DIN => \N__11532\,
            DOUT => \N__11531\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11533\,
            PADOUT => \N__11532\,
            PADIN => \N__11531\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11524\,
            DIN => \N__11523\,
            DOUT => \N__11522\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11524\,
            PADOUT => \N__11523\,
            PADIN => \N__11522\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4239\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11515\,
            DIN => \N__11514\,
            DOUT => \N__11513\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11515\,
            PADOUT => \N__11514\,
            PADIN => \N__11513\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11506\,
            DIN => \N__11505\,
            DOUT => \N__11504\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11506\,
            PADOUT => \N__11505\,
            PADIN => \N__11504\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11497\,
            DIN => \N__11496\,
            DOUT => \N__11495\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11497\,
            PADOUT => \N__11496\,
            PADIN => \N__11495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7935\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11488\,
            DIN => \N__11487\,
            DOUT => \N__11486\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11488\,
            PADOUT => \N__11487\,
            PADIN => \N__11486\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11479\,
            DIN => \N__11478\,
            DOUT => \N__11477\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11479\,
            PADOUT => \N__11478\,
            PADIN => \N__11477\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8496\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11470\,
            DIN => \N__11469\,
            DOUT => \N__11468\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11470\,
            PADOUT => \N__11469\,
            PADIN => \N__11468\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11461\,
            DIN => \N__11460\,
            DOUT => \N__11459\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11461\,
            PADOUT => \N__11460\,
            PADIN => \N__11459\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8880\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11452\,
            DIN => \N__11451\,
            DOUT => \N__11450\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11452\,
            PADOUT => \N__11451\,
            PADIN => \N__11450\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11443\,
            DIN => \N__11442\,
            DOUT => \N__11441\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11443\,
            PADOUT => \N__11442\,
            PADIN => \N__11441\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11434\,
            DIN => \N__11433\,
            DOUT => \N__11432\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11434\,
            PADOUT => \N__11433\,
            PADIN => \N__11432\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11425\,
            DIN => \N__11424\,
            DOUT => \N__11423\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11425\,
            PADOUT => \N__11424\,
            PADIN => \N__11423\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11416\,
            DIN => \N__11415\,
            DOUT => \N__11414\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11416\,
            PADOUT => \N__11415\,
            PADIN => \N__11414\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11407\,
            DIN => \N__11406\,
            DOUT => \N__11405\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11407\,
            PADOUT => \N__11406\,
            PADIN => \N__11405\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4923\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11398\,
            DIN => \N__11397\,
            DOUT => \N__11396\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11398\,
            PADOUT => \N__11397\,
            PADIN => \N__11396\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11389\,
            DIN => \N__11388\,
            DOUT => \N__11387\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11389\,
            PADOUT => \N__11388\,
            PADIN => \N__11387\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11380\,
            DIN => \N__11379\,
            DOUT => \N__11378\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11380\,
            PADOUT => \N__11379\,
            PADIN => \N__11378\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11371\,
            DIN => \N__11370\,
            DOUT => \N__11369\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11371\,
            PADOUT => \N__11370\,
            PADIN => \N__11369\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11362\,
            DIN => \N__11361\,
            DOUT => \N__11360\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11362\,
            PADOUT => \N__11361\,
            PADIN => \N__11360\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6810\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11353\,
            DIN => \N__11352\,
            DOUT => \N__11351\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11353\,
            PADOUT => \N__11352\,
            PADIN => \N__11351\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11344\,
            DIN => \N__11343\,
            DOUT => \N__11342\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11344\,
            PADOUT => \N__11343\,
            PADIN => \N__11342\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9684\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11335\,
            DIN => \N__11334\,
            DOUT => \N__11333\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11335\,
            PADOUT => \N__11334\,
            PADIN => \N__11333\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11326\,
            DIN => \N__11325\,
            DOUT => \N__11324\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11326\,
            PADOUT => \N__11325\,
            PADIN => \N__11324\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6327\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11317\,
            DIN => \N__11316\,
            DOUT => \N__11315\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11317\,
            PADOUT => \N__11316\,
            PADIN => \N__11315\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6806\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11308\,
            DIN => \N__11307\,
            DOUT => \N__11306\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11308\,
            PADOUT => \N__11307\,
            PADIN => \N__11306\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3954\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11299\,
            DIN => \N__11298\,
            DOUT => \N__11297\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11299\,
            PADOUT => \N__11298\,
            PADIN => \N__11297\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11290\,
            DIN => \N__11289\,
            DOUT => \N__11288\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11290\,
            PADOUT => \N__11289\,
            PADIN => \N__11288\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4677\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11281\,
            DIN => \N__11280\,
            DOUT => \N__11279\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11281\,
            PADOUT => \N__11280\,
            PADIN => \N__11279\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6399\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11272\,
            DIN => \N__11271\,
            DOUT => \N__11270\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11272\,
            PADOUT => \N__11271\,
            PADIN => \N__11270\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11263\,
            DIN => \N__11262\,
            DOUT => \N__11261\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11263\,
            PADOUT => \N__11262\,
            PADIN => \N__11261\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11254\,
            DIN => \N__11253\,
            DOUT => \N__11252\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11254\,
            PADOUT => \N__11253\,
            PADIN => \N__11252\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11245\,
            DIN => \N__11244\,
            DOUT => \N__11243\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11245\,
            PADOUT => \N__11244\,
            PADIN => \N__11243\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11236\,
            DIN => \N__11235\,
            DOUT => \N__11234\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11236\,
            PADOUT => \N__11235\,
            PADIN => \N__11234\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8328\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11227\,
            DIN => \N__11226\,
            DOUT => \N__11225\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11227\,
            PADOUT => \N__11226\,
            PADIN => \N__11225\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11218\,
            DIN => \N__11217\,
            DOUT => \N__11216\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11218\,
            PADOUT => \N__11217\,
            PADIN => \N__11216\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6805\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11209\,
            DIN => \N__11208\,
            DOUT => \N__11207\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11209\,
            PADOUT => \N__11208\,
            PADIN => \N__11207\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8304\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11200\,
            DIN => \N__11199\,
            DOUT => \N__11198\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11200\,
            PADOUT => \N__11199\,
            PADIN => \N__11198\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10476\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11191\,
            DIN => \N__11190\,
            DOUT => \N__11189\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11191\,
            PADOUT => \N__11190\,
            PADIN => \N__11189\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4746\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11182\,
            DIN => \N__11181\,
            DOUT => \N__11180\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11182\,
            PADOUT => \N__11181\,
            PADIN => \N__11180\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8106\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11173\,
            DIN => \N__11172\,
            DOUT => \N__11171\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11173\,
            PADOUT => \N__11172\,
            PADIN => \N__11171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4673\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11164\,
            DIN => \N__11163\,
            DOUT => \N__11162\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11164\,
            PADOUT => \N__11163\,
            PADIN => \N__11162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11155\,
            DIN => \N__11154\,
            DOUT => \N__11153\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11155\,
            PADOUT => \N__11154\,
            PADIN => \N__11153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11146\,
            DIN => \N__11145\,
            DOUT => \N__11144\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11146\,
            PADOUT => \N__11145\,
            PADIN => \N__11144\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4521\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11137\,
            DIN => \N__11136\,
            DOUT => \N__11135\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11137\,
            PADOUT => \N__11136\,
            PADIN => \N__11135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8535\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11128\,
            DIN => \N__11127\,
            DOUT => \N__11126\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11128\,
            PADOUT => \N__11127\,
            PADIN => \N__11126\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4587\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11119\,
            DIN => \N__11118\,
            DOUT => \N__11117\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11119\,
            PADOUT => \N__11118\,
            PADIN => \N__11117\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7308\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11110\,
            DIN => \N__11109\,
            DOUT => \N__11108\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11110\,
            PADOUT => \N__11109\,
            PADIN => \N__11108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11101\,
            DIN => \N__11100\,
            DOUT => \N__11099\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11101\,
            PADOUT => \N__11100\,
            PADIN => \N__11099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11092\,
            DIN => \N__11091\,
            DOUT => \N__11090\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11092\,
            PADOUT => \N__11091\,
            PADIN => \N__11090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11083\,
            DIN => \N__11082\,
            DOUT => \N__11081\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11083\,
            PADOUT => \N__11082\,
            PADIN => \N__11081\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11074\,
            DIN => \N__11073\,
            DOUT => \N__11072\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11074\,
            PADOUT => \N__11073\,
            PADIN => \N__11072\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6435\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11065\,
            DIN => \N__11064\,
            DOUT => \N__11063\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11065\,
            PADOUT => \N__11064\,
            PADIN => \N__11063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8865\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11056\,
            DIN => \N__11055\,
            DOUT => \N__11054\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11056\,
            PADOUT => \N__11055\,
            PADIN => \N__11054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11047\,
            DIN => \N__11046\,
            DOUT => \N__11045\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11047\,
            PADOUT => \N__11046\,
            PADIN => \N__11045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7332\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11038\,
            DIN => \N__11037\,
            DOUT => \N__11036\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11038\,
            PADOUT => \N__11037\,
            PADIN => \N__11036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4014\,
            DIN0 => OPEN,
            DOUT0 => \N__4545\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11029\,
            DIN => \N__11028\,
            DOUT => \N__11027\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11029\,
            PADOUT => \N__11028\,
            PADIN => \N__11027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6417\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11020\,
            DIN => \N__11019\,
            DOUT => \N__11018\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11020\,
            PADOUT => \N__11019\,
            PADIN => \N__11018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11011\,
            DIN => \N__11010\,
            DOUT => \N__11009\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11011\,
            PADOUT => \N__11010\,
            PADIN => \N__11009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11002\,
            DIN => \N__11001\,
            DOUT => \N__11000\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11002\,
            PADOUT => \N__11001\,
            PADIN => \N__11000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7542\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10993\,
            DIN => \N__10992\,
            DOUT => \N__10991\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10993\,
            PADOUT => \N__10992\,
            PADIN => \N__10991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10984\,
            DIN => \N__10983\,
            DOUT => \N__10982\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10984\,
            PADOUT => \N__10983\,
            PADIN => \N__10982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10975\,
            DIN => \N__10974\,
            DOUT => \N__10973\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10975\,
            PADOUT => \N__10974\,
            PADIN => \N__10973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10966\,
            DIN => \N__10965\,
            DOUT => \N__10964\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10966\,
            PADOUT => \N__10965\,
            PADIN => \N__10964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10957\,
            DIN => \N__10956\,
            DOUT => \N__10955\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10957\,
            PADOUT => \N__10956\,
            PADIN => \N__10955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7500\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10948\,
            DIN => \N__10947\,
            DOUT => \N__10946\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10948\,
            PADOUT => \N__10947\,
            PADIN => \N__10946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7803\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10939\,
            DIN => \N__10938\,
            DOUT => \N__10937\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10939\,
            PADOUT => \N__10938\,
            PADIN => \N__10937\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9783\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10930\,
            DIN => \N__10929\,
            DOUT => \N__10928\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10930\,
            PADOUT => \N__10929\,
            PADIN => \N__10928\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7881\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10921\,
            DIN => \N__10920\,
            DOUT => \N__10919\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10921\,
            PADOUT => \N__10920\,
            PADIN => \N__10919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10912\,
            DIN => \N__10911\,
            DOUT => \N__10910\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10912\,
            PADOUT => \N__10911\,
            PADIN => \N__10910\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10903\,
            DIN => \N__10902\,
            DOUT => \N__10901\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10903\,
            PADOUT => \N__10902\,
            PADIN => \N__10901\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8169\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10894\,
            DIN => \N__10893\,
            DOUT => \N__10892\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10894\,
            PADOUT => \N__10893\,
            PADIN => \N__10892\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10885\,
            DIN => \N__10884\,
            DOUT => \N__10883\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10885\,
            PADOUT => \N__10884\,
            PADIN => \N__10883\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10876\,
            DIN => \N__10875\,
            DOUT => \N__10874\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10876\,
            PADOUT => \N__10875\,
            PADIN => \N__10874\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5178\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10867\,
            DIN => \N__10866\,
            DOUT => \N__10865\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10867\,
            PADOUT => \N__10866\,
            PADIN => \N__10865\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7578\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2647\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10839\
        );

    \I__2646\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10836\
        );

    \I__2645\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10833\
        );

    \I__2644\ : InMux
    port map (
            O => \N__10845\,
            I => \N__10830\
        );

    \I__2643\ : InMux
    port map (
            O => \N__10844\,
            I => \N__10823\
        );

    \I__2642\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10823\
        );

    \I__2641\ : InMux
    port map (
            O => \N__10842\,
            I => \N__10823\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__10839\,
            I => \N__10809\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__10836\,
            I => \N__10795\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__10833\,
            I => \N__10792\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__10830\,
            I => \N__10780\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__10823\,
            I => \N__10777\
        );

    \I__2635\ : SRMux
    port map (
            O => \N__10822\,
            I => \N__10680\
        );

    \I__2634\ : SRMux
    port map (
            O => \N__10821\,
            I => \N__10680\
        );

    \I__2633\ : SRMux
    port map (
            O => \N__10820\,
            I => \N__10680\
        );

    \I__2632\ : SRMux
    port map (
            O => \N__10819\,
            I => \N__10680\
        );

    \I__2631\ : SRMux
    port map (
            O => \N__10818\,
            I => \N__10680\
        );

    \I__2630\ : SRMux
    port map (
            O => \N__10817\,
            I => \N__10680\
        );

    \I__2629\ : SRMux
    port map (
            O => \N__10816\,
            I => \N__10680\
        );

    \I__2628\ : SRMux
    port map (
            O => \N__10815\,
            I => \N__10680\
        );

    \I__2627\ : SRMux
    port map (
            O => \N__10814\,
            I => \N__10680\
        );

    \I__2626\ : SRMux
    port map (
            O => \N__10813\,
            I => \N__10680\
        );

    \I__2625\ : SRMux
    port map (
            O => \N__10812\,
            I => \N__10680\
        );

    \I__2624\ : Glb2LocalMux
    port map (
            O => \N__10809\,
            I => \N__10680\
        );

    \I__2623\ : SRMux
    port map (
            O => \N__10808\,
            I => \N__10680\
        );

    \I__2622\ : SRMux
    port map (
            O => \N__10807\,
            I => \N__10680\
        );

    \I__2621\ : SRMux
    port map (
            O => \N__10806\,
            I => \N__10680\
        );

    \I__2620\ : SRMux
    port map (
            O => \N__10805\,
            I => \N__10680\
        );

    \I__2619\ : SRMux
    port map (
            O => \N__10804\,
            I => \N__10680\
        );

    \I__2618\ : SRMux
    port map (
            O => \N__10803\,
            I => \N__10680\
        );

    \I__2617\ : SRMux
    port map (
            O => \N__10802\,
            I => \N__10680\
        );

    \I__2616\ : SRMux
    port map (
            O => \N__10801\,
            I => \N__10680\
        );

    \I__2615\ : SRMux
    port map (
            O => \N__10800\,
            I => \N__10680\
        );

    \I__2614\ : SRMux
    port map (
            O => \N__10799\,
            I => \N__10680\
        );

    \I__2613\ : SRMux
    port map (
            O => \N__10798\,
            I => \N__10680\
        );

    \I__2612\ : Glb2LocalMux
    port map (
            O => \N__10795\,
            I => \N__10680\
        );

    \I__2611\ : Glb2LocalMux
    port map (
            O => \N__10792\,
            I => \N__10680\
        );

    \I__2610\ : SRMux
    port map (
            O => \N__10791\,
            I => \N__10680\
        );

    \I__2609\ : SRMux
    port map (
            O => \N__10790\,
            I => \N__10680\
        );

    \I__2608\ : SRMux
    port map (
            O => \N__10789\,
            I => \N__10680\
        );

    \I__2607\ : SRMux
    port map (
            O => \N__10788\,
            I => \N__10680\
        );

    \I__2606\ : SRMux
    port map (
            O => \N__10787\,
            I => \N__10680\
        );

    \I__2605\ : SRMux
    port map (
            O => \N__10786\,
            I => \N__10680\
        );

    \I__2604\ : SRMux
    port map (
            O => \N__10785\,
            I => \N__10680\
        );

    \I__2603\ : SRMux
    port map (
            O => \N__10784\,
            I => \N__10680\
        );

    \I__2602\ : SRMux
    port map (
            O => \N__10783\,
            I => \N__10680\
        );

    \I__2601\ : Glb2LocalMux
    port map (
            O => \N__10780\,
            I => \N__10680\
        );

    \I__2600\ : Glb2LocalMux
    port map (
            O => \N__10777\,
            I => \N__10680\
        );

    \I__2599\ : SRMux
    port map (
            O => \N__10776\,
            I => \N__10680\
        );

    \I__2598\ : SRMux
    port map (
            O => \N__10775\,
            I => \N__10680\
        );

    \I__2597\ : SRMux
    port map (
            O => \N__10774\,
            I => \N__10680\
        );

    \I__2596\ : SRMux
    port map (
            O => \N__10773\,
            I => \N__10680\
        );

    \I__2595\ : SRMux
    port map (
            O => \N__10772\,
            I => \N__10680\
        );

    \I__2594\ : SRMux
    port map (
            O => \N__10771\,
            I => \N__10680\
        );

    \I__2593\ : SRMux
    port map (
            O => \N__10770\,
            I => \N__10680\
        );

    \I__2592\ : SRMux
    port map (
            O => \N__10769\,
            I => \N__10680\
        );

    \I__2591\ : GlobalMux
    port map (
            O => \N__10680\,
            I => \N__10677\
        );

    \I__2590\ : gio2CtrlBuf
    port map (
            O => \N__10677\,
            I => \RESETn_c_i_g\
        );

    \I__2589\ : InMux
    port map (
            O => \N__10674\,
            I => \N__10670\
        );

    \I__2588\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10667\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__10670\,
            I => \N__10663\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__10667\,
            I => \N__10660\
        );

    \I__2585\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10657\
        );

    \I__2584\ : Span12Mux_v
    port map (
            O => \N__10663\,
            I => \N__10654\
        );

    \I__2583\ : Span4Mux_h
    port map (
            O => \N__10660\,
            I => \N__10650\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__10657\,
            I => \N__10647\
        );

    \I__2581\ : Span12Mux_h
    port map (
            O => \N__10654\,
            I => \N__10644\
        );

    \I__2580\ : InMux
    port map (
            O => \N__10653\,
            I => \N__10641\
        );

    \I__2579\ : Span4Mux_v
    port map (
            O => \N__10650\,
            I => \N__10636\
        );

    \I__2578\ : Span4Mux_h
    port map (
            O => \N__10647\,
            I => \N__10636\
        );

    \I__2577\ : Odrv12
    port map (
            O => \N__10644\,
            I => \REG_CYCLEm\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__10641\,
            I => \REG_CYCLEm\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__10636\,
            I => \REG_CYCLEm\
        );

    \I__2574\ : InMux
    port map (
            O => \N__10629\,
            I => \N__10625\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__10628\,
            I => \N__10621\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__10625\,
            I => \N__10617\
        );

    \I__2571\ : InMux
    port map (
            O => \N__10624\,
            I => \N__10614\
        );

    \I__2570\ : InMux
    port map (
            O => \N__10621\,
            I => \N__10611\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__10620\,
            I => \N__10608\
        );

    \I__2568\ : Span4Mux_v
    port map (
            O => \N__10617\,
            I => \N__10603\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__10614\,
            I => \N__10603\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__10611\,
            I => \N__10600\
        );

    \I__2565\ : InMux
    port map (
            O => \N__10608\,
            I => \N__10597\
        );

    \I__2564\ : Span4Mux_v
    port map (
            O => \N__10603\,
            I => \N__10593\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__10600\,
            I => \N__10588\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__10597\,
            I => \N__10588\
        );

    \I__2561\ : InMux
    port map (
            O => \N__10596\,
            I => \N__10585\
        );

    \I__2560\ : Span4Mux_h
    port map (
            O => \N__10593\,
            I => \N__10582\
        );

    \I__2559\ : Span4Mux_v
    port map (
            O => \N__10588\,
            I => \N__10576\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__10585\,
            I => \N__10576\
        );

    \I__2557\ : Span4Mux_h
    port map (
            O => \N__10582\,
            I => \N__10573\
        );

    \I__2556\ : InMux
    port map (
            O => \N__10581\,
            I => \N__10570\
        );

    \I__2555\ : Sp12to4
    port map (
            O => \N__10576\,
            I => \N__10567\
        );

    \I__2554\ : Span4Mux_h
    port map (
            O => \N__10573\,
            I => \N__10562\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__10570\,
            I => \N__10562\
        );

    \I__2552\ : Span12Mux_v
    port map (
            O => \N__10567\,
            I => \N__10559\
        );

    \I__2551\ : Span4Mux_h
    port map (
            O => \N__10562\,
            I => \N__10556\
        );

    \I__2550\ : Span12Mux_h
    port map (
            O => \N__10559\,
            I => \N__10553\
        );

    \I__2549\ : Span4Mux_v
    port map (
            O => \N__10556\,
            I => \N__10550\
        );

    \I__2548\ : Odrv12
    port map (
            O => \N__10553\,
            I => \CASUn_c\
        );

    \I__2547\ : Odrv4
    port map (
            O => \N__10550\,
            I => \CASUn_c\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__10545\,
            I => \N__10540\
        );

    \I__2545\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10537\
        );

    \I__2544\ : InMux
    port map (
            O => \N__10543\,
            I => \N__10534\
        );

    \I__2543\ : InMux
    port map (
            O => \N__10540\,
            I => \N__10531\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__10537\,
            I => \N__10525\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__10534\,
            I => \N__10525\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__10531\,
            I => \N__10522\
        );

    \I__2539\ : InMux
    port map (
            O => \N__10530\,
            I => \N__10519\
        );

    \I__2538\ : Span4Mux_v
    port map (
            O => \N__10525\,
            I => \N__10511\
        );

    \I__2537\ : Span4Mux_v
    port map (
            O => \N__10522\,
            I => \N__10511\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10519\,
            I => \N__10511\
        );

    \I__2535\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10508\
        );

    \I__2534\ : Span4Mux_h
    port map (
            O => \N__10511\,
            I => \N__10503\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10508\,
            I => \N__10503\
        );

    \I__2532\ : Span4Mux_v
    port map (
            O => \N__10503\,
            I => \N__10500\
        );

    \I__2531\ : Span4Mux_v
    port map (
            O => \N__10500\,
            I => \N__10496\
        );

    \I__2530\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10493\
        );

    \I__2529\ : Sp12to4
    port map (
            O => \N__10496\,
            I => \N__10490\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__10493\,
            I => \N__10487\
        );

    \I__2527\ : Span12Mux_h
    port map (
            O => \N__10490\,
            I => \N__10484\
        );

    \I__2526\ : Span12Mux_v
    port map (
            O => \N__10487\,
            I => \N__10481\
        );

    \I__2525\ : Odrv12
    port map (
            O => \N__10484\,
            I => \CASLn_c\
        );

    \I__2524\ : Odrv12
    port map (
            O => \N__10481\,
            I => \CASLn_c\
        );

    \I__2523\ : IoInMux
    port map (
            O => \N__10476\,
            I => \N__10473\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__10473\,
            I => \N__10470\
        );

    \I__2521\ : Span12Mux_s7_v
    port map (
            O => \N__10470\,
            I => \N__10467\
        );

    \I__2520\ : Odrv12
    port map (
            O => \N__10467\,
            I => \DRDENn_c\
        );

    \I__2519\ : InMux
    port map (
            O => \N__10464\,
            I => \N__10461\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__10461\,
            I => \N__10457\
        );

    \I__2517\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10454\
        );

    \I__2516\ : Span12Mux_h
    port map (
            O => \N__10457\,
            I => \N__10451\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__10454\,
            I => \N__10448\
        );

    \I__2514\ : Odrv12
    port map (
            O => \N__10451\,
            I => \DBRn_c_i\
        );

    \I__2513\ : Odrv4
    port map (
            O => \N__10448\,
            I => \DBRn_c_i\
        );

    \I__2512\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10439\
        );

    \I__2511\ : InMux
    port map (
            O => \N__10442\,
            I => \N__10436\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10439\,
            I => \N__10433\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__10436\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2508\ : Odrv12
    port map (
            O => \N__10433\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2507\ : InMux
    port map (
            O => \N__10428\,
            I => \N__10425\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__10425\,
            I => \N__10422\
        );

    \I__2505\ : Span4Mux_v
    port map (
            O => \N__10422\,
            I => \N__10419\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__10419\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2503\ : InMux
    port map (
            O => \N__10416\,
            I => \N__10409\
        );

    \I__2502\ : InMux
    port map (
            O => \N__10415\,
            I => \N__10409\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10405\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__10409\,
            I => \N__10402\
        );

    \I__2499\ : InMux
    port map (
            O => \N__10408\,
            I => \N__10399\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__10405\,
            I => \N__10396\
        );

    \I__2497\ : Span4Mux_v
    port map (
            O => \N__10402\,
            I => \N__10391\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10399\,
            I => \N__10391\
        );

    \I__2495\ : Span4Mux_v
    port map (
            O => \N__10396\,
            I => \N__10388\
        );

    \I__2494\ : Span4Mux_h
    port map (
            O => \N__10391\,
            I => \N__10385\
        );

    \I__2493\ : Span4Mux_v
    port map (
            O => \N__10388\,
            I => \N__10382\
        );

    \I__2492\ : Span4Mux_v
    port map (
            O => \N__10385\,
            I => \N__10379\
        );

    \I__2491\ : Sp12to4
    port map (
            O => \N__10382\,
            I => \N__10374\
        );

    \I__2490\ : Sp12to4
    port map (
            O => \N__10379\,
            I => \N__10374\
        );

    \I__2489\ : Odrv12
    port map (
            O => \N__10374\,
            I => \DRA_c_5\
        );

    \I__2488\ : InMux
    port map (
            O => \N__10371\,
            I => \N__10366\
        );

    \I__2487\ : InMux
    port map (
            O => \N__10370\,
            I => \N__10363\
        );

    \I__2486\ : InMux
    port map (
            O => \N__10369\,
            I => \N__10359\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__10366\,
            I => \N__10354\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__10363\,
            I => \N__10354\
        );

    \I__2483\ : InMux
    port map (
            O => \N__10362\,
            I => \N__10351\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__10359\,
            I => \N__10344\
        );

    \I__2481\ : Span4Mux_v
    port map (
            O => \N__10354\,
            I => \N__10344\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__10351\,
            I => \N__10344\
        );

    \I__2479\ : Span4Mux_h
    port map (
            O => \N__10344\,
            I => \N__10341\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__10341\,
            I => \N__10338\
        );

    \I__2477\ : Sp12to4
    port map (
            O => \N__10338\,
            I => \N__10335\
        );

    \I__2476\ : Odrv12
    port map (
            O => \N__10335\,
            I => \DRA_c_6\
        );

    \I__2475\ : InMux
    port map (
            O => \N__10332\,
            I => \N__10329\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__10329\,
            I => \N__10326\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__10326\,
            I => \N__10323\
        );

    \I__2472\ : Odrv4
    port map (
            O => \N__10323\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2471\ : InMux
    port map (
            O => \N__10320\,
            I => \N__10314\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10314\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__10314\,
            I => \N__10310\
        );

    \I__2468\ : InMux
    port map (
            O => \N__10313\,
            I => \N__10307\
        );

    \I__2467\ : Span4Mux_h
    port map (
            O => \N__10310\,
            I => \N__10301\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10307\,
            I => \N__10301\
        );

    \I__2465\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10298\
        );

    \I__2464\ : Sp12to4
    port map (
            O => \N__10301\,
            I => \N__10293\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__10298\,
            I => \N__10293\
        );

    \I__2462\ : Span12Mux_v
    port map (
            O => \N__10293\,
            I => \N__10290\
        );

    \I__2461\ : Span12Mux_h
    port map (
            O => \N__10290\,
            I => \N__10287\
        );

    \I__2460\ : Odrv12
    port map (
            O => \N__10287\,
            I => \DRA_c_4\
        );

    \I__2459\ : InMux
    port map (
            O => \N__10284\,
            I => \N__10279\
        );

    \I__2458\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10276\
        );

    \I__2457\ : InMux
    port map (
            O => \N__10282\,
            I => \N__10272\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__10279\,
            I => \N__10267\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__10276\,
            I => \N__10267\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10264\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__10272\,
            I => \N__10261\
        );

    \I__2452\ : Span4Mux_v
    port map (
            O => \N__10267\,
            I => \N__10256\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__10264\,
            I => \N__10256\
        );

    \I__2450\ : Span4Mux_v
    port map (
            O => \N__10261\,
            I => \N__10253\
        );

    \I__2449\ : Span4Mux_h
    port map (
            O => \N__10256\,
            I => \N__10250\
        );

    \I__2448\ : Span4Mux_v
    port map (
            O => \N__10253\,
            I => \N__10247\
        );

    \I__2447\ : Span4Mux_v
    port map (
            O => \N__10250\,
            I => \N__10244\
        );

    \I__2446\ : Sp12to4
    port map (
            O => \N__10247\,
            I => \N__10239\
        );

    \I__2445\ : Sp12to4
    port map (
            O => \N__10244\,
            I => \N__10239\
        );

    \I__2444\ : Odrv12
    port map (
            O => \N__10239\,
            I => \DRA_c_3\
        );

    \I__2443\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10233\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__10233\,
            I => \N__10230\
        );

    \I__2441\ : Span4Mux_h
    port map (
            O => \N__10230\,
            I => \N__10227\
        );

    \I__2440\ : Span4Mux_h
    port map (
            O => \N__10227\,
            I => \N__10224\
        );

    \I__2439\ : Odrv4
    port map (
            O => \N__10224\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2438\ : InMux
    port map (
            O => \N__10221\,
            I => \N__10218\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10218\,
            I => \N__10215\
        );

    \I__2436\ : Span4Mux_h
    port map (
            O => \N__10215\,
            I => \N__10212\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__10212\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10209\,
            I => \N__10206\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__10206\,
            I => \N__10203\
        );

    \I__2432\ : Span4Mux_h
    port map (
            O => \N__10203\,
            I => \N__10200\
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__10200\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2430\ : InMux
    port map (
            O => \N__10197\,
            I => \N__10191\
        );

    \I__2429\ : InMux
    port map (
            O => \N__10196\,
            I => \N__10188\
        );

    \I__2428\ : InMux
    port map (
            O => \N__10195\,
            I => \N__10185\
        );

    \I__2427\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10182\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__10191\,
            I => \N__10173\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10188\,
            I => \N__10173\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__10185\,
            I => \N__10173\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__10182\,
            I => \N__10173\
        );

    \I__2422\ : Span12Mux_h
    port map (
            O => \N__10173\,
            I => \N__10170\
        );

    \I__2421\ : Odrv12
    port map (
            O => \N__10170\,
            I => \DRA_c_7\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10167\,
            I => \N__10161\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10166\,
            I => \N__10158\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10165\,
            I => \N__10155\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10152\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__10161\,
            I => \N__10149\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__10158\,
            I => \N__10142\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__10155\,
            I => \N__10142\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__10152\,
            I => \N__10142\
        );

    \I__2412\ : Span4Mux_v
    port map (
            O => \N__10149\,
            I => \N__10137\
        );

    \I__2411\ : Span4Mux_v
    port map (
            O => \N__10142\,
            I => \N__10137\
        );

    \I__2410\ : Sp12to4
    port map (
            O => \N__10137\,
            I => \N__10134\
        );

    \I__2409\ : Odrv12
    port map (
            O => \N__10134\,
            I => \DRA_c_8\
        );

    \I__2408\ : CascadeMux
    port map (
            O => \N__10131\,
            I => \N__10128\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10128\,
            I => \N__10125\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__10125\,
            I => \N__10122\
        );

    \I__2405\ : Odrv12
    port map (
            O => \N__10122\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2404\ : InMux
    port map (
            O => \N__10119\,
            I => \N__10115\
        );

    \I__2403\ : CascadeMux
    port map (
            O => \N__10118\,
            I => \N__10111\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__10115\,
            I => \N__10108\
        );

    \I__2401\ : InMux
    port map (
            O => \N__10114\,
            I => \N__10105\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10111\,
            I => \N__10102\
        );

    \I__2399\ : Span4Mux_h
    port map (
            O => \N__10108\,
            I => \N__10097\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__10105\,
            I => \N__10097\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__10102\,
            I => \N__10094\
        );

    \I__2396\ : Span4Mux_v
    port map (
            O => \N__10097\,
            I => \N__10090\
        );

    \I__2395\ : Span4Mux_v
    port map (
            O => \N__10094\,
            I => \N__10087\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10093\,
            I => \N__10084\
        );

    \I__2393\ : Sp12to4
    port map (
            O => \N__10090\,
            I => \N__10079\
        );

    \I__2392\ : Sp12to4
    port map (
            O => \N__10087\,
            I => \N__10079\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__10084\,
            I => \N__10076\
        );

    \I__2390\ : Span12Mux_h
    port map (
            O => \N__10079\,
            I => \N__10073\
        );

    \I__2389\ : Span12Mux_v
    port map (
            O => \N__10076\,
            I => \N__10070\
        );

    \I__2388\ : Span12Mux_v
    port map (
            O => \N__10073\,
            I => \N__10067\
        );

    \I__2387\ : Span12Mux_v
    port map (
            O => \N__10070\,
            I => \N__10064\
        );

    \I__2386\ : Odrv12
    port map (
            O => \N__10067\,
            I => \DRA_c_9\
        );

    \I__2385\ : Odrv12
    port map (
            O => \N__10064\,
            I => \DRA_c_9\
        );

    \I__2384\ : InMux
    port map (
            O => \N__10059\,
            I => \N__10056\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__10056\,
            I => \N__10053\
        );

    \I__2382\ : Odrv12
    port map (
            O => \N__10053\,
            I => \RAS0n_c\
        );

    \I__2381\ : InMux
    port map (
            O => \N__10050\,
            I => \N__10045\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__10049\,
            I => \N__10036\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__10048\,
            I => \N__10028\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10045\,
            I => \N__10023\
        );

    \I__2377\ : InMux
    port map (
            O => \N__10044\,
            I => \N__10018\
        );

    \I__2376\ : InMux
    port map (
            O => \N__10043\,
            I => \N__10018\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10042\,
            I => \N__10015\
        );

    \I__2374\ : InMux
    port map (
            O => \N__10041\,
            I => \N__10012\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10040\,
            I => \N__10008\
        );

    \I__2372\ : InMux
    port map (
            O => \N__10039\,
            I => \N__10001\
        );

    \I__2371\ : InMux
    port map (
            O => \N__10036\,
            I => \N__10001\
        );

    \I__2370\ : InMux
    port map (
            O => \N__10035\,
            I => \N__10001\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10034\,
            I => \N__9994\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10033\,
            I => \N__9994\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10032\,
            I => \N__9994\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10031\,
            I => \N__9989\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10028\,
            I => \N__9984\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10027\,
            I => \N__9984\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10026\,
            I => \N__9981\
        );

    \I__2362\ : Span4Mux_v
    port map (
            O => \N__10023\,
            I => \N__9974\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__10018\,
            I => \N__9974\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__10015\,
            I => \N__9974\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10012\,
            I => \N__9971\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10011\,
            I => \N__9968\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10008\,
            I => \N__9964\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__10001\,
            I => \N__9959\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__9994\,
            I => \N__9959\
        );

    \I__2354\ : InMux
    port map (
            O => \N__9993\,
            I => \N__9956\
        );

    \I__2353\ : InMux
    port map (
            O => \N__9992\,
            I => \N__9953\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__9989\,
            I => \N__9950\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__9984\,
            I => \N__9945\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__9981\,
            I => \N__9945\
        );

    \I__2349\ : Span4Mux_h
    port map (
            O => \N__9974\,
            I => \N__9939\
        );

    \I__2348\ : Span4Mux_v
    port map (
            O => \N__9971\,
            I => \N__9939\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__9968\,
            I => \N__9936\
        );

    \I__2346\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9933\
        );

    \I__2345\ : Span4Mux_v
    port map (
            O => \N__9964\,
            I => \N__9930\
        );

    \I__2344\ : Span4Mux_v
    port map (
            O => \N__9959\,
            I => \N__9923\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__9956\,
            I => \N__9923\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__9953\,
            I => \N__9923\
        );

    \I__2341\ : Span4Mux_v
    port map (
            O => \N__9950\,
            I => \N__9918\
        );

    \I__2340\ : Span4Mux_v
    port map (
            O => \N__9945\,
            I => \N__9918\
        );

    \I__2339\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9915\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__9939\,
            I => \N__9910\
        );

    \I__2337\ : Span4Mux_v
    port map (
            O => \N__9936\,
            I => \N__9910\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__9933\,
            I => \N__9907\
        );

    \I__2335\ : Span4Mux_h
    port map (
            O => \N__9930\,
            I => \N__9902\
        );

    \I__2334\ : Span4Mux_v
    port map (
            O => \N__9923\,
            I => \N__9902\
        );

    \I__2333\ : Sp12to4
    port map (
            O => \N__9918\,
            I => \N__9897\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__9915\,
            I => \N__9897\
        );

    \I__2331\ : Span4Mux_h
    port map (
            O => \N__9910\,
            I => \N__9894\
        );

    \I__2330\ : Span12Mux_v
    port map (
            O => \N__9907\,
            I => \N__9891\
        );

    \I__2329\ : Sp12to4
    port map (
            O => \N__9902\,
            I => \N__9888\
        );

    \I__2328\ : Span12Mux_h
    port map (
            O => \N__9897\,
            I => \N__9883\
        );

    \I__2327\ : Sp12to4
    port map (
            O => \N__9894\,
            I => \N__9883\
        );

    \I__2326\ : Span12Mux_h
    port map (
            O => \N__9891\,
            I => \N__9880\
        );

    \I__2325\ : Span12Mux_h
    port map (
            O => \N__9888\,
            I => \N__9877\
        );

    \I__2324\ : Span12Mux_v
    port map (
            O => \N__9883\,
            I => \N__9874\
        );

    \I__2323\ : Odrv12
    port map (
            O => \N__9880\,
            I => \AGNUS_REV_c\
        );

    \I__2322\ : Odrv12
    port map (
            O => \N__9877\,
            I => \AGNUS_REV_c\
        );

    \I__2321\ : Odrv12
    port map (
            O => \N__9874\,
            I => \AGNUS_REV_c\
        );

    \I__2320\ : InMux
    port map (
            O => \N__9867\,
            I => \N__9864\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__9864\,
            I => \N__9861\
        );

    \I__2318\ : Odrv12
    port map (
            O => \N__9861\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2317\ : ClkMux
    port map (
            O => \N__9858\,
            I => \N__9834\
        );

    \I__2316\ : ClkMux
    port map (
            O => \N__9857\,
            I => \N__9834\
        );

    \I__2315\ : ClkMux
    port map (
            O => \N__9856\,
            I => \N__9834\
        );

    \I__2314\ : ClkMux
    port map (
            O => \N__9855\,
            I => \N__9834\
        );

    \I__2313\ : ClkMux
    port map (
            O => \N__9854\,
            I => \N__9834\
        );

    \I__2312\ : ClkMux
    port map (
            O => \N__9853\,
            I => \N__9834\
        );

    \I__2311\ : ClkMux
    port map (
            O => \N__9852\,
            I => \N__9834\
        );

    \I__2310\ : ClkMux
    port map (
            O => \N__9851\,
            I => \N__9834\
        );

    \I__2309\ : GlobalMux
    port map (
            O => \N__9834\,
            I => \N__9831\
        );

    \I__2308\ : gio2CtrlBuf
    port map (
            O => \N__9831\,
            I => \C3_c_g\
        );

    \I__2307\ : CEMux
    port map (
            O => \N__9828\,
            I => \N__9789\
        );

    \I__2306\ : CEMux
    port map (
            O => \N__9827\,
            I => \N__9789\
        );

    \I__2305\ : CEMux
    port map (
            O => \N__9826\,
            I => \N__9789\
        );

    \I__2304\ : CEMux
    port map (
            O => \N__9825\,
            I => \N__9789\
        );

    \I__2303\ : CEMux
    port map (
            O => \N__9824\,
            I => \N__9789\
        );

    \I__2302\ : CEMux
    port map (
            O => \N__9823\,
            I => \N__9789\
        );

    \I__2301\ : CEMux
    port map (
            O => \N__9822\,
            I => \N__9789\
        );

    \I__2300\ : CEMux
    port map (
            O => \N__9821\,
            I => \N__9789\
        );

    \I__2299\ : CEMux
    port map (
            O => \N__9820\,
            I => \N__9789\
        );

    \I__2298\ : CEMux
    port map (
            O => \N__9819\,
            I => \N__9789\
        );

    \I__2297\ : CEMux
    port map (
            O => \N__9818\,
            I => \N__9789\
        );

    \I__2296\ : CEMux
    port map (
            O => \N__9817\,
            I => \N__9789\
        );

    \I__2295\ : CEMux
    port map (
            O => \N__9816\,
            I => \N__9789\
        );

    \I__2294\ : GlobalMux
    port map (
            O => \N__9789\,
            I => \N__9786\
        );

    \I__2293\ : gio2CtrlBuf
    port map (
            O => \N__9786\,
            I => \DBRn_c_i_0_g\
        );

    \I__2292\ : IoInMux
    port map (
            O => \N__9783\,
            I => \N__9780\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__9780\,
            I => \N__9777\
        );

    \I__2290\ : Span4Mux_s2_v
    port map (
            O => \N__9777\,
            I => \N__9774\
        );

    \I__2289\ : Span4Mux_h
    port map (
            O => \N__9774\,
            I => \N__9771\
        );

    \I__2288\ : Span4Mux_v
    port map (
            O => \N__9771\,
            I => \N__9768\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__9768\,
            I => \N_216_i\
        );

    \I__2286\ : InMux
    port map (
            O => \N__9765\,
            I => \N__9761\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__9764\,
            I => \N__9758\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__9761\,
            I => \N__9755\
        );

    \I__2283\ : InMux
    port map (
            O => \N__9758\,
            I => \N__9752\
        );

    \I__2282\ : Span4Mux_v
    port map (
            O => \N__9755\,
            I => \N__9744\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__9752\,
            I => \N__9744\
        );

    \I__2280\ : InMux
    port map (
            O => \N__9751\,
            I => \N__9741\
        );

    \I__2279\ : InMux
    port map (
            O => \N__9750\,
            I => \N__9738\
        );

    \I__2278\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9735\
        );

    \I__2277\ : Span4Mux_h
    port map (
            O => \N__9744\,
            I => \N__9730\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__9741\,
            I => \N__9727\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__9738\,
            I => \N__9722\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__9735\,
            I => \N__9722\
        );

    \I__2273\ : InMux
    port map (
            O => \N__9734\,
            I => \N__9719\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__9733\,
            I => \N__9716\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__9730\,
            I => \N__9713\
        );

    \I__2270\ : Span4Mux_v
    port map (
            O => \N__9727\,
            I => \N__9710\
        );

    \I__2269\ : Span4Mux_h
    port map (
            O => \N__9722\,
            I => \N__9705\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__9719\,
            I => \N__9705\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9702\
        );

    \I__2266\ : Span4Mux_h
    port map (
            O => \N__9713\,
            I => \N__9699\
        );

    \I__2265\ : Span4Mux_h
    port map (
            O => \N__9710\,
            I => \N__9696\
        );

    \I__2264\ : Span4Mux_h
    port map (
            O => \N__9705\,
            I => \N__9693\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__9702\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__9699\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__9696\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__9693\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2259\ : IoInMux
    port map (
            O => \N__9684\,
            I => \N__9681\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__9681\,
            I => \N__9678\
        );

    \I__2257\ : IoSpan4Mux
    port map (
            O => \N__9678\,
            I => \N__9675\
        );

    \I__2256\ : Span4Mux_s2_v
    port map (
            O => \N__9675\,
            I => \N__9672\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__9672\,
            I => \N__9669\
        );

    \I__2254\ : Span4Mux_v
    port map (
            O => \N__9669\,
            I => \N__9666\
        );

    \I__2253\ : Odrv4
    port map (
            O => \N__9666\,
            I => \RASn_c\
        );

    \I__2252\ : InMux
    port map (
            O => \N__9663\,
            I => \N__9660\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__9660\,
            I => \N__9626\
        );

    \I__2250\ : ClkMux
    port map (
            O => \N__9659\,
            I => \N__9531\
        );

    \I__2249\ : ClkMux
    port map (
            O => \N__9658\,
            I => \N__9531\
        );

    \I__2248\ : ClkMux
    port map (
            O => \N__9657\,
            I => \N__9531\
        );

    \I__2247\ : ClkMux
    port map (
            O => \N__9656\,
            I => \N__9531\
        );

    \I__2246\ : ClkMux
    port map (
            O => \N__9655\,
            I => \N__9531\
        );

    \I__2245\ : ClkMux
    port map (
            O => \N__9654\,
            I => \N__9531\
        );

    \I__2244\ : ClkMux
    port map (
            O => \N__9653\,
            I => \N__9531\
        );

    \I__2243\ : ClkMux
    port map (
            O => \N__9652\,
            I => \N__9531\
        );

    \I__2242\ : ClkMux
    port map (
            O => \N__9651\,
            I => \N__9531\
        );

    \I__2241\ : ClkMux
    port map (
            O => \N__9650\,
            I => \N__9531\
        );

    \I__2240\ : ClkMux
    port map (
            O => \N__9649\,
            I => \N__9531\
        );

    \I__2239\ : ClkMux
    port map (
            O => \N__9648\,
            I => \N__9531\
        );

    \I__2238\ : ClkMux
    port map (
            O => \N__9647\,
            I => \N__9531\
        );

    \I__2237\ : ClkMux
    port map (
            O => \N__9646\,
            I => \N__9531\
        );

    \I__2236\ : ClkMux
    port map (
            O => \N__9645\,
            I => \N__9531\
        );

    \I__2235\ : ClkMux
    port map (
            O => \N__9644\,
            I => \N__9531\
        );

    \I__2234\ : ClkMux
    port map (
            O => \N__9643\,
            I => \N__9531\
        );

    \I__2233\ : ClkMux
    port map (
            O => \N__9642\,
            I => \N__9531\
        );

    \I__2232\ : ClkMux
    port map (
            O => \N__9641\,
            I => \N__9531\
        );

    \I__2231\ : ClkMux
    port map (
            O => \N__9640\,
            I => \N__9531\
        );

    \I__2230\ : ClkMux
    port map (
            O => \N__9639\,
            I => \N__9531\
        );

    \I__2229\ : ClkMux
    port map (
            O => \N__9638\,
            I => \N__9531\
        );

    \I__2228\ : ClkMux
    port map (
            O => \N__9637\,
            I => \N__9531\
        );

    \I__2227\ : ClkMux
    port map (
            O => \N__9636\,
            I => \N__9531\
        );

    \I__2226\ : ClkMux
    port map (
            O => \N__9635\,
            I => \N__9531\
        );

    \I__2225\ : ClkMux
    port map (
            O => \N__9634\,
            I => \N__9531\
        );

    \I__2224\ : ClkMux
    port map (
            O => \N__9633\,
            I => \N__9531\
        );

    \I__2223\ : ClkMux
    port map (
            O => \N__9632\,
            I => \N__9531\
        );

    \I__2222\ : ClkMux
    port map (
            O => \N__9631\,
            I => \N__9531\
        );

    \I__2221\ : ClkMux
    port map (
            O => \N__9630\,
            I => \N__9531\
        );

    \I__2220\ : ClkMux
    port map (
            O => \N__9629\,
            I => \N__9531\
        );

    \I__2219\ : Glb2LocalMux
    port map (
            O => \N__9626\,
            I => \N__9531\
        );

    \I__2218\ : ClkMux
    port map (
            O => \N__9625\,
            I => \N__9531\
        );

    \I__2217\ : ClkMux
    port map (
            O => \N__9624\,
            I => \N__9531\
        );

    \I__2216\ : ClkMux
    port map (
            O => \N__9623\,
            I => \N__9531\
        );

    \I__2215\ : ClkMux
    port map (
            O => \N__9622\,
            I => \N__9531\
        );

    \I__2214\ : ClkMux
    port map (
            O => \N__9621\,
            I => \N__9531\
        );

    \I__2213\ : ClkMux
    port map (
            O => \N__9620\,
            I => \N__9531\
        );

    \I__2212\ : ClkMux
    port map (
            O => \N__9619\,
            I => \N__9531\
        );

    \I__2211\ : ClkMux
    port map (
            O => \N__9618\,
            I => \N__9531\
        );

    \I__2210\ : ClkMux
    port map (
            O => \N__9617\,
            I => \N__9531\
        );

    \I__2209\ : ClkMux
    port map (
            O => \N__9616\,
            I => \N__9531\
        );

    \I__2208\ : GlobalMux
    port map (
            O => \N__9531\,
            I => \CLK80_PLL\
        );

    \I__2207\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9522\
        );

    \I__2206\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9522\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__9522\,
            I => \N__9519\
        );

    \I__2204\ : Odrv12
    port map (
            O => \N__9519\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9516\,
            I => \N__9513\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__9513\,
            I => \N__9510\
        );

    \I__2201\ : Odrv4
    port map (
            O => \N__9510\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__9507\,
            I => \N__9504\
        );

    \I__2199\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9501\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__9501\,
            I => \N__9498\
        );

    \I__2197\ : Span4Mux_h
    port map (
            O => \N__9498\,
            I => \N__9495\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__9495\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9489\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__9489\,
            I => \N__9486\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__9486\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9480\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__9480\,
            I => \N__9477\
        );

    \I__2190\ : Span4Mux_h
    port map (
            O => \N__9477\,
            I => \N__9474\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__9474\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9468\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__9468\,
            I => \N__9465\
        );

    \I__2186\ : Span4Mux_h
    port map (
            O => \N__9465\,
            I => \N__9462\
        );

    \I__2185\ : Odrv4
    port map (
            O => \N__9462\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9459\,
            I => \N__9454\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9451\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9457\,
            I => \N__9448\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9454\,
            I => \N__9445\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__9451\,
            I => \N__9439\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9448\,
            I => \N__9439\
        );

    \I__2178\ : Span4Mux_v
    port map (
            O => \N__9445\,
            I => \N__9436\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9444\,
            I => \N__9433\
        );

    \I__2176\ : Span4Mux_h
    port map (
            O => \N__9439\,
            I => \N__9430\
        );

    \I__2175\ : Span4Mux_v
    port map (
            O => \N__9436\,
            I => \N__9427\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__9433\,
            I => \N__9424\
        );

    \I__2173\ : Sp12to4
    port map (
            O => \N__9430\,
            I => \N__9421\
        );

    \I__2172\ : Sp12to4
    port map (
            O => \N__9427\,
            I => \N__9416\
        );

    \I__2171\ : Span12Mux_v
    port map (
            O => \N__9424\,
            I => \N__9416\
        );

    \I__2170\ : Span12Mux_v
    port map (
            O => \N__9421\,
            I => \N__9413\
        );

    \I__2169\ : Span12Mux_h
    port map (
            O => \N__9416\,
            I => \N__9410\
        );

    \I__2168\ : Odrv12
    port map (
            O => \N__9413\,
            I => \DRA_c_2\
        );

    \I__2167\ : Odrv12
    port map (
            O => \N__9410\,
            I => \DRA_c_2\
        );

    \I__2166\ : InMux
    port map (
            O => \N__9405\,
            I => \N__9402\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9402\,
            I => \N__9399\
        );

    \I__2164\ : Span4Mux_h
    port map (
            O => \N__9399\,
            I => \N__9396\
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__9396\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__9393\,
            I => \N__9384\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9380\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__9391\,
            I => \N__9375\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9390\,
            I => \N__9372\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__9389\,
            I => \N__9366\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9388\,
            I => \N__9360\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9387\,
            I => \N__9360\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9384\,
            I => \N__9356\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9383\,
            I => \N__9353\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__9380\,
            I => \N__9350\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9379\,
            I => \N__9347\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9378\,
            I => \N__9341\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9341\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9372\,
            I => \N__9337\
        );

    \I__2148\ : InMux
    port map (
            O => \N__9371\,
            I => \N__9332\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9332\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9369\,
            I => \N__9329\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9366\,
            I => \N__9325\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9365\,
            I => \N__9322\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9360\,
            I => \N__9318\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9315\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9356\,
            I => \N__9311\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__9353\,
            I => \N__9308\
        );

    \I__2139\ : Span4Mux_v
    port map (
            O => \N__9350\,
            I => \N__9301\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9347\,
            I => \N__9301\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9346\,
            I => \N__9298\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9341\,
            I => \N__9295\
        );

    \I__2135\ : InMux
    port map (
            O => \N__9340\,
            I => \N__9290\
        );

    \I__2134\ : Span4Mux_v
    port map (
            O => \N__9337\,
            I => \N__9285\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__9332\,
            I => \N__9285\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9329\,
            I => \N__9282\
        );

    \I__2131\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9279\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__9325\,
            I => \N__9274\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__9322\,
            I => \N__9274\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9271\
        );

    \I__2127\ : Span4Mux_v
    port map (
            O => \N__9318\,
            I => \N__9266\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__9315\,
            I => \N__9266\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9263\
        );

    \I__2124\ : Span4Mux_h
    port map (
            O => \N__9311\,
            I => \N__9258\
        );

    \I__2123\ : Span4Mux_h
    port map (
            O => \N__9308\,
            I => \N__9258\
        );

    \I__2122\ : InMux
    port map (
            O => \N__9307\,
            I => \N__9253\
        );

    \I__2121\ : InMux
    port map (
            O => \N__9306\,
            I => \N__9253\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__9301\,
            I => \N__9246\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__9298\,
            I => \N__9246\
        );

    \I__2118\ : Span4Mux_v
    port map (
            O => \N__9295\,
            I => \N__9246\
        );

    \I__2117\ : InMux
    port map (
            O => \N__9294\,
            I => \N__9241\
        );

    \I__2116\ : InMux
    port map (
            O => \N__9293\,
            I => \N__9241\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9290\,
            I => \N__9236\
        );

    \I__2114\ : Span4Mux_h
    port map (
            O => \N__9285\,
            I => \N__9236\
        );

    \I__2113\ : Span12Mux_h
    port map (
            O => \N__9282\,
            I => \N__9227\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__9279\,
            I => \N__9227\
        );

    \I__2111\ : Span12Mux_h
    port map (
            O => \N__9274\,
            I => \N__9227\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9271\,
            I => \N__9227\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__9266\,
            I => \CPU_CYCLEm\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__9263\,
            I => \CPU_CYCLEm\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__9258\,
            I => \CPU_CYCLEm\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__9253\,
            I => \CPU_CYCLEm\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__9246\,
            I => \CPU_CYCLEm\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9241\,
            I => \CPU_CYCLEm\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__9236\,
            I => \CPU_CYCLEm\
        );

    \I__2102\ : Odrv12
    port map (
            O => \N__9227\,
            I => \CPU_CYCLEm\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9210\,
            I => \N__9207\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__9207\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__2099\ : InMux
    port map (
            O => \N__9204\,
            I => \N__9196\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9203\,
            I => \N__9191\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__9202\,
            I => \N__9188\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__9201\,
            I => \N__9185\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__9200\,
            I => \N__9182\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__9199\,
            I => \N__9177\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9196\,
            I => \N__9170\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9195\,
            I => \N__9167\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9194\,
            I => \N__9164\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9191\,
            I => \N__9161\
        );

    \I__2089\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9158\
        );

    \I__2088\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9155\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9150\
        );

    \I__2086\ : InMux
    port map (
            O => \N__9181\,
            I => \N__9144\
        );

    \I__2085\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9144\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9177\,
            I => \N__9137\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9176\,
            I => \N__9137\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9175\,
            I => \N__9137\
        );

    \I__2081\ : InMux
    port map (
            O => \N__9174\,
            I => \N__9130\
        );

    \I__2080\ : InMux
    port map (
            O => \N__9173\,
            I => \N__9130\
        );

    \I__2079\ : Span4Mux_h
    port map (
            O => \N__9170\,
            I => \N__9122\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__9167\,
            I => \N__9122\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__9164\,
            I => \N__9113\
        );

    \I__2076\ : Span4Mux_v
    port map (
            O => \N__9161\,
            I => \N__9113\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__9158\,
            I => \N__9113\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__9155\,
            I => \N__9113\
        );

    \I__2073\ : InMux
    port map (
            O => \N__9154\,
            I => \N__9108\
        );

    \I__2072\ : InMux
    port map (
            O => \N__9153\,
            I => \N__9108\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__9150\,
            I => \N__9105\
        );

    \I__2070\ : InMux
    port map (
            O => \N__9149\,
            I => \N__9101\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__9144\,
            I => \N__9098\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9137\,
            I => \N__9095\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9090\
        );

    \I__2066\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9090\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9130\,
            I => \N__9087\
        );

    \I__2064\ : InMux
    port map (
            O => \N__9129\,
            I => \N__9082\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9128\,
            I => \N__9082\
        );

    \I__2062\ : InMux
    port map (
            O => \N__9127\,
            I => \N__9079\
        );

    \I__2061\ : Span4Mux_h
    port map (
            O => \N__9122\,
            I => \N__9075\
        );

    \I__2060\ : Span4Mux_v
    port map (
            O => \N__9113\,
            I => \N__9072\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9108\,
            I => \N__9069\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__9105\,
            I => \N__9066\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9063\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__9101\,
            I => \N__9048\
        );

    \I__2055\ : Span4Mux_v
    port map (
            O => \N__9098\,
            I => \N__9048\
        );

    \I__2054\ : Span4Mux_v
    port map (
            O => \N__9095\,
            I => \N__9048\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9090\,
            I => \N__9048\
        );

    \I__2052\ : Span4Mux_h
    port map (
            O => \N__9087\,
            I => \N__9048\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__9082\,
            I => \N__9048\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9079\,
            I => \N__9048\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9078\,
            I => \N__9045\
        );

    \I__2048\ : Span4Mux_v
    port map (
            O => \N__9075\,
            I => \N__9042\
        );

    \I__2047\ : Span4Mux_h
    port map (
            O => \N__9072\,
            I => \N__9037\
        );

    \I__2046\ : Span4Mux_v
    port map (
            O => \N__9069\,
            I => \N__9037\
        );

    \I__2045\ : Sp12to4
    port map (
            O => \N__9066\,
            I => \N__9032\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__9063\,
            I => \N__9032\
        );

    \I__2043\ : Span4Mux_h
    port map (
            O => \N__9048\,
            I => \N__9029\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__9045\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2041\ : Odrv4
    port map (
            O => \N__9042\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__9037\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2039\ : Odrv12
    port map (
            O => \N__9032\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__9029\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9018\,
            I => \N__9015\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9015\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9012\,
            I => \N__9009\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9009\,
            I => \N__9006\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__9006\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9003\,
            I => \N__9000\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9000\,
            I => \N__8997\
        );

    \I__2030\ : Span4Mux_h
    port map (
            O => \N__8997\,
            I => \N__8994\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__8994\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2028\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8987\
        );

    \I__2027\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8984\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__8987\,
            I => \N__8981\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__8984\,
            I => \N__8978\
        );

    \I__2024\ : Span4Mux_h
    port map (
            O => \N__8981\,
            I => \N__8975\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__8978\,
            I => \N__8972\
        );

    \I__2022\ : Sp12to4
    port map (
            O => \N__8975\,
            I => \N__8969\
        );

    \I__2021\ : Sp12to4
    port map (
            O => \N__8972\,
            I => \N__8966\
        );

    \I__2020\ : Span12Mux_v
    port map (
            O => \N__8969\,
            I => \N__8963\
        );

    \I__2019\ : Span12Mux_h
    port map (
            O => \N__8966\,
            I => \N__8960\
        );

    \I__2018\ : Span12Mux_h
    port map (
            O => \N__8963\,
            I => \N__8955\
        );

    \I__2017\ : Span12Mux_v
    port map (
            O => \N__8960\,
            I => \N__8955\
        );

    \I__2016\ : Odrv12
    port map (
            O => \N__8955\,
            I => \DRA_c_0\
        );

    \I__2015\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8949\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__8949\,
            I => \N__8946\
        );

    \I__2013\ : Odrv12
    port map (
            O => \N__8946\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2012\ : InMux
    port map (
            O => \N__8943\,
            I => \N__8940\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__8940\,
            I => \N__8934\
        );

    \I__2010\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8929\
        );

    \I__2009\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8929\
        );

    \I__2008\ : InMux
    port map (
            O => \N__8937\,
            I => \N__8926\
        );

    \I__2007\ : Sp12to4
    port map (
            O => \N__8934\,
            I => \N__8919\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__8929\,
            I => \N__8919\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__8926\,
            I => \N__8919\
        );

    \I__2004\ : Span12Mux_v
    port map (
            O => \N__8919\,
            I => \N__8916\
        );

    \I__2003\ : Span12Mux_h
    port map (
            O => \N__8916\,
            I => \N__8913\
        );

    \I__2002\ : Odrv12
    port map (
            O => \N__8913\,
            I => \DRA_c_1\
        );

    \I__2001\ : InMux
    port map (
            O => \N__8910\,
            I => \N__8904\
        );

    \I__2000\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8904\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__8904\,
            I => \N__8901\
        );

    \I__1998\ : Span4Mux_v
    port map (
            O => \N__8901\,
            I => \N__8898\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__8898\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1996\ : IoInMux
    port map (
            O => \N__8895\,
            I => \N__8892\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__8892\,
            I => \N__8889\
        );

    \I__1994\ : Span4Mux_s0_v
    port map (
            O => \N__8889\,
            I => \N__8886\
        );

    \I__1993\ : Span4Mux_v
    port map (
            O => \N__8886\,
            I => \N__8883\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__8883\,
            I => \U712_BYTE_ENABLE_UUBE_i\
        );

    \I__1991\ : IoInMux
    port map (
            O => \N__8880\,
            I => \N__8877\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__8877\,
            I => \N__8874\
        );

    \I__1989\ : Span4Mux_s2_v
    port map (
            O => \N__8874\,
            I => \N__8871\
        );

    \I__1988\ : Span4Mux_v
    port map (
            O => \N__8871\,
            I => \N__8868\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__8868\,
            I => \N_215_i\
        );

    \I__1986\ : IoInMux
    port map (
            O => \N__8865\,
            I => \N__8862\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__8862\,
            I => \N__8859\
        );

    \I__1984\ : IoSpan4Mux
    port map (
            O => \N__8859\,
            I => \N__8856\
        );

    \I__1983\ : Span4Mux_s3_v
    port map (
            O => \N__8856\,
            I => \N__8853\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__8853\,
            I => \N_217_i\
        );

    \I__1981\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8844\
        );

    \I__1980\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8835\
        );

    \I__1979\ : InMux
    port map (
            O => \N__8848\,
            I => \N__8835\
        );

    \I__1978\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8835\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__8844\,
            I => \N__8832\
        );

    \I__1976\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8829\
        );

    \I__1975\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8826\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__8835\,
            I => \N__8823\
        );

    \I__1973\ : Span4Mux_h
    port map (
            O => \N__8832\,
            I => \N__8817\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__8829\,
            I => \N__8817\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__8826\,
            I => \N__8813\
        );

    \I__1970\ : Span4Mux_v
    port map (
            O => \N__8823\,
            I => \N__8810\
        );

    \I__1969\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8807\
        );

    \I__1968\ : Span4Mux_h
    port map (
            O => \N__8817\,
            I => \N__8804\
        );

    \I__1967\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8801\
        );

    \I__1966\ : Span12Mux_v
    port map (
            O => \N__8813\,
            I => \N__8798\
        );

    \I__1965\ : Sp12to4
    port map (
            O => \N__8810\,
            I => \N__8793\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__8807\,
            I => \N__8793\
        );

    \I__1963\ : Span4Mux_v
    port map (
            O => \N__8804\,
            I => \N__8790\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__8801\,
            I => \N__8787\
        );

    \I__1961\ : Span12Mux_h
    port map (
            O => \N__8798\,
            I => \N__8784\
        );

    \I__1960\ : Span12Mux_h
    port map (
            O => \N__8793\,
            I => \N__8777\
        );

    \I__1959\ : Sp12to4
    port map (
            O => \N__8790\,
            I => \N__8777\
        );

    \I__1958\ : Span12Mux_v
    port map (
            O => \N__8787\,
            I => \N__8777\
        );

    \I__1957\ : Odrv12
    port map (
            O => \N__8784\,
            I => \A_c_1\
        );

    \I__1956\ : Odrv12
    port map (
            O => \N__8777\,
            I => \A_c_1\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8772\,
            I => \N__8759\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8771\,
            I => \N__8759\
        );

    \I__1953\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8759\
        );

    \I__1952\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8756\
        );

    \I__1951\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8753\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8767\,
            I => \N__8750\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8747\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__8759\,
            I => \N__8741\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8756\,
            I => \N__8741\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__8753\,
            I => \N__8736\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__8750\,
            I => \N__8736\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__8747\,
            I => \N__8733\
        );

    \I__1943\ : InMux
    port map (
            O => \N__8746\,
            I => \N__8729\
        );

    \I__1942\ : Span4Mux_v
    port map (
            O => \N__8741\,
            I => \N__8725\
        );

    \I__1941\ : Span4Mux_v
    port map (
            O => \N__8736\,
            I => \N__8720\
        );

    \I__1940\ : Span4Mux_v
    port map (
            O => \N__8733\,
            I => \N__8720\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8732\,
            I => \N__8717\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__8729\,
            I => \N__8714\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8728\,
            I => \N__8711\
        );

    \I__1936\ : Sp12to4
    port map (
            O => \N__8725\,
            I => \N__8704\
        );

    \I__1935\ : Sp12to4
    port map (
            O => \N__8720\,
            I => \N__8704\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8717\,
            I => \N__8704\
        );

    \I__1933\ : Span4Mux_v
    port map (
            O => \N__8714\,
            I => \N__8701\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__8711\,
            I => \N__8698\
        );

    \I__1931\ : Span12Mux_h
    port map (
            O => \N__8704\,
            I => \N__8695\
        );

    \I__1930\ : Sp12to4
    port map (
            O => \N__8701\,
            I => \N__8690\
        );

    \I__1929\ : Span12Mux_v
    port map (
            O => \N__8698\,
            I => \N__8690\
        );

    \I__1928\ : Odrv12
    port map (
            O => \N__8695\,
            I => \A_c_0\
        );

    \I__1927\ : Odrv12
    port map (
            O => \N__8690\,
            I => \A_c_0\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__8685\,
            I => \N__8679\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__8684\,
            I => \N__8675\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__8683\,
            I => \N__8672\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__8682\,
            I => \N__8669\
        );

    \I__1922\ : InMux
    port map (
            O => \N__8679\,
            I => \N__8665\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8678\,
            I => \N__8662\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8655\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8655\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8655\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__8668\,
            I => \N__8652\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__8665\,
            I => \N__8649\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__8662\,
            I => \N__8646\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8655\,
            I => \N__8643\
        );

    \I__1913\ : InMux
    port map (
            O => \N__8652\,
            I => \N__8640\
        );

    \I__1912\ : Span4Mux_h
    port map (
            O => \N__8649\,
            I => \N__8634\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__8646\,
            I => \N__8634\
        );

    \I__1910\ : Span4Mux_h
    port map (
            O => \N__8643\,
            I => \N__8629\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__8640\,
            I => \N__8629\
        );

    \I__1908\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8626\
        );

    \I__1907\ : Span4Mux_v
    port map (
            O => \N__8634\,
            I => \N__8621\
        );

    \I__1906\ : Span4Mux_h
    port map (
            O => \N__8629\,
            I => \N__8621\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8626\,
            I => \N__8618\
        );

    \I__1904\ : Span4Mux_v
    port map (
            O => \N__8621\,
            I => \N__8615\
        );

    \I__1903\ : Span12Mux_v
    port map (
            O => \N__8618\,
            I => \N__8610\
        );

    \I__1902\ : Sp12to4
    port map (
            O => \N__8615\,
            I => \N__8610\
        );

    \I__1901\ : Odrv12
    port map (
            O => \N__8610\,
            I => \SIZ_c_0\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__8607\,
            I => \N__8602\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__8606\,
            I => \N__8599\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8605\,
            I => \N__8593\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8602\,
            I => \N__8590\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8599\,
            I => \N__8587\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8598\,
            I => \N__8580\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8597\,
            I => \N__8580\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8580\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__8593\,
            I => \N__8576\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__8590\,
            I => \N__8573\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__8587\,
            I => \N__8570\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8580\,
            I => \N__8567\
        );

    \I__1888\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8564\
        );

    \I__1887\ : Span4Mux_h
    port map (
            O => \N__8576\,
            I => \N__8557\
        );

    \I__1886\ : Span4Mux_v
    port map (
            O => \N__8573\,
            I => \N__8557\
        );

    \I__1885\ : Span4Mux_v
    port map (
            O => \N__8570\,
            I => \N__8557\
        );

    \I__1884\ : Span4Mux_h
    port map (
            O => \N__8567\,
            I => \N__8552\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__8564\,
            I => \N__8552\
        );

    \I__1882\ : Span4Mux_v
    port map (
            O => \N__8557\,
            I => \N__8547\
        );

    \I__1881\ : Span4Mux_h
    port map (
            O => \N__8552\,
            I => \N__8547\
        );

    \I__1880\ : Span4Mux_v
    port map (
            O => \N__8547\,
            I => \N__8544\
        );

    \I__1879\ : Span4Mux_h
    port map (
            O => \N__8544\,
            I => \N__8541\
        );

    \I__1878\ : Sp12to4
    port map (
            O => \N__8541\,
            I => \N__8538\
        );

    \I__1877\ : Odrv12
    port map (
            O => \N__8538\,
            I => \SIZ_c_1\
        );

    \I__1876\ : IoInMux
    port map (
            O => \N__8535\,
            I => \N__8532\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__8532\,
            I => \N__8529\
        );

    \I__1874\ : Span4Mux_s3_h
    port map (
            O => \N__8529\,
            I => \N__8526\
        );

    \I__1873\ : Span4Mux_v
    port map (
            O => \N__8526\,
            I => \N__8523\
        );

    \I__1872\ : Sp12to4
    port map (
            O => \N__8523\,
            I => \N__8520\
        );

    \I__1871\ : Span12Mux_h
    port map (
            O => \N__8520\,
            I => \N__8517\
        );

    \I__1870\ : Odrv12
    port map (
            O => \N__8517\,
            I => \WEn_c\
        );

    \I__1869\ : IoInMux
    port map (
            O => \N__8514\,
            I => \N__8511\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8511\,
            I => \N__8508\
        );

    \I__1867\ : Span4Mux_s0_v
    port map (
            O => \N__8508\,
            I => \N__8505\
        );

    \I__1866\ : Sp12to4
    port map (
            O => \N__8505\,
            I => \N__8502\
        );

    \I__1865\ : Span12Mux_h
    port map (
            O => \N__8502\,
            I => \N__8499\
        );

    \I__1864\ : Odrv12
    port map (
            O => \N__8499\,
            I => \CASn_c\
        );

    \I__1863\ : IoInMux
    port map (
            O => \N__8496\,
            I => \N__8493\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__8493\,
            I => \N__8490\
        );

    \I__1861\ : IoSpan4Mux
    port map (
            O => \N__8490\,
            I => \N__8487\
        );

    \I__1860\ : Span4Mux_s2_v
    port map (
            O => \N__8487\,
            I => \N__8484\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__8484\,
            I => \N__8481\
        );

    \I__1858\ : Span4Mux_v
    port map (
            O => \N__8481\,
            I => \N__8478\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__8478\,
            I => \CRCSn_c\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8472\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__8472\,
            I => \N__8469\
        );

    \I__1854\ : Odrv12
    port map (
            O => \N__8469\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8466\,
            I => \N__8461\
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__8465\,
            I => \N__8458\
        );

    \I__1851\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8454\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8461\,
            I => \N__8451\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8458\,
            I => \N__8448\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__8457\,
            I => \N__8445\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__8454\,
            I => \N__8442\
        );

    \I__1846\ : Span4Mux_h
    port map (
            O => \N__8451\,
            I => \N__8439\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8448\,
            I => \N__8436\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8445\,
            I => \N__8433\
        );

    \I__1843\ : Sp12to4
    port map (
            O => \N__8442\,
            I => \N__8429\
        );

    \I__1842\ : Span4Mux_v
    port map (
            O => \N__8439\,
            I => \N__8422\
        );

    \I__1841\ : Span4Mux_h
    port map (
            O => \N__8436\,
            I => \N__8422\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8433\,
            I => \N__8422\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8419\
        );

    \I__1838\ : Span12Mux_v
    port map (
            O => \N__8429\,
            I => \N__8416\
        );

    \I__1837\ : Span4Mux_h
    port map (
            O => \N__8422\,
            I => \N__8413\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__8419\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1835\ : Odrv12
    port map (
            O => \N__8416\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__8413\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8406\,
            I => \N__8400\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8405\,
            I => \N__8397\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8394\
        );

    \I__1830\ : InMux
    port map (
            O => \N__8403\,
            I => \N__8391\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__8400\,
            I => \N__8386\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__8397\,
            I => \N__8383\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8394\,
            I => \N__8380\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8391\,
            I => \N__8377\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8374\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__8389\,
            I => \N__8370\
        );

    \I__1823\ : Span4Mux_v
    port map (
            O => \N__8386\,
            I => \N__8367\
        );

    \I__1822\ : Span12Mux_h
    port map (
            O => \N__8383\,
            I => \N__8364\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__8380\,
            I => \N__8357\
        );

    \I__1820\ : Span4Mux_h
    port map (
            O => \N__8377\,
            I => \N__8357\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8374\,
            I => \N__8357\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8373\,
            I => \N__8354\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8351\
        );

    \I__1816\ : Span4Mux_h
    port map (
            O => \N__8367\,
            I => \N__8348\
        );

    \I__1815\ : Span12Mux_v
    port map (
            O => \N__8364\,
            I => \N__8345\
        );

    \I__1814\ : Span4Mux_h
    port map (
            O => \N__8357\,
            I => \N__8342\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8354\,
            I => \N__8339\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8351\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__8348\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1810\ : Odrv12
    port map (
            O => \N__8345\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__8342\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1808\ : Odrv12
    port map (
            O => \N__8339\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1807\ : IoInMux
    port map (
            O => \N__8328\,
            I => \N__8325\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8325\,
            I => \N__8322\
        );

    \I__1805\ : Span4Mux_s3_v
    port map (
            O => \N__8322\,
            I => \N__8319\
        );

    \I__1804\ : Sp12to4
    port map (
            O => \N__8319\,
            I => \N__8316\
        );

    \I__1803\ : Span12Mux_h
    port map (
            O => \N__8316\,
            I => \N__8313\
        );

    \I__1802\ : Odrv12
    port map (
            O => \N__8313\,
            I => \CMA_c_10\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8310\,
            I => \N__8307\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8307\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1799\ : IoInMux
    port map (
            O => \N__8304\,
            I => \N__8301\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8301\,
            I => \N__8298\
        );

    \I__1797\ : Span4Mux_s3_h
    port map (
            O => \N__8298\,
            I => \N__8295\
        );

    \I__1796\ : Span4Mux_v
    port map (
            O => \N__8295\,
            I => \N__8292\
        );

    \I__1795\ : Sp12to4
    port map (
            O => \N__8292\,
            I => \N__8289\
        );

    \I__1794\ : Span12Mux_h
    port map (
            O => \N__8289\,
            I => \N__8286\
        );

    \I__1793\ : Odrv12
    port map (
            O => \N__8286\,
            I => \CMA_c_4\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8283\,
            I => \N__8279\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8282\,
            I => \N__8276\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8279\,
            I => \N__8273\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8276\,
            I => \N__8270\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__8273\,
            I => \N__8263\
        );

    \I__1787\ : Span4Mux_h
    port map (
            O => \N__8270\,
            I => \N__8260\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8269\,
            I => \N__8255\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8268\,
            I => \N__8255\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8267\,
            I => \N__8250\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8266\,
            I => \N__8250\
        );

    \I__1782\ : Odrv4
    port map (
            O => \N__8263\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__8260\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8255\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8250\,
            I => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__8241\,
            I => \N__8238\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8238\,
            I => \N__8231\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__8237\,
            I => \N__8227\
        );

    \I__1775\ : CascadeMux
    port map (
            O => \N__8236\,
            I => \N__8223\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__8235\,
            I => \N__8220\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8234\,
            I => \N__8216\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8231\,
            I => \N__8213\
        );

    \I__1771\ : CascadeMux
    port map (
            O => \N__8230\,
            I => \N__8210\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8227\,
            I => \N__8207\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8226\,
            I => \N__8204\
        );

    \I__1768\ : InMux
    port map (
            O => \N__8223\,
            I => \N__8201\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8220\,
            I => \N__8198\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8219\,
            I => \N__8195\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8216\,
            I => \N__8192\
        );

    \I__1764\ : Span4Mux_v
    port map (
            O => \N__8213\,
            I => \N__8189\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8210\,
            I => \N__8186\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__8207\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8204\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__8201\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__8198\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__8195\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1757\ : Odrv12
    port map (
            O => \N__8192\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__8189\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__8186\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1754\ : IoInMux
    port map (
            O => \N__8169\,
            I => \N__8166\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__8166\,
            I => \N__8163\
        );

    \I__1752\ : Span4Mux_s2_h
    port map (
            O => \N__8163\,
            I => \N__8160\
        );

    \I__1751\ : Sp12to4
    port map (
            O => \N__8160\,
            I => \N__8157\
        );

    \I__1750\ : Span12Mux_s9_v
    port map (
            O => \N__8157\,
            I => \N__8154\
        );

    \I__1749\ : Span12Mux_h
    port map (
            O => \N__8154\,
            I => \N__8151\
        );

    \I__1748\ : Odrv12
    port map (
            O => \N__8151\,
            I => \CMA_c_6\
        );

    \I__1747\ : InMux
    port map (
            O => \N__8148\,
            I => \N__8145\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__8145\,
            I => \N__8140\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8144\,
            I => \N__8137\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8143\,
            I => \N__8134\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__8140\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__8137\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__8134\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8127\,
            I => \N__8124\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8124\,
            I => \N__8121\
        );

    \I__1738\ : Span4Mux_h
    port map (
            O => \N__8121\,
            I => \N__8118\
        );

    \I__1737\ : Sp12to4
    port map (
            O => \N__8118\,
            I => \N__8115\
        );

    \I__1736\ : Span12Mux_v
    port map (
            O => \N__8115\,
            I => \N__8112\
        );

    \I__1735\ : Span12Mux_h
    port map (
            O => \N__8112\,
            I => \N__8109\
        );

    \I__1734\ : Odrv12
    port map (
            O => \N__8109\,
            I => \A_c_19\
        );

    \I__1733\ : IoInMux
    port map (
            O => \N__8106\,
            I => \N__8103\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8103\,
            I => \N__8100\
        );

    \I__1731\ : IoSpan4Mux
    port map (
            O => \N__8100\,
            I => \N__8097\
        );

    \I__1730\ : Span4Mux_s0_h
    port map (
            O => \N__8097\,
            I => \N__8094\
        );

    \I__1729\ : Sp12to4
    port map (
            O => \N__8094\,
            I => \N__8091\
        );

    \I__1728\ : Span12Mux_h
    port map (
            O => \N__8091\,
            I => \N__8088\
        );

    \I__1727\ : Odrv12
    port map (
            O => \N__8088\,
            I => \CMA_c_9\
        );

    \I__1726\ : CEMux
    port map (
            O => \N__8085\,
            I => \N__8077\
        );

    \I__1725\ : CEMux
    port map (
            O => \N__8084\,
            I => \N__8074\
        );

    \I__1724\ : CEMux
    port map (
            O => \N__8083\,
            I => \N__8070\
        );

    \I__1723\ : CEMux
    port map (
            O => \N__8082\,
            I => \N__8067\
        );

    \I__1722\ : CEMux
    port map (
            O => \N__8081\,
            I => \N__8064\
        );

    \I__1721\ : CEMux
    port map (
            O => \N__8080\,
            I => \N__8061\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8077\,
            I => \N__8056\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8074\,
            I => \N__8056\
        );

    \I__1718\ : CEMux
    port map (
            O => \N__8073\,
            I => \N__8053\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8070\,
            I => \N__8050\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__8067\,
            I => \N__8047\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8064\,
            I => \N__8044\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8061\,
            I => \N__8041\
        );

    \I__1713\ : Span4Mux_v
    port map (
            O => \N__8056\,
            I => \N__8036\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__8053\,
            I => \N__8036\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__8050\,
            I => \N__8031\
        );

    \I__1710\ : Span4Mux_h
    port map (
            O => \N__8047\,
            I => \N__8031\
        );

    \I__1709\ : Span4Mux_h
    port map (
            O => \N__8044\,
            I => \N__8026\
        );

    \I__1708\ : Span4Mux_h
    port map (
            O => \N__8041\,
            I => \N__8026\
        );

    \I__1707\ : Span4Mux_v
    port map (
            O => \N__8036\,
            I => \N__8023\
        );

    \I__1706\ : Odrv4
    port map (
            O => \N__8031\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__8026\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__8023\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8016\,
            I => \N__8010\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8015\,
            I => \N__8010\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8010\,
            I => \N__8007\
        );

    \I__1700\ : Sp12to4
    port map (
            O => \N__8007\,
            I => \N__8004\
        );

    \I__1699\ : Span12Mux_v
    port map (
            O => \N__8004\,
            I => \N__8001\
        );

    \I__1698\ : Span12Mux_h
    port map (
            O => \N__8001\,
            I => \N__7998\
        );

    \I__1697\ : Odrv12
    port map (
            O => \N__7998\,
            I => \A_c_14\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__7995\,
            I => \U712_CHIP_RAM.CMA_5_0_8_cascade_\
        );

    \I__1695\ : InMux
    port map (
            O => \N__7992\,
            I => \N__7989\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__7989\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1693\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7983\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__7983\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i\
        );

    \I__1691\ : InMux
    port map (
            O => \N__7980\,
            I => \N__7977\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__7977\,
            I => \N__7974\
        );

    \I__1689\ : Span4Mux_v
    port map (
            O => \N__7974\,
            I => \N__7971\
        );

    \I__1688\ : Sp12to4
    port map (
            O => \N__7971\,
            I => \N__7968\
        );

    \I__1687\ : Span12Mux_h
    port map (
            O => \N__7968\,
            I => \N__7965\
        );

    \I__1686\ : Span12Mux_v
    port map (
            O => \N__7965\,
            I => \N__7962\
        );

    \I__1685\ : Odrv12
    port map (
            O => \N__7962\,
            I => \A_c_15\
        );

    \I__1684\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7956\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__7956\,
            I => \N__7953\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__7953\,
            I => \N__7950\
        );

    \I__1681\ : Sp12to4
    port map (
            O => \N__7950\,
            I => \N__7947\
        );

    \I__1680\ : Span12Mux_h
    port map (
            O => \N__7947\,
            I => \N__7944\
        );

    \I__1679\ : Odrv12
    port map (
            O => \N__7944\,
            I => \A_c_8\
        );

    \I__1678\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7938\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__7938\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1676\ : IoInMux
    port map (
            O => \N__7935\,
            I => \N__7932\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__7932\,
            I => \N__7929\
        );

    \I__1674\ : Span12Mux_s3_v
    port map (
            O => \N__7929\,
            I => \N__7926\
        );

    \I__1673\ : Span12Mux_v
    port map (
            O => \N__7926\,
            I => \N__7923\
        );

    \I__1672\ : Odrv12
    port map (
            O => \N__7923\,
            I => \CMA_c_0\
        );

    \I__1671\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7917\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__7917\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1669\ : IoInMux
    port map (
            O => \N__7914\,
            I => \N__7911\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__7911\,
            I => \N__7908\
        );

    \I__1667\ : IoSpan4Mux
    port map (
            O => \N__7908\,
            I => \N__7905\
        );

    \I__1666\ : Span4Mux_s2_h
    port map (
            O => \N__7905\,
            I => \N__7902\
        );

    \I__1665\ : Sp12to4
    port map (
            O => \N__7902\,
            I => \N__7899\
        );

    \I__1664\ : Span12Mux_h
    port map (
            O => \N__7899\,
            I => \N__7896\
        );

    \I__1663\ : Odrv12
    port map (
            O => \N__7896\,
            I => \CMA_c_7\
        );

    \I__1662\ : InMux
    port map (
            O => \N__7893\,
            I => \N__7890\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__7890\,
            I => \U712_CHIP_RAM.CLK_EN_6_0_a5_2\
        );

    \I__1660\ : InMux
    port map (
            O => \N__7887\,
            I => \N__7884\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__7884\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\
        );

    \I__1658\ : IoInMux
    port map (
            O => \N__7881\,
            I => \N__7878\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__7878\,
            I => \N__7875\
        );

    \I__1656\ : IoSpan4Mux
    port map (
            O => \N__7875\,
            I => \N__7872\
        );

    \I__1655\ : IoSpan4Mux
    port map (
            O => \N__7872\,
            I => \N__7869\
        );

    \I__1654\ : Span4Mux_s2_h
    port map (
            O => \N__7869\,
            I => \N__7866\
        );

    \I__1653\ : Sp12to4
    port map (
            O => \N__7866\,
            I => \N__7863\
        );

    \I__1652\ : Span12Mux_h
    port map (
            O => \N__7863\,
            I => \N__7859\
        );

    \I__1651\ : InMux
    port map (
            O => \N__7862\,
            I => \N__7856\
        );

    \I__1650\ : Odrv12
    port map (
            O => \N__7859\,
            I => \CLK_EN_c\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__7856\,
            I => \CLK_EN_c\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7851\,
            I => \N__7848\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__7848\,
            I => \N__7845\
        );

    \I__1646\ : Odrv4
    port map (
            O => \N__7845\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1645\ : InMux
    port map (
            O => \N__7842\,
            I => \N__7839\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__7839\,
            I => \N__7835\
        );

    \I__1643\ : InMux
    port map (
            O => \N__7838\,
            I => \N__7832\
        );

    \I__1642\ : Span4Mux_v
    port map (
            O => \N__7835\,
            I => \N__7829\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7832\,
            I => \N__7826\
        );

    \I__1640\ : Span4Mux_h
    port map (
            O => \N__7829\,
            I => \N__7823\
        );

    \I__1639\ : Span4Mux_v
    port map (
            O => \N__7826\,
            I => \N__7820\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__7823\,
            I => \N__7816\
        );

    \I__1637\ : Span4Mux_h
    port map (
            O => \N__7820\,
            I => \N__7813\
        );

    \I__1636\ : InMux
    port map (
            O => \N__7819\,
            I => \N__7810\
        );

    \I__1635\ : Odrv4
    port map (
            O => \N__7816\,
            I => \DS_ENm\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__7813\,
            I => \DS_ENm\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7810\,
            I => \DS_ENm\
        );

    \I__1632\ : IoInMux
    port map (
            O => \N__7803\,
            I => \N__7800\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__7800\,
            I => \N__7797\
        );

    \I__1630\ : Span4Mux_s2_v
    port map (
            O => \N__7797\,
            I => \N__7794\
        );

    \I__1629\ : Span4Mux_h
    port map (
            O => \N__7794\,
            I => \N__7791\
        );

    \I__1628\ : Span4Mux_h
    port map (
            O => \N__7791\,
            I => \N__7788\
        );

    \I__1627\ : Span4Mux_v
    port map (
            O => \N__7788\,
            I => \N__7785\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__7785\,
            I => \U712_BYTE_ENABLE_un1_UDSn_i\
        );

    \I__1625\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7774\
        );

    \I__1624\ : InMux
    port map (
            O => \N__7781\,
            I => \N__7771\
        );

    \I__1623\ : InMux
    port map (
            O => \N__7780\,
            I => \N__7768\
        );

    \I__1622\ : InMux
    port map (
            O => \N__7779\,
            I => \N__7765\
        );

    \I__1621\ : InMux
    port map (
            O => \N__7778\,
            I => \N__7762\
        );

    \I__1620\ : InMux
    port map (
            O => \N__7777\,
            I => \N__7759\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7774\,
            I => \N__7736\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__7771\,
            I => \N__7736\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__7768\,
            I => \N__7729\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__7765\,
            I => \N__7729\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__7762\,
            I => \N__7729\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7759\,
            I => \N__7726\
        );

    \I__1613\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7721\
        );

    \I__1612\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7721\
        );

    \I__1611\ : InMux
    port map (
            O => \N__7756\,
            I => \N__7718\
        );

    \I__1610\ : InMux
    port map (
            O => \N__7755\,
            I => \N__7715\
        );

    \I__1609\ : InMux
    port map (
            O => \N__7754\,
            I => \N__7712\
        );

    \I__1608\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7709\
        );

    \I__1607\ : InMux
    port map (
            O => \N__7752\,
            I => \N__7706\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7751\,
            I => \N__7699\
        );

    \I__1605\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7699\
        );

    \I__1604\ : InMux
    port map (
            O => \N__7749\,
            I => \N__7699\
        );

    \I__1603\ : InMux
    port map (
            O => \N__7748\,
            I => \N__7696\
        );

    \I__1602\ : InMux
    port map (
            O => \N__7747\,
            I => \N__7693\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7684\
        );

    \I__1600\ : InMux
    port map (
            O => \N__7745\,
            I => \N__7684\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7744\,
            I => \N__7684\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7743\,
            I => \N__7684\
        );

    \I__1597\ : InMux
    port map (
            O => \N__7742\,
            I => \N__7681\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7678\
        );

    \I__1595\ : Span4Mux_v
    port map (
            O => \N__7736\,
            I => \N__7673\
        );

    \I__1594\ : Span4Mux_v
    port map (
            O => \N__7729\,
            I => \N__7673\
        );

    \I__1593\ : Span4Mux_v
    port map (
            O => \N__7726\,
            I => \N__7660\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__7721\,
            I => \N__7660\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__7718\,
            I => \N__7660\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__7715\,
            I => \N__7660\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7712\,
            I => \N__7660\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__7709\,
            I => \N__7660\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__7706\,
            I => \N__7657\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__7699\,
            I => \N__7654\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7696\,
            I => \N__7647\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7693\,
            I => \N__7647\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__7684\,
            I => \N__7647\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7681\,
            I => \N__7641\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7678\,
            I => \N__7638\
        );

    \I__1580\ : Span4Mux_h
    port map (
            O => \N__7673\,
            I => \N__7631\
        );

    \I__1579\ : Span4Mux_v
    port map (
            O => \N__7660\,
            I => \N__7631\
        );

    \I__1578\ : Span4Mux_v
    port map (
            O => \N__7657\,
            I => \N__7631\
        );

    \I__1577\ : Span4Mux_v
    port map (
            O => \N__7654\,
            I => \N__7626\
        );

    \I__1576\ : Span4Mux_v
    port map (
            O => \N__7647\,
            I => \N__7626\
        );

    \I__1575\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7623\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7645\,
            I => \N__7620\
        );

    \I__1573\ : InMux
    port map (
            O => \N__7644\,
            I => \N__7617\
        );

    \I__1572\ : Span12Mux_v
    port map (
            O => \N__7641\,
            I => \N__7610\
        );

    \I__1571\ : Span12Mux_h
    port map (
            O => \N__7638\,
            I => \N__7610\
        );

    \I__1570\ : Sp12to4
    port map (
            O => \N__7631\,
            I => \N__7610\
        );

    \I__1569\ : Sp12to4
    port map (
            O => \N__7626\,
            I => \N__7601\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7623\,
            I => \N__7601\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__7620\,
            I => \N__7601\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7617\,
            I => \N__7601\
        );

    \I__1565\ : Span12Mux_h
    port map (
            O => \N__7610\,
            I => \N__7598\
        );

    \I__1564\ : Span12Mux_h
    port map (
            O => \N__7601\,
            I => \N__7595\
        );

    \I__1563\ : Odrv12
    port map (
            O => \N__7598\,
            I => \RESETn_c\
        );

    \I__1562\ : Odrv12
    port map (
            O => \N__7595\,
            I => \RESETn_c\
        );

    \I__1561\ : IoInMux
    port map (
            O => \N__7590\,
            I => \N__7587\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__7587\,
            I => \N__7584\
        );

    \I__1559\ : Span12Mux_s2_v
    port map (
            O => \N__7584\,
            I => \N__7581\
        );

    \I__1558\ : Odrv12
    port map (
            O => \N__7581\,
            I => \RESETn_c_i\
        );

    \I__1557\ : IoInMux
    port map (
            O => \N__7578\,
            I => \N__7575\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7575\,
            I => \N__7572\
        );

    \I__1555\ : Span12Mux_s11_v
    port map (
            O => \N__7572\,
            I => \N__7569\
        );

    \I__1554\ : Span12Mux_h
    port map (
            O => \N__7569\,
            I => \N__7566\
        );

    \I__1553\ : Odrv12
    port map (
            O => \N__7566\,
            I => \N_163\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7563\,
            I => \N__7560\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7560\,
            I => \N__7557\
        );

    \I__1550\ : Span4Mux_v
    port map (
            O => \N__7557\,
            I => \N__7554\
        );

    \I__1549\ : Span4Mux_v
    port map (
            O => \N__7554\,
            I => \N__7551\
        );

    \I__1548\ : Sp12to4
    port map (
            O => \N__7551\,
            I => \N__7548\
        );

    \I__1547\ : Span12Mux_h
    port map (
            O => \N__7548\,
            I => \N__7545\
        );

    \I__1546\ : Odrv12
    port map (
            O => \N__7545\,
            I => \A_c_17\
        );

    \I__1545\ : IoInMux
    port map (
            O => \N__7542\,
            I => \N__7539\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7539\,
            I => \N__7536\
        );

    \I__1543\ : Span12Mux_s3_h
    port map (
            O => \N__7536\,
            I => \N__7533\
        );

    \I__1542\ : Span12Mux_h
    port map (
            O => \N__7533\,
            I => \N__7530\
        );

    \I__1541\ : Odrv12
    port map (
            O => \N__7530\,
            I => \CMA_c_8\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__7527\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7521\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7521\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7518\,
            I => \N__7515\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7515\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7509\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7509\,
            I => \N__7506\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__7506\,
            I => \U712_CHIP_RAM.N_146\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__7503\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5_cascade_\
        );

    \I__1531\ : IoInMux
    port map (
            O => \N__7500\,
            I => \N__7497\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7497\,
            I => \N__7494\
        );

    \I__1529\ : Span4Mux_s3_h
    port map (
            O => \N__7494\,
            I => \N__7491\
        );

    \I__1528\ : Sp12to4
    port map (
            O => \N__7491\,
            I => \N__7488\
        );

    \I__1527\ : Span12Mux_s8_v
    port map (
            O => \N__7488\,
            I => \N__7485\
        );

    \I__1526\ : Span12Mux_h
    port map (
            O => \N__7485\,
            I => \N__7482\
        );

    \I__1525\ : Odrv12
    port map (
            O => \N__7482\,
            I => \CMA_c_5\
        );

    \I__1524\ : InMux
    port map (
            O => \N__7479\,
            I => \N__7476\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7476\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1522\ : CascadeMux
    port map (
            O => \N__7473\,
            I => \N__7468\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7465\
        );

    \I__1520\ : InMux
    port map (
            O => \N__7471\,
            I => \N__7462\
        );

    \I__1519\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7459\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7465\,
            I => \N__7454\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__7462\,
            I => \N__7454\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__7459\,
            I => \REG_TACK\
        );

    \I__1515\ : Odrv12
    port map (
            O => \N__7454\,
            I => \REG_TACK\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7449\,
            I => \N__7445\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7448\,
            I => \N__7441\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__7445\,
            I => \N__7438\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7444\,
            I => \N__7435\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7441\,
            I => \N__7432\
        );

    \I__1509\ : Span4Mux_h
    port map (
            O => \N__7438\,
            I => \N__7427\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7435\,
            I => \N__7427\
        );

    \I__1507\ : Odrv12
    port map (
            O => \N__7432\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1506\ : Odrv4
    port map (
            O => \N__7427\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7422\,
            I => \N__7416\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7421\,
            I => \N__7413\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7420\,
            I => \N__7409\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7406\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7416\,
            I => \N__7399\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7413\,
            I => \N__7399\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7412\,
            I => \N__7396\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7409\,
            I => \N__7393\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7406\,
            I => \N__7389\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7405\,
            I => \N__7384\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7404\,
            I => \N__7384\
        );

    \I__1494\ : Span4Mux_v
    port map (
            O => \N__7399\,
            I => \N__7379\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__7396\,
            I => \N__7379\
        );

    \I__1492\ : Span4Mux_h
    port map (
            O => \N__7393\,
            I => \N__7376\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7392\,
            I => \N__7373\
        );

    \I__1490\ : Odrv12
    port map (
            O => \N__7389\,
            I => \WRITE_CYCLEm\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__7384\,
            I => \WRITE_CYCLEm\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__7379\,
            I => \WRITE_CYCLEm\
        );

    \I__1487\ : Odrv4
    port map (
            O => \N__7376\,
            I => \WRITE_CYCLEm\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7373\,
            I => \WRITE_CYCLEm\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__7362\,
            I => \N__7359\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7359\,
            I => \N__7356\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7356\,
            I => \N__7353\
        );

    \I__1482\ : Span4Mux_h
    port map (
            O => \N__7353\,
            I => \N__7349\
        );

    \I__1481\ : InMux
    port map (
            O => \N__7352\,
            I => \N__7346\
        );

    \I__1480\ : Odrv4
    port map (
            O => \N__7349\,
            I => \CPU_TACKm\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7346\,
            I => \CPU_TACKm\
        );

    \I__1478\ : CEMux
    port map (
            O => \N__7341\,
            I => \N__7338\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__7338\,
            I => \N__7335\
        );

    \I__1476\ : Odrv4
    port map (
            O => \N__7335\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\
        );

    \I__1475\ : IoInMux
    port map (
            O => \N__7332\,
            I => \N__7329\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7329\,
            I => \N__7326\
        );

    \I__1473\ : IoSpan4Mux
    port map (
            O => \N__7326\,
            I => \N__7323\
        );

    \I__1472\ : Span4Mux_s3_h
    port map (
            O => \N__7323\,
            I => \N__7320\
        );

    \I__1471\ : Sp12to4
    port map (
            O => \N__7320\,
            I => \N__7317\
        );

    \I__1470\ : Span12Mux_s8_h
    port map (
            O => \N__7317\,
            I => \N__7314\
        );

    \I__1469\ : Span12Mux_v
    port map (
            O => \N__7314\,
            I => \N__7311\
        );

    \I__1468\ : Odrv12
    port map (
            O => \N__7311\,
            I => \N_118_i\
        );

    \I__1467\ : IoInMux
    port map (
            O => \N__7308\,
            I => \N__7305\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7305\,
            I => \N__7302\
        );

    \I__1465\ : Span4Mux_s0_h
    port map (
            O => \N__7302\,
            I => \N__7299\
        );

    \I__1464\ : Sp12to4
    port map (
            O => \N__7299\,
            I => \N__7296\
        );

    \I__1463\ : Span12Mux_s6_v
    port map (
            O => \N__7296\,
            I => \N__7293\
        );

    \I__1462\ : Span12Mux_h
    port map (
            O => \N__7293\,
            I => \N__7290\
        );

    \I__1461\ : Span12Mux_v
    port map (
            O => \N__7290\,
            I => \N__7287\
        );

    \I__1460\ : Odrv12
    port map (
            O => \N__7287\,
            I => \N_119_i\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7284\,
            I => \N__7281\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7281\,
            I => \N__7277\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7274\
        );

    \I__1456\ : Span4Mux_h
    port map (
            O => \N__7277\,
            I => \N__7268\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7274\,
            I => \N__7265\
        );

    \I__1454\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7262\
        );

    \I__1453\ : InMux
    port map (
            O => \N__7272\,
            I => \N__7257\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7257\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__7268\,
            I => \U712_CHIP_RAM.N_323\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__7265\,
            I => \U712_CHIP_RAM.N_323\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7262\,
            I => \U712_CHIP_RAM.N_323\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7257\,
            I => \U712_CHIP_RAM.N_323\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7248\,
            I => \N__7242\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__7247\,
            I => \N__7238\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7246\,
            I => \N__7230\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7230\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7242\,
            I => \N__7226\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7241\,
            I => \N__7218\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7218\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__7237\,
            I => \N__7213\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7236\,
            I => \N__7210\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7207\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7230\,
            I => \N__7204\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7229\,
            I => \N__7201\
        );

    \I__1435\ : Span4Mux_h
    port map (
            O => \N__7226\,
            I => \N__7198\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7225\,
            I => \N__7191\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7224\,
            I => \N__7191\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7223\,
            I => \N__7191\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__7218\,
            I => \N__7188\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7217\,
            I => \N__7183\
        );

    \I__1429\ : InMux
    port map (
            O => \N__7216\,
            I => \N__7183\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7180\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__7210\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__7207\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1425\ : Odrv4
    port map (
            O => \N__7204\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7201\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1423\ : Odrv4
    port map (
            O => \N__7198\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7191\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1421\ : Odrv4
    port map (
            O => \N__7188\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7183\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__7180\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__7161\,
            I => \N__7156\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7160\,
            I => \N__7152\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7149\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7142\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__7155\,
            I => \N__7138\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7152\,
            I => \N__7135\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7149\,
            I => \N__7132\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7148\,
            I => \N__7127\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7147\,
            I => \N__7127\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__7146\,
            I => \N__7124\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7118\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7142\,
            I => \N__7115\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7141\,
            I => \N__7112\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7138\,
            I => \N__7109\
        );

    \I__1404\ : Span4Mux_v
    port map (
            O => \N__7135\,
            I => \N__7102\
        );

    \I__1403\ : Span4Mux_v
    port map (
            O => \N__7132\,
            I => \N__7102\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__7127\,
            I => \N__7102\
        );

    \I__1401\ : InMux
    port map (
            O => \N__7124\,
            I => \N__7097\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7097\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7122\,
            I => \N__7094\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7121\,
            I => \N__7091\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__7118\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1396\ : Odrv4
    port map (
            O => \N__7115\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7112\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7109\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__7102\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7097\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7094\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7091\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1389\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7071\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__7071\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_a5_0_1_0\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__7068\,
            I => \N__7065\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7065\,
            I => \N__7062\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7062\,
            I => \U712_CHIP_RAM.N_287\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7059\,
            I => \N__7053\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7058\,
            I => \N__7050\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7057\,
            I => \N__7047\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7056\,
            I => \N__7044\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7053\,
            I => \N__7041\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__7050\,
            I => \N__7038\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__7047\,
            I => \N__7033\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7044\,
            I => \N__7030\
        );

    \I__1376\ : Span4Mux_v
    port map (
            O => \N__7041\,
            I => \N__7024\
        );

    \I__1375\ : Span4Mux_v
    port map (
            O => \N__7038\,
            I => \N__7024\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7037\,
            I => \N__7019\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7036\,
            I => \N__7019\
        );

    \I__1372\ : Span4Mux_v
    port map (
            O => \N__7033\,
            I => \N__7014\
        );

    \I__1371\ : Span4Mux_v
    port map (
            O => \N__7030\,
            I => \N__7014\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7029\,
            I => \N__7011\
        );

    \I__1369\ : Odrv4
    port map (
            O => \N__7024\,
            I => \DMA_CYCLEm\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7019\,
            I => \DMA_CYCLEm\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__7014\,
            I => \DMA_CYCLEm\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7011\,
            I => \DMA_CYCLEm\
        );

    \I__1365\ : IoInMux
    port map (
            O => \N__7002\,
            I => \N__6999\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__6999\,
            I => \N__6995\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6998\,
            I => \N__6992\
        );

    \I__1362\ : Span12Mux_s4_v
    port map (
            O => \N__6995\,
            I => \N__6989\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6992\,
            I => \N__6986\
        );

    \I__1360\ : Span12Mux_v
    port map (
            O => \N__6989\,
            I => \N__6981\
        );

    \I__1359\ : Span4Mux_v
    port map (
            O => \N__6986\,
            I => \N__6978\
        );

    \I__1358\ : InMux
    port map (
            O => \N__6985\,
            I => \N__6975\
        );

    \I__1357\ : InMux
    port map (
            O => \N__6984\,
            I => \N__6972\
        );

    \I__1356\ : Odrv12
    port map (
            O => \N__6981\,
            I => \DBENn_c\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__6978\,
            I => \DBENn_c\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6975\,
            I => \DBENn_c\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__6972\,
            I => \DBENn_c\
        );

    \I__1352\ : InMux
    port map (
            O => \N__6963\,
            I => \N__6957\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6962\,
            I => \N__6957\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6957\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_a5_0Z0Z_0\
        );

    \I__1349\ : CascadeMux
    port map (
            O => \N__6954\,
            I => \N__6951\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6951\,
            I => \N__6948\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__6948\,
            I => \N__6945\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__6945\,
            I => \U712_BYTE_ENABLE.UUBE\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6939\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__6939\,
            I => \N__6936\
        );

    \I__1343\ : Odrv4
    port map (
            O => \N__6936\,
            I => \U712_BYTE_ENABLE.N_216\
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__6933\,
            I => \N__6930\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6930\,
            I => \N__6927\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__6927\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6921\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6921\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6918\,
            I => \N__6915\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__6915\,
            I => \N__6912\
        );

    \I__1335\ : Span12Mux_h
    port map (
            O => \N__6912\,
            I => \N__6909\
        );

    \I__1334\ : Odrv12
    port map (
            O => \N__6909\,
            I => \A_c_9\
        );

    \I__1333\ : InMux
    port map (
            O => \N__6906\,
            I => \N__6903\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6903\,
            I => \N__6900\
        );

    \I__1331\ : Span12Mux_v
    port map (
            O => \N__6900\,
            I => \N__6897\
        );

    \I__1330\ : Span12Mux_h
    port map (
            O => \N__6897\,
            I => \N__6894\
        );

    \I__1329\ : Odrv12
    port map (
            O => \N__6894\,
            I => \A_c_2\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__6891\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\
        );

    \I__1327\ : InMux
    port map (
            O => \N__6888\,
            I => \N__6885\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__6885\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1325\ : InMux
    port map (
            O => \N__6882\,
            I => \N__6879\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6879\,
            I => \N__6876\
        );

    \I__1323\ : Span12Mux_v
    port map (
            O => \N__6876\,
            I => \N__6873\
        );

    \I__1322\ : Span12Mux_h
    port map (
            O => \N__6873\,
            I => \N__6870\
        );

    \I__1321\ : Odrv12
    port map (
            O => \N__6870\,
            I => \A_c_7\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6867\,
            I => \N__6862\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__6866\,
            I => \N__6859\
        );

    \I__1318\ : InMux
    port map (
            O => \N__6865\,
            I => \N__6856\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__6862\,
            I => \N__6853\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6859\,
            I => \N__6850\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__6856\,
            I => \N__6846\
        );

    \I__1314\ : Span4Mux_h
    port map (
            O => \N__6853\,
            I => \N__6841\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6850\,
            I => \N__6841\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6838\
        );

    \I__1311\ : Span4Mux_v
    port map (
            O => \N__6846\,
            I => \N__6833\
        );

    \I__1310\ : Span4Mux_h
    port map (
            O => \N__6841\,
            I => \N__6833\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6838\,
            I => \N__6830\
        );

    \I__1308\ : Span4Mux_v
    port map (
            O => \N__6833\,
            I => \N__6827\
        );

    \I__1307\ : Span12Mux_h
    port map (
            O => \N__6830\,
            I => \N__6824\
        );

    \I__1306\ : Span4Mux_v
    port map (
            O => \N__6827\,
            I => \N__6821\
        );

    \I__1305\ : Span12Mux_v
    port map (
            O => \N__6824\,
            I => \N__6818\
        );

    \I__1304\ : Span4Mux_v
    port map (
            O => \N__6821\,
            I => \N__6815\
        );

    \I__1303\ : Odrv12
    port map (
            O => \N__6818\,
            I => \CLK40_PLL_i\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__6815\,
            I => \CLK40_PLL_i\
        );

    \I__1301\ : IoInMux
    port map (
            O => \N__6810\,
            I => \N__6807\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6807\,
            I => \N__6802\
        );

    \I__1299\ : IoInMux
    port map (
            O => \N__6806\,
            I => \N__6799\
        );

    \I__1298\ : IoInMux
    port map (
            O => \N__6805\,
            I => \N__6796\
        );

    \I__1297\ : Span4Mux_s1_v
    port map (
            O => \N__6802\,
            I => \N__6793\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__6799\,
            I => \N__6790\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__6796\,
            I => \N__6787\
        );

    \I__1294\ : Span4Mux_h
    port map (
            O => \N__6793\,
            I => \N__6784\
        );

    \I__1293\ : Span4Mux_s1_v
    port map (
            O => \N__6790\,
            I => \N__6781\
        );

    \I__1292\ : Span4Mux_s3_h
    port map (
            O => \N__6787\,
            I => \N__6778\
        );

    \I__1291\ : Sp12to4
    port map (
            O => \N__6784\,
            I => \N__6773\
        );

    \I__1290\ : Sp12to4
    port map (
            O => \N__6781\,
            I => \N__6773\
        );

    \I__1289\ : Span4Mux_h
    port map (
            O => \N__6778\,
            I => \N__6770\
        );

    \I__1288\ : Span12Mux_h
    port map (
            O => \N__6773\,
            I => \N__6767\
        );

    \I__1287\ : Span4Mux_h
    port map (
            O => \N__6770\,
            I => \N__6764\
        );

    \I__1286\ : Span12Mux_v
    port map (
            O => \N__6767\,
            I => \N__6761\
        );

    \I__1285\ : Span4Mux_h
    port map (
            O => \N__6764\,
            I => \N__6758\
        );

    \I__1284\ : Odrv12
    port map (
            O => \N__6761\,
            I => \CLK40_PLL_i_i\
        );

    \I__1283\ : Odrv4
    port map (
            O => \N__6758\,
            I => \CLK40_PLL_i_i\
        );

    \I__1282\ : InMux
    port map (
            O => \N__6753\,
            I => \N__6750\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6750\,
            I => \N__6744\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6749\,
            I => \N__6741\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6734\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6731\
        );

    \I__1277\ : Span4Mux_h
    port map (
            O => \N__6744\,
            I => \N__6726\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__6741\,
            I => \N__6726\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6740\,
            I => \N__6723\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6739\,
            I => \N__6720\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6738\,
            I => \N__6715\
        );

    \I__1272\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6715\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__6734\,
            I => \U712_CHIP_RAM.N_327\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__6731\,
            I => \U712_CHIP_RAM.N_327\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__6726\,
            I => \U712_CHIP_RAM.N_327\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6723\,
            I => \U712_CHIP_RAM.N_327\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__6720\,
            I => \U712_CHIP_RAM.N_327\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__6715\,
            I => \U712_CHIP_RAM.N_327\
        );

    \I__1265\ : InMux
    port map (
            O => \N__6702\,
            I => \N__6697\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6701\,
            I => \N__6694\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6700\,
            I => \N__6691\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__6697\,
            I => \U712_CHIP_RAM.N_339\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6694\,
            I => \U712_CHIP_RAM.N_339\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6691\,
            I => \U712_CHIP_RAM.N_339\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__6684\,
            I => \N__6680\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__6683\,
            I => \N__6677\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6669\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6677\,
            I => \N__6669\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6676\,
            I => \N__6664\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6664\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__6674\,
            I => \N__6658\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6669\,
            I => \N__6651\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__6664\,
            I => \N__6651\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6663\,
            I => \N__6646\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__6662\,
            I => \N__6642\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6661\,
            I => \N__6636\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6658\,
            I => \N__6636\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6657\,
            I => \N__6630\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6656\,
            I => \N__6627\
        );

    \I__1244\ : Span4Mux_v
    port map (
            O => \N__6651\,
            I => \N__6624\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6650\,
            I => \N__6619\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6649\,
            I => \N__6619\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6646\,
            I => \N__6616\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6645\,
            I => \N__6613\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6642\,
            I => \N__6608\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6641\,
            I => \N__6608\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6636\,
            I => \N__6605\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6600\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6600\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6633\,
            I => \N__6597\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6630\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6627\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1231\ : Odrv4
    port map (
            O => \N__6624\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__6619\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__6616\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__6613\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6608\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1226\ : Odrv12
    port map (
            O => \N__6605\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6600\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6597\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__6576\,
            I => \N__6568\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__6575\,
            I => \N__6565\
        );

    \I__1221\ : CascadeMux
    port map (
            O => \N__6574\,
            I => \N__6558\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__6573\,
            I => \N__6555\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6551\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6542\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6568\,
            I => \N__6542\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6565\,
            I => \N__6542\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6564\,
            I => \N__6539\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6535\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6530\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6561\,
            I => \N__6530\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6558\,
            I => \N__6527\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6524\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6521\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6551\,
            I => \N__6518\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6513\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6513\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6542\,
            I => \N__6510\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6539\,
            I => \N__6507\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6538\,
            I => \N__6504\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6535\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6530\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6527\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6524\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6521\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1197\ : Odrv4
    port map (
            O => \N__6518\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6513\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__6510\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1194\ : Odrv4
    port map (
            O => \N__6507\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6504\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__6483\,
            I => \N__6480\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6477\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__6477\,
            I => \U712_CHIP_RAM.un3_DMA_CYCLE_START\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6471\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6471\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6462\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6467\,
            I => \N__6462\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6462\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1184\ : IoInMux
    port map (
            O => \N__6459\,
            I => \N__6456\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6456\,
            I => \N__6453\
        );

    \I__1182\ : IoSpan4Mux
    port map (
            O => \N__6453\,
            I => \N__6450\
        );

    \I__1181\ : Span4Mux_s3_v
    port map (
            O => \N__6450\,
            I => \N__6447\
        );

    \I__1180\ : Span4Mux_v
    port map (
            O => \N__6447\,
            I => \N__6444\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__6444\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6441\,
            I => \N__6438\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6438\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1176\ : IoInMux
    port map (
            O => \N__6435\,
            I => \N__6432\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6432\,
            I => \N__6429\
        );

    \I__1174\ : Span12Mux_s5_v
    port map (
            O => \N__6429\,
            I => \N__6426\
        );

    \I__1173\ : Odrv12
    port map (
            O => \N__6426\,
            I => \CMA_c_1\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6423\,
            I => \N__6420\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6420\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1170\ : IoInMux
    port map (
            O => \N__6417\,
            I => \N__6414\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6414\,
            I => \N__6411\
        );

    \I__1168\ : IoSpan4Mux
    port map (
            O => \N__6411\,
            I => \N__6408\
        );

    \I__1167\ : Span4Mux_s3_v
    port map (
            O => \N__6408\,
            I => \N__6405\
        );

    \I__1166\ : Sp12to4
    port map (
            O => \N__6405\,
            I => \N__6402\
        );

    \I__1165\ : Odrv12
    port map (
            O => \N__6402\,
            I => \CMA_c_2\
        );

    \I__1164\ : IoInMux
    port map (
            O => \N__6399\,
            I => \N__6396\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6396\,
            I => \N__6393\
        );

    \I__1162\ : Span12Mux_s6_h
    port map (
            O => \N__6393\,
            I => \N__6390\
        );

    \I__1161\ : Span12Mux_v
    port map (
            O => \N__6390\,
            I => \N__6387\
        );

    \I__1160\ : Odrv12
    port map (
            O => \N__6387\,
            I => \CMA_c_3\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6384\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__1158\ : CEMux
    port map (
            O => \N__6381\,
            I => \N__6378\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6378\,
            I => \N__6375\
        );

    \I__1156\ : Span4Mux_v
    port map (
            O => \N__6375\,
            I => \N__6371\
        );

    \I__1155\ : CEMux
    port map (
            O => \N__6374\,
            I => \N__6368\
        );

    \I__1154\ : Span4Mux_h
    port map (
            O => \N__6371\,
            I => \N__6365\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6368\,
            I => \N__6362\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__6365\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__6362\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6354\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6354\,
            I => \N__6351\
        );

    \I__1148\ : Span4Mux_v
    port map (
            O => \N__6351\,
            I => \N__6348\
        );

    \I__1147\ : Sp12to4
    port map (
            O => \N__6348\,
            I => \N__6345\
        );

    \I__1146\ : Span12Mux_h
    port map (
            O => \N__6345\,
            I => \N__6342\
        );

    \I__1145\ : Odrv12
    port map (
            O => \N__6342\,
            I => \A_c_20\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__6339\,
            I => \U712_CHIP_RAM.N_289_cascade_\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6333\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__6333\,
            I => \N__6330\
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__6330\,
            I => \U712_CHIP_RAM.N_288\
        );

    \I__1140\ : IoInMux
    port map (
            O => \N__6327\,
            I => \N__6324\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6324\,
            I => \N__6321\
        );

    \I__1138\ : IoSpan4Mux
    port map (
            O => \N__6321\,
            I => \N__6318\
        );

    \I__1137\ : Sp12to4
    port map (
            O => \N__6318\,
            I => \N__6315\
        );

    \I__1136\ : Span12Mux_s7_v
    port map (
            O => \N__6315\,
            I => \N__6311\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6308\
        );

    \I__1134\ : Odrv12
    port map (
            O => \N__6311\,
            I => \BANK0_c\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6308\,
            I => \BANK0_c\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6303\,
            I => \N__6299\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6302\,
            I => \N__6296\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6299\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a5_0\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6296\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a5_0\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6287\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__6290\,
            I => \N__6283\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6287\,
            I => \N__6280\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6286\,
            I => \N__6277\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6283\,
            I => \N__6274\
        );

    \I__1123\ : Odrv4
    port map (
            O => \N__6280\,
            I => \U712_CHIP_RAM.N_186\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6277\,
            I => \U712_CHIP_RAM.N_186\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6274\,
            I => \U712_CHIP_RAM.N_186\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6264\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6264\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0\
        );

    \I__1118\ : InMux
    port map (
            O => \N__6261\,
            I => \N__6257\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6254\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6257\,
            I => \N__6251\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__6254\,
            I => \N__6247\
        );

    \I__1114\ : Span4Mux_v
    port map (
            O => \N__6251\,
            I => \N__6244\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6250\,
            I => \N__6241\
        );

    \I__1112\ : Span4Mux_h
    port map (
            O => \N__6247\,
            I => \N__6238\
        );

    \I__1111\ : Odrv4
    port map (
            O => \N__6244\,
            I => \U712_CHIP_RAM.N_341\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6241\,
            I => \U712_CHIP_RAM.N_341\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__6238\,
            I => \U712_CHIP_RAM.N_341\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6231\,
            I => \N__6228\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6228\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6222\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6222\,
            I => \U712_CHIP_RAM.N_331\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6219\,
            I => \N__6214\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6218\,
            I => \N__6211\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6208\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__6214\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6211\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6208\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6196\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6200\,
            I => \N__6193\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6190\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__6196\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6193\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6190\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__6183\,
            I => \U712_CHIP_RAM.N_331_cascade_\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6180\,
            I => \N__6175\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6179\,
            I => \N__6172\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6178\,
            I => \N__6169\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6175\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__6172\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6169\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1085\ : CascadeMux
    port map (
            O => \N__6162\,
            I => \N__6158\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6153\
        );

    \I__1083\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6150\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6147\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6156\,
            I => \N__6143\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__6153\,
            I => \N__6138\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__6150\,
            I => \N__6138\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6147\,
            I => \N__6135\
        );

    \I__1077\ : InMux
    port map (
            O => \N__6146\,
            I => \N__6130\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__6143\,
            I => \N__6125\
        );

    \I__1075\ : Span4Mux_v
    port map (
            O => \N__6138\,
            I => \N__6120\
        );

    \I__1074\ : Span4Mux_v
    port map (
            O => \N__6135\,
            I => \N__6120\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6134\,
            I => \N__6117\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6114\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__6130\,
            I => \N__6111\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6129\,
            I => \N__6106\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6128\,
            I => \N__6106\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__6125\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__6120\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6117\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__6114\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1064\ : Odrv4
    port map (
            O => \N__6111\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6106\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__6093\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6087\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6087\,
            I => \N__6082\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6086\,
            I => \N__6075\
        );

    \I__1058\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6075\
        );

    \I__1057\ : Span4Mux_h
    port map (
            O => \N__6082\,
            I => \N__6072\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6067\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6080\,
            I => \N__6067\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6075\,
            I => \U712_CHIP_RAM.N_337\
        );

    \I__1053\ : Odrv4
    port map (
            O => \N__6072\,
            I => \U712_CHIP_RAM.N_337\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6067\,
            I => \U712_CHIP_RAM.N_337\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6055\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6059\,
            I => \N__6052\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6058\,
            I => \N__6045\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6055\,
            I => \N__6040\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6052\,
            I => \N__6040\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6037\
        );

    \I__1045\ : InMux
    port map (
            O => \N__6050\,
            I => \N__6032\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6029\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6048\,
            I => \N__6025\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6045\,
            I => \N__6022\
        );

    \I__1041\ : Span4Mux_v
    port map (
            O => \N__6040\,
            I => \N__6017\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6037\,
            I => \N__6017\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6014\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6011\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6032\,
            I => \N__6006\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6029\,
            I => \N__6006\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6003\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6025\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1033\ : Odrv12
    port map (
            O => \N__6022\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1032\ : Odrv4
    port map (
            O => \N__6017\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6014\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6011\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1029\ : Odrv4
    port map (
            O => \N__6006\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__6003\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__5988\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5985\,
            I => \N__5982\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5982\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5979\,
            I => \bfn_11_12_0_\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5976\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5973\,
            I => \N__5970\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__5970\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5967\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5964\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__1018\ : CascadeMux
    port map (
            O => \N__5961\,
            I => \N__5956\
        );

    \I__1017\ : InMux
    port map (
            O => \N__5960\,
            I => \N__5953\
        );

    \I__1016\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5950\
        );

    \I__1015\ : InMux
    port map (
            O => \N__5956\,
            I => \N__5947\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5953\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5950\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5947\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5940\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5937\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5934\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__1008\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5915\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5930\,
            I => \N__5915\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5929\,
            I => \N__5915\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5928\,
            I => \N__5915\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5910\
        );

    \I__1003\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5910\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5905\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5924\,
            I => \N__5905\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5915\,
            I => \U712_CHIP_RAM.N_181\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5910\,
            I => \U712_CHIP_RAM.N_181\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5905\,
            I => \U712_CHIP_RAM.N_181\
        );

    \I__997\ : InMux
    port map (
            O => \N__5898\,
            I => \N__5895\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__5895\,
            I => \N__5892\
        );

    \I__995\ : Sp12to4
    port map (
            O => \N__5892\,
            I => \N__5889\
        );

    \I__994\ : Span12Mux_v
    port map (
            O => \N__5889\,
            I => \N__5886\
        );

    \I__993\ : Span12Mux_h
    port map (
            O => \N__5886\,
            I => \N__5883\
        );

    \I__992\ : Odrv12
    port map (
            O => \N__5883\,
            I => \A_c_5\
        );

    \I__991\ : InMux
    port map (
            O => \N__5880\,
            I => \N__5877\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5877\,
            I => \N__5874\
        );

    \I__989\ : Span4Mux_v
    port map (
            O => \N__5874\,
            I => \N__5871\
        );

    \I__988\ : Sp12to4
    port map (
            O => \N__5871\,
            I => \N__5868\
        );

    \I__987\ : Span12Mux_h
    port map (
            O => \N__5868\,
            I => \N__5865\
        );

    \I__986\ : Odrv12
    port map (
            O => \N__5865\,
            I => \A_c_12\
        );

    \I__985\ : InMux
    port map (
            O => \N__5862\,
            I => \N__5859\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5859\,
            I => \N__5856\
        );

    \I__983\ : Span4Mux_h
    port map (
            O => \N__5856\,
            I => \N__5853\
        );

    \I__982\ : Span4Mux_h
    port map (
            O => \N__5853\,
            I => \N__5850\
        );

    \I__981\ : Sp12to4
    port map (
            O => \N__5850\,
            I => \N__5847\
        );

    \I__980\ : Span12Mux_v
    port map (
            O => \N__5847\,
            I => \N__5844\
        );

    \I__979\ : Odrv12
    port map (
            O => \N__5844\,
            I => \A_c_16\
        );

    \I__978\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5838\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5838\,
            I => \N__5835\
        );

    \I__976\ : Span4Mux_v
    port map (
            O => \N__5835\,
            I => \N__5832\
        );

    \I__975\ : Sp12to4
    port map (
            O => \N__5832\,
            I => \N__5829\
        );

    \I__974\ : Span12Mux_h
    port map (
            O => \N__5829\,
            I => \N__5826\
        );

    \I__973\ : Span12Mux_v
    port map (
            O => \N__5826\,
            I => \N__5823\
        );

    \I__972\ : Odrv12
    port map (
            O => \N__5823\,
            I => \A_c_18\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__5820\,
            I => \N__5817\
        );

    \I__970\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5811\
        );

    \I__969\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5808\
        );

    \I__968\ : InMux
    port map (
            O => \N__5815\,
            I => \N__5805\
        );

    \I__967\ : InMux
    port map (
            O => \N__5814\,
            I => \N__5802\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5811\,
            I => \N__5797\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__5808\,
            I => \N__5797\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5805\,
            I => \N__5794\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__5802\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__962\ : Odrv4
    port map (
            O => \N__5797\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__961\ : Odrv12
    port map (
            O => \N__5794\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__5787\,
            I => \N__5784\
        );

    \I__959\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5781\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5781\,
            I => \N__5778\
        );

    \I__957\ : Span4Mux_v
    port map (
            O => \N__5778\,
            I => \N__5774\
        );

    \I__956\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5771\
        );

    \I__955\ : Span4Mux_h
    port map (
            O => \N__5774\,
            I => \N__5768\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5771\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__5768\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__5763\,
            I => \U712_CYCLE_TERM.N_211_i_0_en_cascade_\
        );

    \I__951\ : CEMux
    port map (
            O => \N__5760\,
            I => \N__5757\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__5757\,
            I => \N__5754\
        );

    \I__949\ : Odrv12
    port map (
            O => \N__5754\,
            I => \U712_CYCLE_TERM.N_211_i_0_en_0\
        );

    \I__948\ : InMux
    port map (
            O => \N__5751\,
            I => \N__5748\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__5748\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0\
        );

    \I__946\ : CEMux
    port map (
            O => \N__5745\,
            I => \N__5742\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5742\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0\
        );

    \I__944\ : CascadeMux
    port map (
            O => \N__5739\,
            I => \U712_CHIP_RAM.N_339_cascade_\
        );

    \I__943\ : InMux
    port map (
            O => \N__5736\,
            I => \N__5732\
        );

    \I__942\ : InMux
    port map (
            O => \N__5735\,
            I => \N__5727\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5732\,
            I => \N__5724\
        );

    \I__940\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5720\
        );

    \I__939\ : InMux
    port map (
            O => \N__5730\,
            I => \N__5717\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5727\,
            I => \N__5712\
        );

    \I__937\ : Span4Mux_h
    port map (
            O => \N__5724\,
            I => \N__5712\
        );

    \I__936\ : InMux
    port map (
            O => \N__5723\,
            I => \N__5709\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5720\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5717\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__5712\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__5709\,
            I => \U712_CHIP_RAM.N_335\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__5700\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_1_cascade_\
        );

    \I__930\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5693\
        );

    \I__929\ : InMux
    port map (
            O => \N__5696\,
            I => \N__5690\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5693\,
            I => \U712_CHIP_RAM.N_296\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__5690\,
            I => \U712_CHIP_RAM.N_296\
        );

    \I__926\ : CascadeMux
    port map (
            O => \N__5685\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_i_a5_0_1_cascade_\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__5682\,
            I => \U712_CHIP_RAM.N_257_cascade_\
        );

    \I__924\ : InMux
    port map (
            O => \N__5679\,
            I => \N__5676\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5676\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_i_0\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__5673\,
            I => \U712_CHIP_RAM.N_338_cascade_\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__5670\,
            I => \N__5658\
        );

    \I__920\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5655\
        );

    \I__919\ : InMux
    port map (
            O => \N__5668\,
            I => \N__5648\
        );

    \I__918\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5648\
        );

    \I__917\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5648\
        );

    \I__916\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5642\
        );

    \I__915\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5637\
        );

    \I__914\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5637\
        );

    \I__913\ : InMux
    port map (
            O => \N__5662\,
            I => \N__5632\
        );

    \I__912\ : InMux
    port map (
            O => \N__5661\,
            I => \N__5632\
        );

    \I__911\ : InMux
    port map (
            O => \N__5658\,
            I => \N__5629\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5655\,
            I => \N__5624\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5648\,
            I => \N__5624\
        );

    \I__908\ : InMux
    port map (
            O => \N__5647\,
            I => \N__5617\
        );

    \I__907\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5617\
        );

    \I__906\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5617\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5642\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5637\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5632\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5629\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__901\ : Odrv4
    port map (
            O => \N__5624\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__5617\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__899\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5601\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__5601\,
            I => \U712_CHIP_RAM.N_284_2\
        );

    \I__897\ : InMux
    port map (
            O => \N__5598\,
            I => \N__5594\
        );

    \I__896\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5591\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__5594\,
            I => \N__5588\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__5591\,
            I => \N__5585\
        );

    \I__893\ : Odrv4
    port map (
            O => \N__5588\,
            I => \U712_CHIP_RAM.N_253\
        );

    \I__892\ : Odrv4
    port map (
            O => \N__5585\,
            I => \U712_CHIP_RAM.N_253\
        );

    \I__891\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5577\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5577\,
            I => \N__5571\
        );

    \I__889\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5566\
        );

    \I__888\ : InMux
    port map (
            O => \N__5575\,
            I => \N__5566\
        );

    \I__887\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5563\
        );

    \I__886\ : Span4Mux_v
    port map (
            O => \N__5571\,
            I => \N__5556\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5566\,
            I => \N__5556\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5563\,
            I => \N__5556\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__5556\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__5553\,
            I => \U712_CHIP_RAM.N_284_2_cascade_\
        );

    \I__881\ : InMux
    port map (
            O => \N__5550\,
            I => \N__5547\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5547\,
            I => \U712_CHIP_RAM.N_254\
        );

    \I__879\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5541\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__5541\,
            I => \U712_CHIP_RAM.N_322\
        );

    \I__877\ : InMux
    port map (
            O => \N__5538\,
            I => \N__5535\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5535\,
            I => \N__5532\
        );

    \I__875\ : Odrv4
    port map (
            O => \N__5532\,
            I => \U712_CHIP_RAM.N_206\
        );

    \I__874\ : InMux
    port map (
            O => \N__5529\,
            I => \N__5525\
        );

    \I__873\ : InMux
    port map (
            O => \N__5528\,
            I => \N__5520\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5525\,
            I => \N__5517\
        );

    \I__871\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5512\
        );

    \I__870\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5512\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5520\,
            I => \U712_CHIP_RAM.N_338\
        );

    \I__868\ : Odrv4
    port map (
            O => \N__5517\,
            I => \U712_CHIP_RAM.N_338\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5512\,
            I => \U712_CHIP_RAM.N_338\
        );

    \I__866\ : InMux
    port map (
            O => \N__5505\,
            I => \N__5502\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5502\,
            I => \U712_CHIP_RAM.N_256\
        );

    \I__864\ : InMux
    port map (
            O => \N__5499\,
            I => \N__5496\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5496\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__5493\,
            I => \N__5490\
        );

    \I__861\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5487\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__5487\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__859\ : InMux
    port map (
            O => \N__5484\,
            I => \N__5481\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5481\,
            I => \U712_CHIP_RAM.N_284\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__5478\,
            I => \U712_CHIP_RAM.N_284_cascade_\
        );

    \I__856\ : InMux
    port map (
            O => \N__5475\,
            I => \N__5467\
        );

    \I__855\ : InMux
    port map (
            O => \N__5474\,
            I => \N__5467\
        );

    \I__854\ : InMux
    port map (
            O => \N__5473\,
            I => \N__5462\
        );

    \I__853\ : InMux
    port map (
            O => \N__5472\,
            I => \N__5462\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5467\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5462\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__5457\,
            I => \N__5453\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__5456\,
            I => \N__5450\
        );

    \I__848\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5445\
        );

    \I__847\ : InMux
    port map (
            O => \N__5450\,
            I => \N__5445\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5445\,
            I => \N__5440\
        );

    \I__845\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5437\
        );

    \I__844\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5434\
        );

    \I__843\ : Span4Mux_v
    port map (
            O => \N__5440\,
            I => \N__5429\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5437\,
            I => \N__5429\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5434\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__5429\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__839\ : InMux
    port map (
            O => \N__5424\,
            I => \N__5421\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5421\,
            I => \U712_CHIP_RAM.N_218\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__5418\,
            I => \U712_CHIP_RAM.N_218_cascade_\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__5415\,
            I => \N__5412\
        );

    \I__835\ : InMux
    port map (
            O => \N__5412\,
            I => \N__5409\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5409\,
            I => \N__5405\
        );

    \I__833\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5402\
        );

    \I__832\ : Odrv4
    port map (
            O => \N__5405\,
            I => \U712_CHIP_RAM.N_259\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5402\,
            I => \U712_CHIP_RAM.N_259\
        );

    \I__830\ : CascadeMux
    port map (
            O => \N__5397\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a2_0_a5_0_cascade_\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__5394\,
            I => \U712_CHIP_RAM.N_206_cascade_\
        );

    \I__828\ : InMux
    port map (
            O => \N__5391\,
            I => \N__5388\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5388\,
            I => \U712_CHIP_RAM.N_329\
        );

    \I__826\ : InMux
    port map (
            O => \N__5385\,
            I => \N__5382\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5382\,
            I => \N__5377\
        );

    \I__824\ : InMux
    port map (
            O => \N__5381\,
            I => \N__5374\
        );

    \I__823\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5371\
        );

    \I__822\ : Odrv4
    port map (
            O => \N__5377\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5374\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5371\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__5364\,
            I => \U712_CHIP_RAM.N_323_cascade_\
        );

    \I__818\ : InMux
    port map (
            O => \N__5361\,
            I => \N__5358\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5358\,
            I => \U712_CHIP_RAM.N_374\
        );

    \I__816\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5350\
        );

    \I__815\ : InMux
    port map (
            O => \N__5354\,
            I => \N__5345\
        );

    \I__814\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5345\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__5350\,
            I => \U712_CHIP_RAM.N_378\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5345\,
            I => \U712_CHIP_RAM.N_378\
        );

    \I__811\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5334\
        );

    \I__810\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5334\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__5334\,
            I => \U712_CHIP_RAM.N_184\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__5331\,
            I => \U712_CHIP_RAM.N_335_cascade_\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__5328\,
            I => \N__5324\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__5327\,
            I => \N__5321\
        );

    \I__805\ : InMux
    port map (
            O => \N__5324\,
            I => \N__5318\
        );

    \I__804\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5315\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5318\,
            I => \U712_CHIP_RAM.N_280\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5315\,
            I => \U712_CHIP_RAM.N_280\
        );

    \I__801\ : SRMux
    port map (
            O => \N__5310\,
            I => \N__5307\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__5307\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__799\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5300\
        );

    \I__798\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5297\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5300\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5297\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__795\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5288\
        );

    \I__794\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5285\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__5288\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5285\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__5280\,
            I => \N__5276\
        );

    \I__790\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5273\
        );

    \I__789\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5270\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5273\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5270\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__786\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5261\
        );

    \I__785\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5258\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__5261\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5258\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__782\ : InMux
    port map (
            O => \N__5253\,
            I => \N__5249\
        );

    \I__781\ : InMux
    port map (
            O => \N__5252\,
            I => \N__5246\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__5249\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5246\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__778\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5237\
        );

    \I__777\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5234\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5237\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5234\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__774\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5225\
        );

    \I__773\ : InMux
    port map (
            O => \N__5228\,
            I => \N__5222\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5225\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5222\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__770\ : InMux
    port map (
            O => \N__5217\,
            I => \N__5213\
        );

    \I__769\ : InMux
    port map (
            O => \N__5216\,
            I => \N__5210\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5213\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__5210\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__5205\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_\
        );

    \I__765\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5199\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5199\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__763\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5193\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__5193\,
            I => \U712_CHIP_RAM.N_340\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__5190\,
            I => \U712_CHIP_RAM.N_340_cascade_\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__5187\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\
        );

    \I__759\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5181\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5181\,
            I => \U712_CHIP_RAM.N_97\
        );

    \I__757\ : IoInMux
    port map (
            O => \N__5178\,
            I => \N__5175\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5175\,
            I => \N__5172\
        );

    \I__755\ : Span12Mux_s3_v
    port map (
            O => \N__5172\,
            I => \N__5169\
        );

    \I__754\ : Span12Mux_v
    port map (
            O => \N__5169\,
            I => \N__5165\
        );

    \I__753\ : InMux
    port map (
            O => \N__5168\,
            I => \N__5162\
        );

    \I__752\ : Odrv12
    port map (
            O => \N__5165\,
            I => \LATCH_CLK_c\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__5162\,
            I => \LATCH_CLK_c\
        );

    \I__750\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5152\
        );

    \I__749\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5148\
        );

    \I__748\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5145\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__5152\,
            I => \N__5142\
        );

    \I__746\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5139\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__5148\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5145\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__5142\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__5139\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__741\ : InMux
    port map (
            O => \N__5130\,
            I => \N__5127\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5127\,
            I => \U712_CYCLE_TERM.N_312\
        );

    \I__739\ : InMux
    port map (
            O => \N__5124\,
            I => \N__5121\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__5121\,
            I => \N__5118\
        );

    \I__737\ : Span12Mux_h
    port map (
            O => \N__5118\,
            I => \N__5115\
        );

    \I__736\ : Span12Mux_v
    port map (
            O => \N__5115\,
            I => \N__5112\
        );

    \I__735\ : Odrv12
    port map (
            O => \N__5112\,
            I => \A_c_3\
        );

    \I__734\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5106\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5106\,
            I => \N__5103\
        );

    \I__732\ : Span12Mux_v
    port map (
            O => \N__5103\,
            I => \N__5100\
        );

    \I__731\ : Span12Mux_h
    port map (
            O => \N__5100\,
            I => \N__5097\
        );

    \I__730\ : Odrv12
    port map (
            O => \N__5097\,
            I => \A_c_10\
        );

    \I__729\ : InMux
    port map (
            O => \N__5094\,
            I => \bfn_10_9_0_\
        );

    \I__728\ : InMux
    port map (
            O => \N__5091\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__727\ : InMux
    port map (
            O => \N__5088\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__726\ : InMux
    port map (
            O => \N__5085\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__725\ : InMux
    port map (
            O => \N__5082\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__724\ : InMux
    port map (
            O => \N__5079\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__723\ : InMux
    port map (
            O => \N__5076\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__722\ : InMux
    port map (
            O => \N__5073\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__721\ : ClkMux
    port map (
            O => \N__5070\,
            I => \N__5049\
        );

    \I__720\ : ClkMux
    port map (
            O => \N__5069\,
            I => \N__5049\
        );

    \I__719\ : ClkMux
    port map (
            O => \N__5068\,
            I => \N__5049\
        );

    \I__718\ : ClkMux
    port map (
            O => \N__5067\,
            I => \N__5049\
        );

    \I__717\ : ClkMux
    port map (
            O => \N__5066\,
            I => \N__5049\
        );

    \I__716\ : ClkMux
    port map (
            O => \N__5065\,
            I => \N__5049\
        );

    \I__715\ : ClkMux
    port map (
            O => \N__5064\,
            I => \N__5049\
        );

    \I__714\ : GlobalMux
    port map (
            O => \N__5049\,
            I => \N__5046\
        );

    \I__713\ : gio2CtrlBuf
    port map (
            O => \N__5046\,
            I => \C1_c_g\
        );

    \I__712\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5040\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5040\,
            I => \U712_CHIP_RAM.N_258\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__5037\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_\
        );

    \I__709\ : IoInMux
    port map (
            O => \N__5034\,
            I => \N__5031\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5031\,
            I => \N__5028\
        );

    \I__707\ : Span4Mux_s0_h
    port map (
            O => \N__5028\,
            I => \N__5025\
        );

    \I__706\ : Span4Mux_h
    port map (
            O => \N__5025\,
            I => \N__5022\
        );

    \I__705\ : Span4Mux_h
    port map (
            O => \N__5022\,
            I => \N__5019\
        );

    \I__704\ : Sp12to4
    port map (
            O => \N__5019\,
            I => \N__5016\
        );

    \I__703\ : Span12Mux_v
    port map (
            O => \N__5016\,
            I => \N__5013\
        );

    \I__702\ : Odrv12
    port map (
            O => \N__5013\,
            I => \N_235\
        );

    \I__701\ : InMux
    port map (
            O => \N__5010\,
            I => \N__5005\
        );

    \I__700\ : InMux
    port map (
            O => \N__5009\,
            I => \N__4999\
        );

    \I__699\ : InMux
    port map (
            O => \N__5008\,
            I => \N__4999\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5005\,
            I => \N__4996\
        );

    \I__697\ : InMux
    port map (
            O => \N__5004\,
            I => \N__4993\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__4999\,
            I => \N__4990\
        );

    \I__695\ : Span4Mux_v
    port map (
            O => \N__4996\,
            I => \N__4985\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4993\,
            I => \N__4985\
        );

    \I__693\ : Span4Mux_v
    port map (
            O => \N__4990\,
            I => \N__4982\
        );

    \I__692\ : Span4Mux_v
    port map (
            O => \N__4985\,
            I => \N__4979\
        );

    \I__691\ : Sp12to4
    port map (
            O => \N__4982\,
            I => \N__4974\
        );

    \I__690\ : Sp12to4
    port map (
            O => \N__4979\,
            I => \N__4974\
        );

    \I__689\ : Span12Mux_h
    port map (
            O => \N__4974\,
            I => \N__4971\
        );

    \I__688\ : Odrv12
    port map (
            O => \N__4971\,
            I => \RnW_c\
        );

    \I__687\ : InMux
    port map (
            O => \N__4968\,
            I => \N__4965\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4965\,
            I => \N__4961\
        );

    \I__685\ : InMux
    port map (
            O => \N__4964\,
            I => \N__4958\
        );

    \I__684\ : Span4Mux_v
    port map (
            O => \N__4961\,
            I => \N__4953\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4958\,
            I => \N__4953\
        );

    \I__682\ : Span4Mux_v
    port map (
            O => \N__4953\,
            I => \N__4950\
        );

    \I__681\ : Sp12to4
    port map (
            O => \N__4950\,
            I => \N__4947\
        );

    \I__680\ : Span12Mux_h
    port map (
            O => \N__4947\,
            I => \N__4944\
        );

    \I__679\ : Odrv12
    port map (
            O => \N__4944\,
            I => \AWEn_c\
        );

    \I__678\ : InMux
    port map (
            O => \N__4941\,
            I => \N__4938\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4938\,
            I => \U712_CHIP_RAM.N_222\
        );

    \I__676\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4932\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__4932\,
            I => \N__4929\
        );

    \I__674\ : Span4Mux_v
    port map (
            O => \N__4929\,
            I => \N__4926\
        );

    \I__673\ : Odrv4
    port map (
            O => \N__4926\,
            I => \U712_BYTE_ENABLE.N_217\
        );

    \I__672\ : IoInMux
    port map (
            O => \N__4923\,
            I => \N__4920\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4920\,
            I => \N__4917\
        );

    \I__670\ : Span4Mux_s3_v
    port map (
            O => \N__4917\,
            I => \N__4914\
        );

    \I__669\ : Span4Mux_h
    port map (
            O => \N__4914\,
            I => \N__4911\
        );

    \I__668\ : Span4Mux_v
    port map (
            O => \N__4911\,
            I => \N__4908\
        );

    \I__667\ : Odrv4
    port map (
            O => \N__4908\,
            I => \DMA_LATCH_EN_c\
        );

    \I__666\ : InMux
    port map (
            O => \N__4905\,
            I => \N__4902\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4902\,
            I => \N__4899\
        );

    \I__664\ : Span4Mux_v
    port map (
            O => \N__4899\,
            I => \N__4896\
        );

    \I__663\ : Sp12to4
    port map (
            O => \N__4896\,
            I => \N__4893\
        );

    \I__662\ : Span12Mux_h
    port map (
            O => \N__4893\,
            I => \N__4890\
        );

    \I__661\ : Odrv12
    port map (
            O => \N__4890\,
            I => \A_c_11\
        );

    \I__660\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4884\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__4884\,
            I => \N__4881\
        );

    \I__658\ : Span12Mux_v
    port map (
            O => \N__4881\,
            I => \N__4878\
        );

    \I__657\ : Span12Mux_h
    port map (
            O => \N__4878\,
            I => \N__4875\
        );

    \I__656\ : Odrv12
    port map (
            O => \N__4875\,
            I => \A_c_4\
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__4872\,
            I => \U712_CHIP_RAM.N_187_cascade_\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__4869\,
            I => \U712_CHIP_RAM.N_316_cascade_\
        );

    \I__653\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4863\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__4863\,
            I => \U712_CHIP_RAM.N_316\
        );

    \I__651\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4857\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4857\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a5_1\
        );

    \I__649\ : CascadeMux
    port map (
            O => \N__4854\,
            I => \U712_CHIP_RAM.N_283_cascade_\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__4851\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\
        );

    \I__647\ : InMux
    port map (
            O => \N__4848\,
            I => \N__4843\
        );

    \I__646\ : InMux
    port map (
            O => \N__4847\,
            I => \N__4838\
        );

    \I__645\ : InMux
    port map (
            O => \N__4846\,
            I => \N__4838\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4843\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4838\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__642\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4830\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__4830\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__4827\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_\
        );

    \I__639\ : CEMux
    port map (
            O => \N__4824\,
            I => \N__4821\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4821\,
            I => \N__4818\
        );

    \I__637\ : Span4Mux_v
    port map (
            O => \N__4818\,
            I => \N__4815\
        );

    \I__636\ : Span4Mux_h
    port map (
            O => \N__4815\,
            I => \N__4812\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__4812\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\
        );

    \I__634\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4806\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4806\,
            I => \N__4803\
        );

    \I__632\ : Span4Mux_h
    port map (
            O => \N__4803\,
            I => \N__4800\
        );

    \I__631\ : Span4Mux_v
    port map (
            O => \N__4800\,
            I => \N__4797\
        );

    \I__630\ : Span4Mux_v
    port map (
            O => \N__4797\,
            I => \N__4794\
        );

    \I__629\ : Span4Mux_v
    port map (
            O => \N__4794\,
            I => \N__4791\
        );

    \I__628\ : Odrv4
    port map (
            O => \N__4791\,
            I => \RAMSPACEn_c\
        );

    \I__627\ : InMux
    port map (
            O => \N__4788\,
            I => \N__4785\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__4785\,
            I => \N__4782\
        );

    \I__625\ : Span4Mux_v
    port map (
            O => \N__4782\,
            I => \N__4778\
        );

    \I__624\ : InMux
    port map (
            O => \N__4781\,
            I => \N__4775\
        );

    \I__623\ : Span4Mux_v
    port map (
            O => \N__4778\,
            I => \N__4772\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__4775\,
            I => \N__4769\
        );

    \I__621\ : Sp12to4
    port map (
            O => \N__4772\,
            I => \N__4766\
        );

    \I__620\ : Span12Mux_h
    port map (
            O => \N__4769\,
            I => \N__4763\
        );

    \I__619\ : Span12Mux_h
    port map (
            O => \N__4766\,
            I => \N__4760\
        );

    \I__618\ : Span12Mux_v
    port map (
            O => \N__4763\,
            I => \N__4757\
        );

    \I__617\ : Odrv12
    port map (
            O => \N__4760\,
            I => \TSn_c\
        );

    \I__616\ : Odrv12
    port map (
            O => \N__4757\,
            I => \TSn_c\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__4752\,
            I => \U712_CHIP_RAM.N_279_cascade_\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__4749\,
            I => \U712_BYTE_ENABLE.N_215_cascade_\
        );

    \I__613\ : IoInMux
    port map (
            O => \N__4746\,
            I => \N__4743\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4743\,
            I => \N__4740\
        );

    \I__611\ : Span12Mux_s11_v
    port map (
            O => \N__4740\,
            I => \N__4737\
        );

    \I__610\ : Odrv12
    port map (
            O => \N__4737\,
            I => \N_167_i\
        );

    \I__609\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4728\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__4733\,
            I => \N__4718\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__4732\,
            I => \N__4715\
        );

    \I__606\ : InMux
    port map (
            O => \N__4731\,
            I => \N__4712\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4728\,
            I => \N__4709\
        );

    \I__604\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4706\
        );

    \I__603\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4697\
        );

    \I__602\ : InMux
    port map (
            O => \N__4725\,
            I => \N__4697\
        );

    \I__601\ : InMux
    port map (
            O => \N__4724\,
            I => \N__4697\
        );

    \I__600\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4697\
        );

    \I__599\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4688\
        );

    \I__598\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4688\
        );

    \I__597\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4688\
        );

    \I__596\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4688\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4712\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__594\ : Odrv4
    port map (
            O => \N__4709\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4706\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__4697\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4688\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__590\ : IoInMux
    port map (
            O => \N__4677\,
            I => \N__4674\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4674\,
            I => \N__4670\
        );

    \I__588\ : IoInMux
    port map (
            O => \N__4673\,
            I => \N__4667\
        );

    \I__587\ : Span4Mux_s2_v
    port map (
            O => \N__4670\,
            I => \N__4664\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__4667\,
            I => \N__4661\
        );

    \I__585\ : Span4Mux_h
    port map (
            O => \N__4664\,
            I => \N__4658\
        );

    \I__584\ : IoSpan4Mux
    port map (
            O => \N__4661\,
            I => \N__4655\
        );

    \I__583\ : Span4Mux_v
    port map (
            O => \N__4658\,
            I => \N__4652\
        );

    \I__582\ : Span4Mux_s3_v
    port map (
            O => \N__4655\,
            I => \N__4649\
        );

    \I__581\ : Span4Mux_v
    port map (
            O => \N__4652\,
            I => \N__4646\
        );

    \I__580\ : Span4Mux_h
    port map (
            O => \N__4649\,
            I => \N__4643\
        );

    \I__579\ : Sp12to4
    port map (
            O => \N__4646\,
            I => \N__4640\
        );

    \I__578\ : Span4Mux_v
    port map (
            O => \N__4643\,
            I => \N__4637\
        );

    \I__577\ : Odrv12
    port map (
            O => \N__4640\,
            I => \ASn_c\
        );

    \I__576\ : Odrv4
    port map (
            O => \N__4637\,
            I => \ASn_c\
        );

    \I__575\ : CEMux
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4629\,
            I => \N__4626\
        );

    \I__573\ : Span4Mux_h
    port map (
            O => \N__4626\,
            I => \N__4623\
        );

    \I__572\ : Odrv4
    port map (
            O => \N__4623\,
            I => \U712_REG_SM.N_219_0_0\
        );

    \I__571\ : InMux
    port map (
            O => \N__4620\,
            I => \N__4617\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4617\,
            I => \N__4614\
        );

    \I__569\ : Sp12to4
    port map (
            O => \N__4614\,
            I => \N__4611\
        );

    \I__568\ : Span12Mux_v
    port map (
            O => \N__4611\,
            I => \N__4608\
        );

    \I__567\ : Span12Mux_h
    port map (
            O => \N__4608\,
            I => \N__4605\
        );

    \I__566\ : Odrv12
    port map (
            O => \N__4605\,
            I => \A_c_6\
        );

    \I__565\ : InMux
    port map (
            O => \N__4602\,
            I => \N__4599\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4599\,
            I => \N__4596\
        );

    \I__563\ : Span4Mux_v
    port map (
            O => \N__4596\,
            I => \N__4593\
        );

    \I__562\ : Sp12to4
    port map (
            O => \N__4593\,
            I => \N__4590\
        );

    \I__561\ : Odrv12
    port map (
            O => \N__4590\,
            I => \A_c_13\
        );

    \I__560\ : IoInMux
    port map (
            O => \N__4587\,
            I => \N__4584\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4584\,
            I => \N__4581\
        );

    \I__558\ : Span4Mux_s3_v
    port map (
            O => \N__4581\,
            I => \N__4578\
        );

    \I__557\ : Span4Mux_v
    port map (
            O => \N__4578\,
            I => \N__4575\
        );

    \I__556\ : Span4Mux_v
    port map (
            O => \N__4575\,
            I => \N__4572\
        );

    \I__555\ : Span4Mux_v
    port map (
            O => \N__4572\,
            I => \N__4568\
        );

    \I__554\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4565\
        );

    \I__553\ : Odrv4
    port map (
            O => \N__4568\,
            I => \DBDIR_c\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__4565\,
            I => \DBDIR_c\
        );

    \I__551\ : InMux
    port map (
            O => \N__4560\,
            I => \N__4555\
        );

    \I__550\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4550\
        );

    \I__549\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4550\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4555\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4550\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__546\ : IoInMux
    port map (
            O => \N__4545\,
            I => \N__4542\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__4542\,
            I => \N__4539\
        );

    \I__544\ : Span4Mux_s1_h
    port map (
            O => \N__4539\,
            I => \N__4536\
        );

    \I__543\ : Sp12to4
    port map (
            O => \N__4536\,
            I => \N__4533\
        );

    \I__542\ : Span12Mux_v
    port map (
            O => \N__4533\,
            I => \N__4529\
        );

    \I__541\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4526\
        );

    \I__540\ : Odrv12
    port map (
            O => \N__4529\,
            I => \TACK_OUTn\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4526\,
            I => \TACK_OUTn\
        );

    \I__538\ : IoInMux
    port map (
            O => \N__4521\,
            I => \N__4518\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__4518\,
            I => \N__4515\
        );

    \I__536\ : IoSpan4Mux
    port map (
            O => \N__4515\,
            I => \N__4512\
        );

    \I__535\ : Sp12to4
    port map (
            O => \N__4512\,
            I => \N__4509\
        );

    \I__534\ : Span12Mux_s7_h
    port map (
            O => \N__4509\,
            I => \N__4506\
        );

    \I__533\ : Span12Mux_h
    port map (
            O => \N__4506\,
            I => \N__4503\
        );

    \I__532\ : Odrv12
    port map (
            O => \N__4503\,
            I => \N_165_i\
        );

    \I__531\ : InMux
    port map (
            O => \N__4500\,
            I => \N__4497\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4497\,
            I => \N__4494\
        );

    \I__529\ : Span4Mux_v
    port map (
            O => \N__4494\,
            I => \N__4490\
        );

    \I__528\ : InMux
    port map (
            O => \N__4493\,
            I => \N__4487\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__4490\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0Z0Z_0\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__4487\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0Z0Z_0\
        );

    \I__525\ : CascadeMux
    port map (
            O => \N__4482\,
            I => \N__4479\
        );

    \I__524\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4476\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4476\,
            I => \N__4473\
        );

    \I__522\ : Span4Mux_h
    port map (
            O => \N__4473\,
            I => \N__4470\
        );

    \I__521\ : Span4Mux_h
    port map (
            O => \N__4470\,
            I => \N__4467\
        );

    \I__520\ : Sp12to4
    port map (
            O => \N__4467\,
            I => \N__4464\
        );

    \I__519\ : Span12Mux_v
    port map (
            O => \N__4464\,
            I => \N__4461\
        );

    \I__518\ : Odrv12
    port map (
            O => \N__4461\,
            I => \REGSPACEn_c\
        );

    \I__517\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4455\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4455\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_i_i_0\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__4452\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_i_i_0_cascade_\
        );

    \I__514\ : InMux
    port map (
            O => \N__4449\,
            I => \N__4446\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4446\,
            I => \U712_CHIP_RAM.N_23\
        );

    \I__512\ : InMux
    port map (
            O => \N__4443\,
            I => \N__4439\
        );

    \I__511\ : InMux
    port map (
            O => \N__4442\,
            I => \N__4436\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__4439\,
            I => \U712_REG_SM.N_219\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4436\,
            I => \U712_REG_SM.N_219\
        );

    \I__508\ : InMux
    port map (
            O => \N__4431\,
            I => \N__4424\
        );

    \I__507\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4424\
        );

    \I__506\ : InMux
    port map (
            O => \N__4429\,
            I => \N__4421\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4424\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__4421\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__503\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4413\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4413\,
            I => \U712_REG_SM.N_261\
        );

    \I__501\ : InMux
    port map (
            O => \N__4410\,
            I => \N__4407\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4407\,
            I => \U712_REG_SM.DS_EN_RNOZ0Z_0\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__4404\,
            I => \N__4401\
        );

    \I__498\ : InMux
    port map (
            O => \N__4401\,
            I => \N__4393\
        );

    \I__497\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4388\
        );

    \I__496\ : InMux
    port map (
            O => \N__4399\,
            I => \N__4388\
        );

    \I__495\ : InMux
    port map (
            O => \N__4398\,
            I => \N__4385\
        );

    \I__494\ : InMux
    port map (
            O => \N__4397\,
            I => \N__4380\
        );

    \I__493\ : InMux
    port map (
            O => \N__4396\,
            I => \N__4380\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__4393\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4388\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4385\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4380\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__488\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4367\
        );

    \I__487\ : InMux
    port map (
            O => \N__4370\,
            I => \N__4364\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__4367\,
            I => \N__4361\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__4364\,
            I => \N__4358\
        );

    \I__484\ : Span4Mux_v
    port map (
            O => \N__4361\,
            I => \N__4355\
        );

    \I__483\ : Span4Mux_v
    port map (
            O => \N__4358\,
            I => \N__4352\
        );

    \I__482\ : Sp12to4
    port map (
            O => \N__4355\,
            I => \N__4349\
        );

    \I__481\ : Span4Mux_h
    port map (
            O => \N__4352\,
            I => \N__4346\
        );

    \I__480\ : Span12Mux_h
    port map (
            O => \N__4349\,
            I => \N__4341\
        );

    \I__479\ : Sp12to4
    port map (
            O => \N__4346\,
            I => \N__4341\
        );

    \I__478\ : Odrv12
    port map (
            O => \N__4341\,
            I => \DBRn_c\
        );

    \I__477\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4335\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4335\,
            I => \N__4332\
        );

    \I__475\ : Odrv4
    port map (
            O => \N__4332\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__474\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4326\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__4326\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__472\ : InMux
    port map (
            O => \N__4323\,
            I => \N__4319\
        );

    \I__471\ : InMux
    port map (
            O => \N__4322\,
            I => \N__4310\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__4319\,
            I => \N__4307\
        );

    \I__469\ : InMux
    port map (
            O => \N__4318\,
            I => \N__4304\
        );

    \I__468\ : InMux
    port map (
            O => \N__4317\,
            I => \N__4299\
        );

    \I__467\ : InMux
    port map (
            O => \N__4316\,
            I => \N__4299\
        );

    \I__466\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4292\
        );

    \I__465\ : InMux
    port map (
            O => \N__4314\,
            I => \N__4292\
        );

    \I__464\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4292\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4310\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__462\ : Odrv4
    port map (
            O => \N__4307\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4304\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4299\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4292\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__458\ : InMux
    port map (
            O => \N__4281\,
            I => \N__4277\
        );

    \I__457\ : IoInMux
    port map (
            O => \N__4280\,
            I => \N__4274\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__4277\,
            I => \N__4271\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4274\,
            I => \N__4268\
        );

    \I__454\ : Span4Mux_v
    port map (
            O => \N__4271\,
            I => \N__4265\
        );

    \I__453\ : IoSpan4Mux
    port map (
            O => \N__4268\,
            I => \N__4262\
        );

    \I__452\ : Sp12to4
    port map (
            O => \N__4265\,
            I => \N__4259\
        );

    \I__451\ : IoSpan4Mux
    port map (
            O => \N__4262\,
            I => \N__4256\
        );

    \I__450\ : Span12Mux_h
    port map (
            O => \N__4259\,
            I => \N__4253\
        );

    \I__449\ : IoSpan4Mux
    port map (
            O => \N__4256\,
            I => \N__4250\
        );

    \I__448\ : Odrv12
    port map (
            O => \N__4253\,
            I => \C1_c\
        );

    \I__447\ : Odrv4
    port map (
            O => \N__4250\,
            I => \C1_c\
        );

    \I__446\ : InMux
    port map (
            O => \N__4245\,
            I => \N__4242\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__4242\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__444\ : IoInMux
    port map (
            O => \N__4239\,
            I => \N__4236\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4236\,
            I => \N__4233\
        );

    \I__442\ : Span12Mux_s11_v
    port map (
            O => \N__4233\,
            I => \N__4230\
        );

    \I__441\ : Odrv12
    port map (
            O => \N__4230\,
            I => \VBENn_c\
        );

    \I__440\ : InMux
    port map (
            O => \N__4227\,
            I => \N__4221\
        );

    \I__439\ : InMux
    port map (
            O => \N__4226\,
            I => \N__4221\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__4221\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__437\ : CascadeMux
    port map (
            O => \N__4218\,
            I => \N__4215\
        );

    \I__436\ : InMux
    port map (
            O => \N__4215\,
            I => \N__4212\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__4212\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a5_0_0_0\
        );

    \I__434\ : InMux
    port map (
            O => \N__4209\,
            I => \N__4204\
        );

    \I__433\ : InMux
    port map (
            O => \N__4208\,
            I => \N__4199\
        );

    \I__432\ : InMux
    port map (
            O => \N__4207\,
            I => \N__4199\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__4204\,
            I => \U712_REG_SM.N_209\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__4199\,
            I => \U712_REG_SM.N_209\
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__4194\,
            I => \U712_REG_SM.STATE_COUNTc_1_0_cascade_\
        );

    \I__428\ : CascadeMux
    port map (
            O => \N__4191\,
            I => \U712_REG_SM.N_272_cascade_\
        );

    \I__427\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4180\
        );

    \I__426\ : InMux
    port map (
            O => \N__4187\,
            I => \N__4173\
        );

    \I__425\ : InMux
    port map (
            O => \N__4186\,
            I => \N__4173\
        );

    \I__424\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4173\
        );

    \I__423\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4170\
        );

    \I__422\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4167\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__4180\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__4173\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__4170\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__4167\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__417\ : CascadeMux
    port map (
            O => \N__4158\,
            I => \N__4155\
        );

    \I__416\ : InMux
    port map (
            O => \N__4155\,
            I => \N__4143\
        );

    \I__415\ : InMux
    port map (
            O => \N__4154\,
            I => \N__4143\
        );

    \I__414\ : InMux
    port map (
            O => \N__4153\,
            I => \N__4143\
        );

    \I__413\ : InMux
    port map (
            O => \N__4152\,
            I => \N__4143\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__4143\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__411\ : InMux
    port map (
            O => \N__4140\,
            I => \N__4137\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__4137\,
            I => \U712_REG_SM.STATE_COUNT_srsts_i_0_a5_0_0_0\
        );

    \I__409\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4131\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__4131\,
            I => \N__4127\
        );

    \I__407\ : InMux
    port map (
            O => \N__4130\,
            I => \N__4124\
        );

    \I__406\ : Odrv4
    port map (
            O => \N__4127\,
            I => \U712_REG_SM.N_207\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__4124\,
            I => \U712_REG_SM.N_207\
        );

    \I__404\ : CascadeMux
    port map (
            O => \N__4119\,
            I => \N__4114\
        );

    \I__403\ : CascadeMux
    port map (
            O => \N__4118\,
            I => \N__4109\
        );

    \I__402\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4105\
        );

    \I__401\ : InMux
    port map (
            O => \N__4114\,
            I => \N__4102\
        );

    \I__400\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4099\
        );

    \I__399\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4096\
        );

    \I__398\ : InMux
    port map (
            O => \N__4109\,
            I => \N__4091\
        );

    \I__397\ : InMux
    port map (
            O => \N__4108\,
            I => \N__4091\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__4105\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4102\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__4099\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__4096\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__4091\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__391\ : InMux
    port map (
            O => \N__4080\,
            I => \N__4077\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__4077\,
            I => \U712_REG_SM.N_191\
        );

    \I__389\ : InMux
    port map (
            O => \N__4074\,
            I => \N__4071\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__4071\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__387\ : CascadeMux
    port map (
            O => \N__4068\,
            I => \U712_REG_SM.N_191_cascade_\
        );

    \I__386\ : IoInMux
    port map (
            O => \N__4065\,
            I => \N__4062\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__4062\,
            I => \N__4059\
        );

    \I__384\ : IoSpan4Mux
    port map (
            O => \N__4059\,
            I => \N__4056\
        );

    \I__383\ : Span4Mux_s3_h
    port map (
            O => \N__4056\,
            I => \N__4053\
        );

    \I__382\ : Span4Mux_v
    port map (
            O => \N__4053\,
            I => \N__4050\
        );

    \I__381\ : Span4Mux_h
    port map (
            O => \N__4050\,
            I => \N__4047\
        );

    \I__380\ : Sp12to4
    port map (
            O => \N__4047\,
            I => \N__4043\
        );

    \I__379\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4040\
        );

    \I__378\ : Span12Mux_h
    port map (
            O => \N__4043\,
            I => \N__4035\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__4040\,
            I => \N__4035\
        );

    \I__376\ : Span12Mux_h
    port map (
            O => \N__4035\,
            I => \N__4032\
        );

    \I__375\ : Odrv12
    port map (
            O => \N__4032\,
            I => \C3_c\
        );

    \I__374\ : InMux
    port map (
            O => \N__4029\,
            I => \N__4026\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__4026\,
            I => \U712_REG_SM.N_85\
        );

    \I__372\ : InMux
    port map (
            O => \N__4023\,
            I => \N__4020\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__4020\,
            I => \N__4017\
        );

    \I__370\ : Odrv4
    port map (
            O => \N__4017\,
            I => \U712_REG_SM.N_263\
        );

    \I__369\ : IoInMux
    port map (
            O => \N__4014\,
            I => \N__4011\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__4011\,
            I => \N__4008\
        );

    \I__367\ : Span12Mux_s8_h
    port map (
            O => \N__4008\,
            I => \N__4005\
        );

    \I__366\ : Odrv12
    port map (
            O => \N__4005\,
            I => \N_812_i\
        );

    \I__365\ : InMux
    port map (
            O => \N__4002\,
            I => \N__3999\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3999\,
            I => \N__3996\
        );

    \I__363\ : Span4Mux_v
    port map (
            O => \N__3996\,
            I => \N__3993\
        );

    \I__362\ : Odrv4
    port map (
            O => \N__3993\,
            I => \TACK_EN_i_ess\
        );

    \I__361\ : IoInMux
    port map (
            O => \N__3990\,
            I => \N__3987\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3987\,
            I => \N__3984\
        );

    \I__359\ : IoSpan4Mux
    port map (
            O => \N__3984\,
            I => \N__3981\
        );

    \I__358\ : Span4Mux_s3_h
    port map (
            O => \N__3981\,
            I => \N__3978\
        );

    \I__357\ : Span4Mux_h
    port map (
            O => \N__3978\,
            I => \N__3975\
        );

    \I__356\ : Odrv4
    port map (
            O => \N__3975\,
            I => \DBRn_c_i_0\
        );

    \I__355\ : CascadeMux
    port map (
            O => \N__3972\,
            I => \U712_REG_SM.N_266_cascade_\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__3969\,
            I => \U712_REG_SM.N_269_cascade_\
        );

    \I__353\ : InMux
    port map (
            O => \N__3966\,
            I => \N__3962\
        );

    \I__352\ : InMux
    port map (
            O => \N__3965\,
            I => \N__3959\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3962\,
            I => \U712_REG_SM.N_233\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__3959\,
            I => \U712_REG_SM.N_233\
        );

    \I__349\ : IoInMux
    port map (
            O => \N__3954\,
            I => \N__3951\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3951\,
            I => \N__3948\
        );

    \I__347\ : Span4Mux_s2_v
    port map (
            O => \N__3948\,
            I => \N__3945\
        );

    \I__346\ : Span4Mux_v
    port map (
            O => \N__3945\,
            I => \N__3942\
        );

    \I__345\ : Odrv4
    port map (
            O => \N__3942\,
            I => \CLK80_PLL_i_i\
        );

    \I__344\ : IoInMux
    port map (
            O => \N__3939\,
            I => \N__3936\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3936\,
            I => \N__3933\
        );

    \I__342\ : IoSpan4Mux
    port map (
            O => \N__3933\,
            I => \N__3930\
        );

    \I__341\ : Span4Mux_s2_v
    port map (
            O => \N__3930\,
            I => \N__3927\
        );

    \I__340\ : Sp12to4
    port map (
            O => \N__3927\,
            I => \N__3924\
        );

    \I__339\ : Span12Mux_v
    port map (
            O => \N__3924\,
            I => \N__3921\
        );

    \I__338\ : Odrv12
    port map (
            O => \N__3921\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__5067\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__5068\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__5070\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__5064\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__5066\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__5065\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_9_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7590\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4280\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3990\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4065\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9663\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4002\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_812_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__7741\,
            in1 => \N__5814\,
            in2 => \_gnd_net_\,
            in3 => \N__7448\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9648\,
            ce => \N__5760\,
            sr => \N__10812\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10848\,
            in2 => \_gnd_net_\,
            in3 => \N__10460\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__5010\,
            in1 => \N__4113\,
            in2 => \_gnd_net_\,
            in3 => \N__3965\,
            lcout => \U712_REG_SM.N_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4400\,
            in1 => \N__4208\,
            in2 => \_gnd_net_\,
            in3 => \N__4725\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_266_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011100010"
        )
    port map (
            in0 => \N__10653\,
            in1 => \N__7780\,
            in2 => \N__3972\,
            in3 => \N__3966\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000101"
        )
    port map (
            in0 => \N__4399\,
            in1 => \_gnd_net_\,
            in2 => \N__4118\,
            in3 => \N__4207\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_269_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100000000"
        )
    port map (
            in0 => \N__4726\,
            in1 => \N__4323\,
            in2 => \N__3969\,
            in3 => \N__7781\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9654\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__4108\,
            in1 => \N__4724\,
            in2 => \_gnd_net_\,
            in3 => \N__4317\,
            lcout => \U712_REG_SM.N_263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__4184\,
            in1 => \N__4316\,
            in2 => \_gnd_net_\,
            in3 => \N__4723\,
            lcout => \U712_REG_SM.N_233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__4185\,
            in1 => \N__5004\,
            in2 => \_gnd_net_\,
            in3 => \N__4398\,
            lcout => \U712_REG_SM.DS_EN_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4370\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__4186\,
            in1 => \N__4318\,
            in2 => \_gnd_net_\,
            in3 => \N__4727\,
            lcout => \U712_REG_SM.N_191\,
            ltout => \U712_REG_SM.N_191_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__4117\,
            in1 => \N__7782\,
            in2 => \N__4068\,
            in3 => \N__4187\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9656\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4046\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9659\,
            ce => 'H',
            sr => \N__10783\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001000100010"
        )
    port map (
            in0 => \N__5777\,
            in1 => \N__5157\,
            in2 => \N__4218\,
            in3 => \N__7449\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9644\,
            ce => 'H',
            sr => \N__10805\
        );

    \U712_REG_SM.REG_TACK_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__4134\,
            in1 => \N__4029\,
            in2 => \N__7473\,
            in3 => \N__4023\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9644\,
            ce => 'H',
            sr => \N__10805\
        );

    \DBR_SYNC_1_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4338\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9649\,
            ce => 'H',
            sr => \N__10799\
        );

    \U712_REG_SM.STATE_COUNT_RNINRSB_1_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4153\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4396\,
            lcout => \U712_REG_SM.N_207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4314\,
            in2 => \_gnd_net_\,
            in3 => \N__5443\,
            lcout => \U712_REG_SM.N_209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101111"
        )
    port map (
            in0 => \N__4315\,
            in1 => \N__4721\,
            in2 => \N__4158\,
            in3 => \N__4397\,
            lcout => OPEN,
            ltout => \U712_REG_SM.STATE_COUNTc_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__7779\,
            in1 => \N__4209\,
            in2 => \N__4194\,
            in3 => \N__4731\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4188\,
            in1 => \N__4431\,
            in2 => \_gnd_net_\,
            in3 => \N__4112\,
            lcout => \U712_REG_SM.STATE_COUNT_srsts_i_0_a5_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__4430\,
            in1 => \N__4154\,
            in2 => \N__4733\,
            in3 => \N__4074\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_272_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__7778\,
            in1 => \N__4322\,
            in2 => \N__4191\,
            in3 => \N__4722\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9653\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIVCF31_1_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__4183\,
            in1 => \N__4313\,
            in2 => \N__4732\,
            in3 => \N__4152\,
            lcout => \U712_REG_SM.N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001000100011"
        )
    port map (
            in0 => \N__4140\,
            in1 => \N__4130\,
            in2 => \N__4119\,
            in3 => \N__4080\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9655\,
            ce => 'H',
            sr => \N__10784\
        );

    \U712_REG_SM.C1_SYNC_1_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4245\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9655\,
            ce => 'H',
            sr => \N__10784\
        );

    \U712_REG_SM.DS_EN_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000110011"
        )
    port map (
            in0 => \N__7819\,
            in1 => \N__4410\,
            in2 => \N__4404\,
            in3 => \N__4443\,
            lcout => \DS_ENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9655\,
            ce => 'H',
            sr => \N__10784\
        );

    \DBR_SYNC_0_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4371\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9655\,
            ce => 'H',
            sr => \N__10784\
        );

    \U712_REG_SM.C3_SYNC_1_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4329\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9655\,
            ce => 'H',
            sr => \N__10784\
        );

    \U712_REG_SM.C1_SYNC_0_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4281\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9657\,
            ce => 'H',
            sr => \N__10773\
        );

    \U712_BUFFERS.un1_VBENn_0_a5_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9369\,
            in2 => \_gnd_net_\,
            in3 => \N__10673\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7749\,
            in1 => \N__6867\,
            in2 => \_gnd_net_\,
            in3 => \N__5156\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4227\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7750\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4559\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7751\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9637\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4558\,
            in2 => \_gnd_net_\,
            in3 => \N__4226\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a5_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__4833\,
            in1 => \N__6984\,
            in2 => \N__6162\,
            in3 => \N__8952\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9640\,
            ce => 'H',
            sr => \N__10800\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5665\,
            in1 => \N__6060\,
            in2 => \_gnd_net_\,
            in3 => \N__6161\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9645\,
            ce => \N__4824\,
            sr => \N__10789\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000010001"
        )
    port map (
            in0 => \N__5043\,
            in1 => \N__4458\,
            in2 => \N__9733\,
            in3 => \N__4847\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__4846\,
            in1 => \N__4449\,
            in2 => \_gnd_net_\,
            in3 => \N__8432\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000010"
        )
    port map (
            in0 => \N__7748\,
            in1 => \N__4781\,
            in2 => \N__4482\,
            in3 => \N__4416\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_0_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6059\,
            in1 => \N__6146\,
            in2 => \_gnd_net_\,
            in3 => \N__10443\,
            lcout => \U712_CHIP_RAM.N_288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIE24B8_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__5597\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6090\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_i_i_0\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_i_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5529\,
            in2 => \N__4452\,
            in3 => \N__5736\,
            lcout => \U712_CHIP_RAM.N_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10845\,
            in2 => \_gnd_net_\,
            in3 => \N__4442\,
            lcout => \U712_REG_SM.N_219_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4429\,
            in2 => \_gnd_net_\,
            in3 => \N__10666\,
            lcout => \U712_REG_SM.N_261\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_i_o5_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110111100101"
        )
    port map (
            in0 => \N__8639\,
            in1 => \N__8816\,
            in2 => \N__8606\,
            in3 => \N__8728\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_167_i_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__4500\,
            in1 => \N__10544\,
            in2 => \N__4749\,
            in3 => \N__9392\,
            lcout => \N_167_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4734\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9658\,
            ce => \N__4632\,
            sr => \N__10770\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4620\,
            in1 => \N__4602\,
            in2 => \_gnd_net_\,
            in3 => \N__9104\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__8373\,
            in1 => \N__9734\,
            in2 => \N__8457\,
            in3 => \N__9127\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__4968\,
            in1 => \N__4571\,
            in2 => \_gnd_net_\,
            in3 => \N__5385\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9634\,
            ce => 'H',
            sr => \N__10801\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__4532\,
            in1 => \N__4560\,
            in2 => \N__6866\,
            in3 => \N__5155\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9634\,
            ce => 'H',
            sr => \N__10801\
        );

    \U712_BYTE_ENABLE.N_165_i_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111110101"
        )
    port map (
            in0 => \N__4493\,
            in1 => \N__4935\,
            in2 => \N__10628\,
            in3 => \N__9379\,
            lcout => \N_165_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7037\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6985\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_a5_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIALFTC_2_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__5196\,
            in1 => \N__6663\,
            in2 => \N__5327\,
            in3 => \N__5380\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4827\,
            in3 => \N__10846\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__7646\,
            in1 => \N__6849\,
            in2 => \N__5820\,
            in3 => \N__5130\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9638\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7036\,
            in2 => \_gnd_net_\,
            in3 => \N__7160\,
            lcout => \U712_CHIP_RAM.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHFLS1_1_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__7241\,
            in1 => \N__7746\,
            in2 => \N__6573\,
            in3 => \N__7148\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9383\,
            in2 => \_gnd_net_\,
            in3 => \N__5473\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__4809\,
            in1 => \N__4788\,
            in2 => \N__4752\,
            in3 => \N__7743\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9641\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5444\,
            in1 => \N__5472\,
            in2 => \_gnd_net_\,
            in3 => \N__5574\,
            lcout => \U712_CHIP_RAM.N_341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_1_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001000100"
        )
    port map (
            in0 => \N__6645\,
            in1 => \N__7147\,
            in2 => \N__7247\,
            in3 => \N__6550\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_187_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7745\,
            in1 => \N__5661\,
            in2 => \N__4872\,
            in3 => \N__7273\,
            lcout => \U712_CHIP_RAM.N_253\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI57LV_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7029\,
            in1 => \N__6641\,
            in2 => \_gnd_net_\,
            in3 => \N__6549\,
            lcout => \U712_CHIP_RAM.N_329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__7744\,
            in1 => \N__5355\,
            in2 => \N__6662\,
            in3 => \N__5662\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9641\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_1_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__7248\,
            in1 => \N__7159\,
            in2 => \N__6576\,
            in3 => \N__6737\,
            lcout => \U712_CHIP_RAM.N_316\,
            ltout => \U712_CHIP_RAM.N_316_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4HBB7_2_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__6635\,
            in1 => \_gnd_net_\,
            in2 => \N__4869\,
            in3 => \N__5353\,
            lcout => \U712_CHIP_RAM.N_259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQQ7R7_1_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__5354\,
            in1 => \N__5523\,
            in2 => \_gnd_net_\,
            in3 => \N__4866\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_283_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVVPHH_1_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__6738\,
            in1 => \N__4860\,
            in2 => \N__4854\,
            in3 => \N__5484\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5544\,
            in2 => \N__4851\,
            in3 => \N__9078\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__5679\,
            in1 => \N__4848\,
            in2 => \N__8389\,
            in3 => \N__5505\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9646\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNILSA11_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6634\,
            in2 => \N__6575\,
            in3 => \N__7392\,
            lcout => \U712_CHIP_RAM.N_184\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5524\,
            in1 => \N__6571\,
            in2 => \_gnd_net_\,
            in3 => \N__5731\,
            lcout => \U712_CHIP_RAM.N_258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6286\,
            in1 => \N__5669\,
            in2 => \_gnd_net_\,
            in3 => \N__6157\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__7404\,
            in1 => \N__4941\,
            in2 => \N__5037\,
            in3 => \N__7747\,
            lcout => \WRITE_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9651\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_0_m2_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001100110011"
        )
    port map (
            in0 => \N__5008\,
            in1 => \N__7405\,
            in2 => \N__10620\,
            in3 => \N__10543\,
            lcout => \N_235\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__5009\,
            in1 => \N__4964\,
            in2 => \_gnd_net_\,
            in3 => \N__6051\,
            lcout => \U712_CHIP_RAM.N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LMBE_i_o5_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001001111"
        )
    port map (
            in0 => \N__8746\,
            in1 => \N__8843\,
            in2 => \N__8607\,
            in3 => \N__8678\,
            lcout => \U712_BYTE_ENABLE.N_217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DMA_LATCH_EN_0_a5_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__10596\,
            in1 => \N__10518\,
            in2 => \_gnd_net_\,
            in3 => \N__7419\,
            lcout => \DMA_LATCH_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9154\,
            in1 => \N__4905\,
            in2 => \_gnd_net_\,
            in3 => \N__4887\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5124\,
            in1 => \N__5109\,
            in2 => \_gnd_net_\,
            in3 => \N__9153\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5304\,
            in2 => \_gnd_net_\,
            in3 => \N__5094\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__5069\,
            ce => 'H',
            sr => \N__5310\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5292\,
            in2 => \_gnd_net_\,
            in3 => \N__5091\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__5069\,
            ce => 'H',
            sr => \N__5310\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5265\,
            in2 => \_gnd_net_\,
            in3 => \N__5088\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__5069\,
            ce => 'H',
            sr => \N__5310\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5217\,
            in2 => \_gnd_net_\,
            in3 => \N__5085\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__5069\,
            ce => 'H',
            sr => \N__5310\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5279\,
            in2 => \_gnd_net_\,
            in3 => \N__5082\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__5069\,
            ce => 'H',
            sr => \N__5310\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5229\,
            in2 => \_gnd_net_\,
            in3 => \N__5079\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__5069\,
            ce => 'H',
            sr => \N__5310\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5241\,
            in2 => \_gnd_net_\,
            in3 => \N__5076\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__5069\,
            ce => 'H',
            sr => \N__5310\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5253\,
            in2 => \_gnd_net_\,
            in3 => \N__5073\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5069\,
            ce => 'H',
            sr => \N__5310\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101111111"
        )
    port map (
            in0 => \N__5303\,
            in1 => \N__5291\,
            in2 => \N__5280\,
            in3 => \N__5264\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5252\,
            in1 => \N__5240\,
            in2 => \_gnd_net_\,
            in3 => \N__5228\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010001010"
        )
    port map (
            in0 => \N__7752\,
            in1 => \N__5216\,
            in2 => \N__5205\,
            in3 => \N__5202\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9632\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__6049\,
            in1 => \_gnd_net_\,
            in2 => \N__5670\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7056\,
            in1 => \N__6739\,
            in2 => \N__6674\,
            in3 => \N__6700\,
            lcout => \U712_CHIP_RAM.N_340\,
            ltout => \U712_CHIP_RAM.N_340_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5381\,
            in2 => \N__5190\,
            in3 => \N__5697\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100011001000"
        )
    port map (
            in0 => \N__5168\,
            in1 => \N__7645\,
            in2 => \N__5187\,
            in3 => \N__5184\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9635\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110111"
        )
    port map (
            in0 => \N__7472\,
            in1 => \N__5816\,
            in2 => \N__7362\,
            in3 => \N__5151\,
            lcout => \U712_CYCLE_TERM.N_312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIM4DI_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7420\,
            in2 => \_gnd_net_\,
            in3 => \N__6572\,
            lcout => \U712_CHIP_RAM.N_206\,
            ltout => \U712_CHIP_RAM.N_206_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_3_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6661\,
            in1 => \N__7229\,
            in2 => \N__5394\,
            in3 => \N__5723\,
            lcout => \U712_CHIP_RAM.N_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOJRU2_1_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__7225\,
            in1 => \N__5340\,
            in2 => \N__7155\,
            in3 => \N__5391\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6050\,
            in1 => \N__5647\,
            in2 => \_gnd_net_\,
            in3 => \N__6128\,
            lcout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6199\,
            in1 => \N__6178\,
            in2 => \N__5961\,
            in3 => \N__6217\,
            lcout => \U712_CHIP_RAM.N_323\,
            ltout => \U712_CHIP_RAM.N_323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5364\,
            in3 => \N__5645\,
            lcout => \U712_CHIP_RAM.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__6129\,
            in1 => \N__5361\,
            in2 => \N__5328\,
            in3 => \N__6250\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7272\,
            in1 => \N__7224\,
            in2 => \N__7146\,
            in3 => \N__6554\,
            lcout => \U712_CHIP_RAM.N_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5646\,
            in1 => \N__7271\,
            in2 => \_gnd_net_\,
            in3 => \N__7123\,
            lcout => \U712_CHIP_RAM.N_335\,
            ltout => \U712_CHIP_RAM.N_335_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_3_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__5339\,
            in1 => \_gnd_net_\,
            in2 => \N__5331\,
            in3 => \N__7223\,
            lcout => \U712_CHIP_RAM.N_280\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__5474\,
            in1 => \N__5575\,
            in2 => \N__5456\,
            in3 => \N__5604\,
            lcout => \U712_CHIP_RAM.N_284\,
            ltout => \U712_CHIP_RAM.N_284_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__5663\,
            in1 => \N__5959\,
            in2 => \N__5478\,
            in3 => \N__6085\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__5475\,
            in1 => \N__5576\,
            in2 => \N__5457\,
            in3 => \N__6035\,
            lcout => \U712_CHIP_RAM.N_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__5424\,
            in1 => \N__5985\,
            in2 => \N__5415\,
            in3 => \N__5926\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9642\,
            ce => \N__6374\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_1_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__7755\,
            in1 => \N__6302\,
            in2 => \_gnd_net_\,
            in3 => \N__6747\,
            lcout => \U712_CHIP_RAM.N_218\,
            ltout => \U712_CHIP_RAM.N_218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQVN9G_2_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__6134\,
            in1 => \_gnd_net_\,
            in2 => \N__5418\,
            in3 => \N__5408\,
            lcout => \U712_CHIP_RAM.N_181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6291\,
            in2 => \_gnd_net_\,
            in3 => \N__5664\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_0_a2_0_a5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__5973\,
            in1 => \N__5927\,
            in2 => \N__5397\,
            in3 => \N__6086\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9642\,
            ce => \N__6374\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6650\,
            in1 => \N__7757\,
            in2 => \_gnd_net_\,
            in3 => \N__5667\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_i_a5_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6562\,
            in1 => \N__7280\,
            in2 => \N__5685\,
            in3 => \N__7246\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_257_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__6081\,
            in1 => \_gnd_net_\,
            in2 => \N__5682\,
            in3 => \N__5668\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIL1QU_2_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7758\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6649\,
            lcout => \U712_CHIP_RAM.N_338\,
            ltout => \U712_CHIP_RAM.N_338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__7245\,
            in1 => \N__6749\,
            in2 => \N__5673\,
            in3 => \N__6561\,
            lcout => \U712_CHIP_RAM.N_254\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5666\,
            in1 => \N__6028\,
            in2 => \_gnd_net_\,
            in3 => \N__6080\,
            lcout => \U712_CHIP_RAM.N_284_2\,
            ltout => \U712_CHIP_RAM.N_284_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__5598\,
            in1 => \N__5580\,
            in2 => \N__5553\,
            in3 => \N__5550\,
            lcout => \U712_CHIP_RAM.N_322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5735\,
            in1 => \N__5538\,
            in2 => \_gnd_net_\,
            in3 => \N__5528\,
            lcout => \U712_CHIP_RAM.N_256\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__5499\,
            in1 => \N__9328\,
            in2 => \N__9200\,
            in3 => \N__9471\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9340\,
            in1 => \N__9195\,
            in2 => \N__5493\,
            in3 => \N__10236\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5898\,
            in1 => \N__5880\,
            in2 => \_gnd_net_\,
            in3 => \N__9136\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9135\,
            in1 => \N__5862\,
            in2 => \_gnd_net_\,
            in3 => \N__5841\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6058\,
            in1 => \N__6261\,
            in2 => \_gnd_net_\,
            in3 => \N__6156\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9629\,
            ce => \N__5745\,
            sr => \N__10785\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__7444\,
            in1 => \N__5815\,
            in2 => \N__5787\,
            in3 => \N__7644\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_211_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10844\,
            in1 => \_gnd_net_\,
            in2 => \N__5763\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_211_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10842\,
            in2 => \_gnd_net_\,
            in3 => \N__5751\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_1_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7216\,
            in1 => \N__7122\,
            in2 => \_gnd_net_\,
            in3 => \N__6564\,
            lcout => \U712_CHIP_RAM.N_339\,
            ltout => \U712_CHIP_RAM.N_339_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101011111"
        )
    port map (
            in0 => \N__6740\,
            in1 => \N__7217\,
            in2 => \N__5739\,
            in3 => \N__6675\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000101"
        )
    port map (
            in0 => \N__6676\,
            in1 => \N__5730\,
            in2 => \N__5700\,
            in3 => \N__5696\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5988\,
            in3 => \N__10843\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6563\,
            in2 => \_gnd_net_\,
            in3 => \N__5979\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5928\,
            in1 => \N__7141\,
            in2 => \_gnd_net_\,
            in3 => \N__5976\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__9636\,
            ce => \N__6381\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6657\,
            in2 => \_gnd_net_\,
            in3 => \N__5967\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5929\,
            in1 => \N__7236\,
            in2 => \_gnd_net_\,
            in3 => \N__5964\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__9636\,
            ce => \N__6381\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5924\,
            in1 => \N__5960\,
            in2 => \_gnd_net_\,
            in3 => \N__5940\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__9636\,
            ce => \N__6381\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5930\,
            in1 => \N__6180\,
            in2 => \_gnd_net_\,
            in3 => \N__5937\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__9636\,
            ce => \N__6381\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5925\,
            in1 => \N__6201\,
            in2 => \_gnd_net_\,
            in3 => \N__5934\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__9636\,
            ce => \N__6381\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5931\,
            in1 => \N__6219\,
            in2 => \_gnd_net_\,
            in3 => \N__6384\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9636\,
            ce => \N__6381\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_1_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6231\,
            in1 => \N__10040\,
            in2 => \_gnd_net_\,
            in3 => \N__6357\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_289_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__6314\,
            in1 => \N__6267\,
            in2 => \N__6339\,
            in3 => \N__6336\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9639\,
            ce => 'H',
            sr => \N__10771\
        );

    \U712_CHIP_RAM.BANK0_RNO_2_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__6225\,
            in1 => \N__6303\,
            in2 => \N__6290\,
            in3 => \N__6748\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6036\,
            in1 => \N__6260\,
            in2 => \_gnd_net_\,
            in3 => \N__6133\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6633\,
            in1 => \N__7121\,
            in2 => \N__7237\,
            in3 => \N__6538\,
            lcout => \U712_CHIP_RAM.N_331\,
            ltout => \U712_CHIP_RAM.N_331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_7_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6218\,
            in1 => \N__6200\,
            in2 => \N__6183\,
            in3 => \N__6179\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER15\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_7_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6093\,
            in3 => \N__7753\,
            lcout => \U712_CHIP_RAM.N_337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011101100"
        )
    port map (
            in0 => \N__7754\,
            in1 => \N__6048\,
            in2 => \N__6483\,
            in3 => \N__7057\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9643\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7412\,
            in1 => \N__6656\,
            in2 => \N__6574\,
            in3 => \N__9321\,
            lcout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_a5_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6474\,
            in2 => \_gnd_net_\,
            in3 => \N__6467\,
            lcout => \U712_CHIP_RAM.un3_DMA_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6468\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7756\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9647\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__7777\,
            in1 => \N__10624\,
            in2 => \_gnd_net_\,
            in3 => \N__10530\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7518\,
            in1 => \N__6441\,
            in2 => \_gnd_net_\,
            in3 => \N__7524\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9618\,
            ce => \N__8080\,
            sr => \N__10798\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8266\,
            in1 => \N__9405\,
            in2 => \N__8236\,
            in3 => \N__6423\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9621\,
            ce => \N__8082\,
            sr => \N__10788\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__8226\,
            in1 => \N__8267\,
            in2 => \N__9507\,
            in3 => \N__6924\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9621\,
            ce => \N__8082\,
            sr => \N__10788\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000111"
        )
    port map (
            in0 => \N__9749\,
            in1 => \N__9128\,
            in2 => \N__8465\,
            in3 => \N__8390\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9294\,
            in1 => \N__9149\,
            in2 => \N__6933\,
            in3 => \N__9483\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9293\,
            in2 => \_gnd_net_\,
            in3 => \N__9129\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9175\,
            in1 => \N__6918\,
            in2 => \_gnd_net_\,
            in3 => \N__6906\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9346\,
            in1 => \N__9176\,
            in2 => \N__6891\,
            in3 => \N__9003\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9307\,
            in1 => \N__6888\,
            in2 => \N__9199\,
            in3 => \N__10209\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6882\,
            in1 => \N__9306\,
            in2 => \_gnd_net_\,
            in3 => \N__9492\,
            lcout => \U712_CHIP_RAM.N_146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_RNI8MQ3_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6865\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__7058\,
            in1 => \N__6753\,
            in2 => \N__6684\,
            in3 => \N__6702\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__6701\,
            in1 => \N__7421\,
            in2 => \N__6683\,
            in3 => \N__9314\,
            lcout => \U712_CHIP_RAM.CLK_EN_6_0_a5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7471\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7352\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__9359\,
            in1 => \N__7145\,
            in2 => \N__7068\,
            in3 => \N__7422\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9631\,
            ce => \N__7341\,
            sr => \N__10769\
        );

    \U712_BYTE_ENABLE.N_118_i_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__10629\,
            in1 => \N__6962\,
            in2 => \N__6954\,
            in3 => \N__9387\,
            lcout => \N_118_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_119_i_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__6942\,
            in1 => \N__6963\,
            in2 => \N__10545\,
            in3 => \N__9388\,
            lcout => \N_119_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7284\,
            in1 => \N__7235\,
            in2 => \N__7161\,
            in3 => \N__7074\,
            lcout => \U712_CHIP_RAM.N_287\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_a5_0_0_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7059\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6998\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_a5_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_0_a2_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8766\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8850\,
            lcout => \U712_BYTE_ENABLE.UUBE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_i_o5_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101001111"
        )
    port map (
            in0 => \N__8842\,
            in1 => \N__8732\,
            in2 => \N__8685\,
            in3 => \N__8605\,
            lcout => \U712_BYTE_ENABLE.N_216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7742\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_LDSn_i_0_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011111111"
        )
    port map (
            in0 => \N__8767\,
            in1 => \N__8579\,
            in2 => \N__8668\,
            in3 => \N__7838\,
            lcout => \N_163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8148\,
            in1 => \N__7563\,
            in2 => \N__9389\,
            in3 => \N__10428\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9619\,
            ce => \N__8073\,
            sr => \N__10813\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9751\,
            in2 => \_gnd_net_\,
            in3 => \N__8404\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011110000"
        )
    port map (
            in0 => \N__9371\,
            in1 => \N__8909\,
            in2 => \N__7527\,
            in3 => \N__9181\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011111111"
        )
    port map (
            in0 => \N__9370\,
            in1 => \N__8910\,
            in2 => \N__8230\,
            in3 => \N__9180\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__9204\,
            in1 => \N__8219\,
            in2 => \_gnd_net_\,
            in3 => \N__7512\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7479\,
            in2 => \N__7503\,
            in3 => \N__7992\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9623\,
            ce => \N__8085\,
            sr => \N__10802\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111010101"
        )
    port map (
            in0 => \N__8143\,
            in1 => \N__8016\,
            in2 => \N__9391\,
            in3 => \N__9528\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__9750\,
            in1 => \N__9173\,
            in2 => \_gnd_net_\,
            in3 => \N__8403\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => \U712_CHIP_RAM.CMA_5_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__9378\,
            in1 => \N__8015\,
            in2 => \N__7995\,
            in3 => \N__9527\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__10847\,
            in1 => \N__7986\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7980\,
            in1 => \N__7959\,
            in2 => \_gnd_net_\,
            in3 => \N__9174\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8268\,
            in1 => \N__7851\,
            in2 => \N__8241\,
            in3 => \N__7941\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9630\,
            ce => \N__8084\,
            sr => \N__10786\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__8234\,
            in1 => \N__8269\,
            in2 => \N__10131\,
            in3 => \N__7920\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9630\,
            ce => \N__8084\,
            sr => \N__10786\
        );

    \U712_CHIP_RAM.CLK_EN_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__7862\,
            in1 => \N__7893\,
            in2 => \_gnd_net_\,
            in3 => \N__7887\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9633\,
            ce => 'H',
            sr => \N__10774\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8943\,
            in1 => \N__8991\,
            in2 => \_gnd_net_\,
            in3 => \N__10050\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9858\,
            ce => \N__9817\,
            sr => \N__10772\
        );

    \U712_BYTE_ENABLE.un1_UDSn_i_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8768\,
            in2 => \_gnd_net_\,
            in3 => \N__7842\,
            lcout => \U712_BYTE_ENABLE_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WEn_LC_14_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8405\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9616\,
            ce => 'H',
            sr => \N__10821\
        );

    \U712_CHIP_RAM.CASn_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9203\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9617\,
            ce => 'H',
            sr => \N__10819\
        );

    \U712_CHIP_RAM.CRCSn_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8466\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9620\,
            ce => 'H',
            sr => \N__10818\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9365\,
            in1 => \N__8475\,
            in2 => \N__9201\,
            in3 => \N__10332\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8464\,
            in1 => \N__9194\,
            in2 => \N__9764\,
            in3 => \N__8406\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9624\,
            ce => \N__8081\,
            sr => \N__10814\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8283\,
            in1 => \N__9516\,
            in2 => \N__8235\,
            in3 => \N__8310\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9624\,
            ce => \N__8081\,
            sr => \N__10814\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__8282\,
            in1 => \N__9012\,
            in2 => \N__8237\,
            in3 => \N__9018\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9625\,
            ce => \N__8083\,
            sr => \N__10806\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8144\,
            in1 => \N__8127\,
            in2 => \N__9393\,
            in3 => \N__9867\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9625\,
            ce => \N__8083\,
            sr => \N__10806\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9390\,
            in1 => \N__9210\,
            in2 => \N__9202\,
            in3 => \N__10221\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10197\,
            in1 => \N__9967\,
            in2 => \_gnd_net_\,
            in3 => \N__10371\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9853\,
            ce => \N__9819\,
            sr => \N__10790\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8939\,
            in1 => \N__10044\,
            in2 => \_gnd_net_\,
            in3 => \N__9458\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9816\,
            sr => \N__10787\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8938\,
            in1 => \N__10043\,
            in2 => \_gnd_net_\,
            in3 => \N__8990\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9816\,
            sr => \N__10787\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9444\,
            in1 => \N__9993\,
            in2 => \_gnd_net_\,
            in3 => \N__8937\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9857\,
            ce => \N__9820\,
            sr => \N__10775\
        );

    \U712_BYTE_ENABLE.UUBE_i_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__8822\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8769\,
            lcout => \U712_BYTE_ENABLE_UUBE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_215_i_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101110000"
        )
    port map (
            in0 => \N__8847\,
            in1 => \N__8770\,
            in2 => \N__8682\,
            in3 => \N__8596\,
            lcout => \N_215_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_217_i_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111010000"
        )
    port map (
            in0 => \N__8849\,
            in1 => \N__8772\,
            in2 => \N__8684\,
            in3 => \N__8598\,
            lcout => \N_217_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_216_i_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010110000"
        )
    port map (
            in0 => \N__8848\,
            in1 => \N__8771\,
            in2 => \N__8683\,
            in3 => \N__8597\,
            lcout => \N_216_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RASn_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9765\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9622\,
            ce => 'H',
            sr => \N__10820\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10416\,
            in1 => \N__10039\,
            in2 => \_gnd_net_\,
            in3 => \N__10369\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9854\,
            ce => \N__9823\,
            sr => \N__10807\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10320\,
            in1 => \_gnd_net_\,
            in2 => \N__10049\,
            in3 => \N__10415\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9854\,
            ce => \N__9823\,
            sr => \N__10807\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10284\,
            in1 => \N__10035\,
            in2 => \_gnd_net_\,
            in3 => \N__10319\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9854\,
            ce => \N__9823\,
            sr => \N__10807\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10034\,
            in1 => \N__10196\,
            in2 => \_gnd_net_\,
            in3 => \N__10370\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__9822\,
            sr => \N__10803\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10313\,
            in1 => \N__10033\,
            in2 => \_gnd_net_\,
            in3 => \N__10408\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__9822\,
            sr => \N__10803\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9459\,
            in1 => \N__10032\,
            in2 => \_gnd_net_\,
            in3 => \N__10283\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__9822\,
            sr => \N__10803\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9457\,
            in1 => \N__10042\,
            in2 => \_gnd_net_\,
            in3 => \N__10275\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9855\,
            ce => \N__9818\,
            sr => \N__10791\
        );

    \U712_CHIP_RAM.DMA_A20_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__9992\,
            in1 => \N__10464\,
            in2 => \N__10118\,
            in3 => \N__10442\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10776\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10031\,
            in1 => \N__10119\,
            in2 => \_gnd_net_\,
            in3 => \N__10167\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9856\,
            ce => \N__9827\,
            sr => \N__10817\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__10414\,
            in1 => \_gnd_net_\,
            in2 => \N__10048\,
            in3 => \N__10362\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__9825\,
            sr => \N__10815\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10306\,
            in1 => \N__10027\,
            in2 => \_gnd_net_\,
            in3 => \N__10282\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__9825\,
            sr => \N__10815\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10165\,
            in1 => \N__10195\,
            in2 => \_gnd_net_\,
            in3 => \N__10026\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__9824\,
            sr => \N__10808\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9944\,
            in1 => \N__10114\,
            in2 => \_gnd_net_\,
            in3 => \N__10166\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__9821\,
            sr => \N__10804\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10194\,
            in1 => \N__10041\,
            in2 => \_gnd_net_\,
            in3 => \N__10164\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9852\,
            ce => \N__9826\,
            sr => \N__10816\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_22_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10093\,
            in1 => \N__10059\,
            in2 => \_gnd_net_\,
            in3 => \N__10011\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9851\,
            ce => \N__9828\,
            sr => \N__10822\
        );

    \U712_BUFFERS.un1_DRDENn_0_a5_LC_24_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__10674\,
            in1 => \N__10581\,
            in2 => \_gnd_net_\,
            in3 => \N__10499\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Sep 14 2025 20:46:27

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    DBRn : in std_logic;
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    PRnW : out std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    BLSn : out std_logic;
    TCIn : out std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__12997\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7443\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4611\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4602\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4395\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \DBRn_c_i_cascade_\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_10_6_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \C3_c\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \N_58_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_352\ : std_logic;
signal \INVU712_CYCLE_TERM.TACK_ENC_net\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_4\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_5\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_6\ : std_logic;
signal \PRnW_c\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\ : std_logic;
signal \BLSn_c\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STARTZ0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_36_0_cascade_\ : std_logic;
signal \TACK_OUT\ : std_logic;
signal \INVU712_CYCLE_TERM.TACK_STATE_0C_net\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.N_455_cascade_\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.N_387\ : std_logic;
signal \U712_REG_SM.N_185_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_7\ : std_logic;
signal \U712_REG_SM.N_368_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_378\ : std_logic;
signal \U712_REG_SM.N_441\ : std_logic;
signal \U712_REG_SM.N_358_cascade_\ : std_logic;
signal \U712_REG_SM.N_368\ : std_logic;
signal \U712_REG_SM.N_366\ : std_logic;
signal \U712_REG_SM.N_366_cascade_\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0\ : std_logic;
signal \CLK40_PLL\ : std_logic;
signal \CLK40_PLL_iso_i\ : std_logic;
signal \U712_REG_SM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_REG_SM.N_375\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_483\ : std_logic;
signal \U712_REG_SM.N_483_cascade_\ : std_logic;
signal \U712_REG_SM.N_367\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_358\ : std_logic;
signal \U712_REG_SM.N_592\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \U712_CYCLE_TERM.TACK_RST_0_i\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_407\ : std_logic;
signal \U712_REG_SM.N_369_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_4\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\ : std_logic;
signal \U712_REG_SM.N_481\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \U712_REG_SM.N_185\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_468\ : std_logic;
signal \N_65_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_343_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_466_cascade_\ : std_logic;
signal \N_67_i\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.N_185_0\ : std_logic;
signal \U712_REG_SM.N_482\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.N_362_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_493_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_503_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_596_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_596\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_i_i_a2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_365\ : std_logic;
signal \U712_CHIP_RAM.N_365_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_7\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1Z0Z_0_cascade_\ : std_logic;
signal \N_62_i\ : std_logic;
signal \U712_CHIP_RAM.N_452_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_2\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_cascade_\ : std_logic;
signal \U712_REG_SM.N_406\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_8\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_445_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_5_iv_0_0\ : std_logic;
signal \U712_BYTE_ENABLE.LMBE_0_i_o3_0_oZ0Z2\ : std_logic;
signal \N_282_i\ : std_logic;
signal \N_219\ : std_logic;
signal \N_60_i\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\ : std_logic;
signal \DBR_SYNC_i_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\ : std_logic;
signal \bfn_15_4_0_\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3\ : std_logic;
signal \U712_CHIP_RAM.N_451_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CAS_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_362\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_165_i_i_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_a2_1_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER19\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_344_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_435\ : std_logic;
signal \U712_CHIP_RAM.N_430\ : std_logic;
signal \U712_CHIP_RAM.N_347_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_590\ : std_logic;
signal \U712_CHIP_RAM.N_590_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_509_cascade_\ : std_logic;
signal \U712_CHIP_RAM.DBENn_8_0_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_CHIP_RAM.N_458_cascade_\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.N_350\ : std_logic;
signal \U712_CHIP_RAM.N_452\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a2_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_344\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_0\ : std_logic;
signal \U712_CHIP_RAM.N_72_cascade_\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CHIP_RAM.N_462\ : std_logic;
signal \U712_CHIP_RAM.N_503\ : std_logic;
signal \U712_CHIP_RAM.N_462_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_510\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\ : std_logic;
signal \N_119_i\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \N_61_i\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.N_431\ : std_logic;
signal \U712_CHIP_RAM.N_359\ : std_logic;
signal \U712_CHIP_RAM.N_595\ : std_logic;
signal \U712_CHIP_RAM.N_348\ : std_logic;
signal \U712_CHIP_RAM.N_595_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_577\ : std_logic;
signal \U712_CHIP_RAM.N_279\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_i_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0\ : std_logic;
signal \bfn_16_6_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.N_132_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_436\ : std_logic;
signal \U712_CHIP_RAM.N_499\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_506_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_147_i_i_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_147_i_i_a2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_500_i\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto7_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_CHIP_RAM.N_509\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_508\ : std_logic;
signal \U712_CHIP_RAM.N_494\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \N_207_i\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \RASn_c\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_354_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_9\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.N_354\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA25_0_i_0\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_2\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \RnW_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \DMA_WRITE_CYCLE\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \N_409\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \PRnW_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \BLSn_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    TCIn <= \TCIn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    PRnW <= \PRnW_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    \C3_wire\ <= C3;
    BLSn <= \BLSn_wire\;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL\,
            REFERENCECLK => \N__4413\,
            RESETB => \N__7416\,
            BYPASS => \GNDG0\,
            PLLOUTCOREA => OPEN,
            SDI => \GNDG0\,
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => \GNDG0\,
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => \GNDG0\
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12997\,
            DIN => \N__12996\,
            DOUT => \N__12995\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12997\,
            PADOUT => \N__12996\,
            PADIN => \N__12995\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6363\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12988\,
            DIN => \N__12987\,
            DOUT => \N__12986\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12988\,
            PADOUT => \N__12987\,
            PADIN => \N__12986\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12979\,
            DIN => \N__12978\,
            DOUT => \N__12977\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12979\,
            PADOUT => \N__12978\,
            PADIN => \N__12977\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9399\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12970\,
            DIN => \N__12969\,
            DOUT => \N__12968\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12970\,
            PADOUT => \N__12969\,
            PADIN => \N__12968\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10707\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12961\,
            DIN => \N__12960\,
            DOUT => \N__12959\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12961\,
            PADOUT => \N__12960\,
            PADIN => \N__12959\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12952\,
            DIN => \N__12951\,
            DOUT => \N__12950\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12952\,
            PADOUT => \N__12951\,
            PADIN => \N__12950\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12943\,
            DIN => \N__12942\,
            DOUT => \N__12941\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12943\,
            PADOUT => \N__12942\,
            PADIN => \N__12941\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12934\,
            DIN => \N__12933\,
            DOUT => \N__12932\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12934\,
            PADOUT => \N__12933\,
            PADIN => \N__12932\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12925\,
            DIN => \N__12924\,
            DOUT => \N__12923\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12925\,
            PADOUT => \N__12924\,
            PADIN => \N__12923\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12916\,
            DIN => \N__12915\,
            DOUT => \N__12914\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12916\,
            PADOUT => \N__12915\,
            PADIN => \N__12914\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12907\,
            DIN => \N__12906\,
            DOUT => \N__12905\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12907\,
            PADOUT => \N__12906\,
            PADIN => \N__12905\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12898\,
            DIN => \N__12897\,
            DOUT => \N__12896\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12898\,
            PADOUT => \N__12897\,
            PADIN => \N__12896\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6033\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12889\,
            DIN => \N__12888\,
            DOUT => \N__12887\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12889\,
            PADOUT => \N__12888\,
            PADIN => \N__12887\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6465\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12880\,
            DIN => \N__12879\,
            DOUT => \N__12878\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12880\,
            PADOUT => \N__12879\,
            PADIN => \N__12878\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12871\,
            DIN => \N__12870\,
            DOUT => \N__12869\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12871\,
            PADOUT => \N__12870\,
            PADIN => \N__12869\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6968\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12862\,
            DIN => \N__12861\,
            DOUT => \N__12860\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12862\,
            PADOUT => \N__12861\,
            PADIN => \N__12860\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12853\,
            DIN => \N__12852\,
            DOUT => \N__12851\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12853\,
            PADOUT => \N__12852\,
            PADIN => \N__12851\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12844\,
            DIN => \N__12843\,
            DOUT => \N__12842\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12844\,
            PADOUT => \N__12843\,
            PADIN => \N__12842\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4989\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12835\,
            DIN => \N__12834\,
            DOUT => \N__12833\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12835\,
            PADOUT => \N__12834\,
            PADIN => \N__12833\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12826\,
            DIN => \N__12825\,
            DOUT => \N__12824\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12826\,
            PADOUT => \N__12825\,
            PADIN => \N__12824\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12817\,
            DIN => \N__12816\,
            DOUT => \N__12815\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12817\,
            PADOUT => \N__12816\,
            PADIN => \N__12815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9222\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12808\,
            DIN => \N__12807\,
            DOUT => \N__12806\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12808\,
            PADOUT => \N__12807\,
            PADIN => \N__12806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12799\,
            DIN => \N__12798\,
            DOUT => \N__12797\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12799\,
            PADOUT => \N__12798\,
            PADIN => \N__12797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9417\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12790\,
            DIN => \N__12789\,
            DOUT => \N__12788\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12790\,
            PADOUT => \N__12789\,
            PADIN => \N__12788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12781\,
            DIN => \N__12780\,
            DOUT => \N__12779\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12781\,
            PADOUT => \N__12780\,
            PADIN => \N__12779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6480\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12772\,
            DIN => \N__12771\,
            DOUT => \N__12770\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12772\,
            PADOUT => \N__12771\,
            PADIN => \N__12770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5257\,
            DIN0 => OPEN,
            DOUT0 => \N__4894\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12763\,
            DIN => \N__12762\,
            DOUT => \N__12761\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12763\,
            PADOUT => \N__12762\,
            PADIN => \N__12761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12754\,
            DIN => \N__12753\,
            DOUT => \N__12752\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12754\,
            PADOUT => \N__12753\,
            PADIN => \N__12752\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12745\,
            DIN => \N__12744\,
            DOUT => \N__12743\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12745\,
            PADOUT => \N__12744\,
            PADIN => \N__12743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12736\,
            DIN => \N__12735\,
            DOUT => \N__12734\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12736\,
            PADOUT => \N__12735\,
            PADIN => \N__12734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12727\,
            DIN => \N__12726\,
            DOUT => \N__12725\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12727\,
            PADOUT => \N__12726\,
            PADIN => \N__12725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12718\,
            DIN => \N__12717\,
            DOUT => \N__12716\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12718\,
            PADOUT => \N__12717\,
            PADIN => \N__12716\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6501\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12709\,
            DIN => \N__12708\,
            DOUT => \N__12707\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12709\,
            PADOUT => \N__12708\,
            PADIN => \N__12707\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12700\,
            DIN => \N__12699\,
            DOUT => \N__12698\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12700\,
            PADOUT => \N__12699\,
            PADIN => \N__12698\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12691\,
            DIN => \N__12690\,
            DOUT => \N__12689\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12691\,
            PADOUT => \N__12690\,
            PADIN => \N__12689\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12682\,
            DIN => \N__12681\,
            DOUT => \N__12680\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12682\,
            PADOUT => \N__12681\,
            PADIN => \N__12680\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12673\,
            DIN => \N__12672\,
            DOUT => \N__12671\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12673\,
            PADOUT => \N__12672\,
            PADIN => \N__12671\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12664\,
            DIN => \N__12663\,
            DOUT => \N__12662\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12664\,
            PADOUT => \N__12663\,
            PADIN => \N__12662\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9432\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12655\,
            DIN => \N__12654\,
            DOUT => \N__12653\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12655\,
            PADOUT => \N__12654\,
            PADIN => \N__12653\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12646\,
            DIN => \N__12645\,
            DOUT => \N__12644\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12646\,
            PADOUT => \N__12645\,
            PADIN => \N__12644\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12637\,
            DIN => \N__12636\,
            DOUT => \N__12635\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12637\,
            PADOUT => \N__12636\,
            PADIN => \N__12635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5817\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12628\,
            DIN => \N__12627\,
            DOUT => \N__12626\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12628\,
            PADOUT => \N__12627\,
            PADIN => \N__12626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7296\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12619\,
            DIN => \N__12618\,
            DOUT => \N__12617\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12619\,
            PADOUT => \N__12618\,
            PADIN => \N__12617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12610\,
            DIN => \N__12609\,
            DOUT => \N__12608\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12610\,
            PADOUT => \N__12609\,
            PADIN => \N__12608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9924\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12601\,
            DIN => \N__12600\,
            DOUT => \N__12599\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12601\,
            PADOUT => \N__12600\,
            PADIN => \N__12599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10134\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12592\,
            DIN => \N__12591\,
            DOUT => \N__12590\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12592\,
            PADOUT => \N__12591\,
            PADIN => \N__12590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4761\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12583\,
            DIN => \N__12582\,
            DOUT => \N__12581\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12583\,
            PADOUT => \N__12582\,
            PADIN => \N__12581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12574\,
            DIN => \N__12573\,
            DOUT => \N__12572\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12574\,
            PADOUT => \N__12573\,
            PADIN => \N__12572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12565\,
            DIN => \N__12564\,
            DOUT => \N__12563\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12565\,
            PADOUT => \N__12564\,
            PADIN => \N__12563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6303\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12556\,
            DIN => \N__12555\,
            DOUT => \N__12554\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12556\,
            PADOUT => \N__12555\,
            PADIN => \N__12554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5262\,
            DIN0 => OPEN,
            DOUT0 => \N__4901\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12547\,
            DIN => \N__12546\,
            DOUT => \N__12545\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12547\,
            PADOUT => \N__12546\,
            PADIN => \N__12545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10572\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12538\,
            DIN => \N__12537\,
            DOUT => \N__12536\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12538\,
            PADOUT => \N__12537\,
            PADIN => \N__12536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4638\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12529\,
            DIN => \N__12528\,
            DOUT => \N__12527\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12529\,
            PADOUT => \N__12528\,
            PADIN => \N__12527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5886\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12520\,
            DIN => \N__12519\,
            DOUT => \N__12518\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12520\,
            PADOUT => \N__12519\,
            PADIN => \N__12518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12511\,
            DIN => \N__12510\,
            DOUT => \N__12509\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12511\,
            PADOUT => \N__12510\,
            PADIN => \N__12509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12502\,
            DIN => \N__12501\,
            DOUT => \N__12500\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12502\,
            PADOUT => \N__12501\,
            PADIN => \N__12500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7359\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12493\,
            DIN => \N__12492\,
            DOUT => \N__12491\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12493\,
            PADOUT => \N__12492\,
            PADIN => \N__12491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12484\,
            DIN => \N__12483\,
            DOUT => \N__12482\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12484\,
            PADOUT => \N__12483\,
            PADIN => \N__12482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12475\,
            DIN => \N__12474\,
            DOUT => \N__12473\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12475\,
            PADOUT => \N__12474\,
            PADIN => \N__12473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5097\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12466\,
            DIN => \N__12465\,
            DOUT => \N__12464\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12466\,
            PADOUT => \N__12465\,
            PADIN => \N__12464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7467\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12457\,
            DIN => \N__12456\,
            DOUT => \N__12455\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12457\,
            PADOUT => \N__12456\,
            PADIN => \N__12455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12448\,
            DIN => \N__12447\,
            DOUT => \N__12446\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12448\,
            PADOUT => \N__12447\,
            PADIN => \N__12446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5832\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12439\,
            DIN => \N__12438\,
            DOUT => \N__12437\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12439\,
            PADOUT => \N__12438\,
            PADIN => \N__12437\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5261\,
            DIN0 => OPEN,
            DOUT0 => \N__4902\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12430\,
            DIN => \N__12429\,
            DOUT => \N__12428\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12430\,
            PADOUT => \N__12429\,
            PADIN => \N__12428\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7455\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12421\,
            DIN => \N__12420\,
            DOUT => \N__12419\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12421\,
            PADOUT => \N__12420\,
            PADIN => \N__12419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12412\,
            DIN => \N__12411\,
            DOUT => \N__12410\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12412\,
            PADOUT => \N__12411\,
            PADIN => \N__12410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12403\,
            DIN => \N__12402\,
            DOUT => \N__12401\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12403\,
            PADOUT => \N__12402\,
            PADIN => \N__12401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6006\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12394\,
            DIN => \N__12393\,
            DOUT => \N__12392\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12394\,
            PADOUT => \N__12393\,
            PADIN => \N__12392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12385\,
            DIN => \N__12384\,
            DOUT => \N__12383\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12385\,
            PADOUT => \N__12384\,
            PADIN => \N__12383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12376\,
            DIN => \N__12375\,
            DOUT => \N__12374\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12376\,
            PADOUT => \N__12375\,
            PADIN => \N__12374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5049\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12367\,
            DIN => \N__12366\,
            DOUT => \N__12365\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12367\,
            PADOUT => \N__12366\,
            PADIN => \N__12365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12358\,
            DIN => \N__12357\,
            DOUT => \N__12356\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12358\,
            PADOUT => \N__12357\,
            PADIN => \N__12356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12349\,
            DIN => \N__12348\,
            DOUT => \N__12347\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12349\,
            PADOUT => \N__12348\,
            PADIN => \N__12347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9660\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12340\,
            DIN => \N__12339\,
            DOUT => \N__12338\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12340\,
            PADOUT => \N__12339\,
            PADIN => \N__12338\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5934\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12331\,
            DIN => \N__12330\,
            DOUT => \N__12329\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12331\,
            PADOUT => \N__12330\,
            PADIN => \N__12329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7839\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12322\,
            DIN => \N__12321\,
            DOUT => \N__12320\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12322\,
            PADOUT => \N__12321\,
            PADIN => \N__12320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6912\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12313\,
            DIN => \N__12312\,
            DOUT => \N__12311\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12313\,
            PADOUT => \N__12312\,
            PADIN => \N__12311\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12304\,
            DIN => \N__12303\,
            DOUT => \N__12302\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12304\,
            PADOUT => \N__12303\,
            PADIN => \N__12302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12295\,
            DIN => \N__12294\,
            DOUT => \N__12293\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12295\,
            PADOUT => \N__12294\,
            PADIN => \N__12293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6063\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12286\,
            DIN => \N__12285\,
            DOUT => \N__12284\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12286\,
            PADOUT => \N__12285\,
            PADIN => \N__12284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12277\,
            DIN => \N__12276\,
            DOUT => \N__12275\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12277\,
            PADOUT => \N__12276\,
            PADIN => \N__12275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12268\,
            DIN => \N__12267\,
            DOUT => \N__12266\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12268\,
            PADOUT => \N__12267\,
            PADIN => \N__12266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7893\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12259\,
            DIN => \N__12258\,
            DOUT => \N__12257\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12259\,
            PADOUT => \N__12258\,
            PADIN => \N__12257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5973\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12250\,
            DIN => \N__12249\,
            DOUT => \N__12248\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12250\,
            PADOUT => \N__12249\,
            PADIN => \N__12248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5505\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PRnW_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12241\,
            DIN => \N__12240\,
            DOUT => \N__12239\,
            PACKAGEPIN => \PRnW_wire\
        );

    \PRnW_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12241\,
            PADOUT => \N__12240\,
            PADIN => \N__12239\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4797\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12232\,
            DIN => \N__12231\,
            DOUT => \N__12230\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12232\,
            PADOUT => \N__12231\,
            PADIN => \N__12230\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12223\,
            DIN => \N__12222\,
            DOUT => \N__12221\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12223\,
            PADOUT => \N__12222\,
            PADIN => \N__12221\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5504\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12214\,
            DIN => \N__12213\,
            DOUT => \N__12212\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12214\,
            PADOUT => \N__12213\,
            PADIN => \N__12212\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4452\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12205\,
            DIN => \N__12204\,
            DOUT => \N__12203\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12205\,
            PADOUT => \N__12204\,
            PADIN => \N__12203\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9633\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12196\,
            DIN => \N__12195\,
            DOUT => \N__12194\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12196\,
            PADOUT => \N__12195\,
            PADIN => \N__12194\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12187\,
            DIN => \N__12186\,
            DOUT => \N__12185\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12187\,
            PADOUT => \N__12186\,
            PADIN => \N__12185\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12178\,
            DIN => \N__12177\,
            DOUT => \N__12176\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12178\,
            PADOUT => \N__12177\,
            PADIN => \N__12176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BLSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12169\,
            DIN => \N__12168\,
            DOUT => \N__12167\,
            PACKAGEPIN => \BLSn_wire\
        );

    \BLSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12169\,
            PADOUT => \N__12168\,
            PADIN => \N__12167\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4760\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12160\,
            DIN => \N__12159\,
            DOUT => \N__12158\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12160\,
            PADOUT => \N__12159\,
            PADIN => \N__12158\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12151\,
            DIN => \N__12150\,
            DOUT => \N__12149\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12151\,
            PADOUT => \N__12150\,
            PADIN => \N__12149\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5479\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12142\,
            DIN => \N__12141\,
            DOUT => \N__12140\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12142\,
            PADOUT => \N__12141\,
            PADIN => \N__12140\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9336\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12133\,
            DIN => \N__12132\,
            DOUT => \N__12131\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12133\,
            PADOUT => \N__12132\,
            PADIN => \N__12131\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4719\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12124\,
            DIN => \N__12123\,
            DOUT => \N__12122\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12124\,
            PADOUT => \N__12123\,
            PADIN => \N__12122\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10323\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2950\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12099\
        );

    \I__2949\ : InMux
    port map (
            O => \N__12104\,
            I => \N__12096\
        );

    \I__2948\ : InMux
    port map (
            O => \N__12103\,
            I => \N__12091\
        );

    \I__2947\ : InMux
    port map (
            O => \N__12102\,
            I => \N__12091\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__12099\,
            I => \N__12088\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__12096\,
            I => \N__12083\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__12091\,
            I => \N__12083\
        );

    \I__2943\ : Span4Mux_v
    port map (
            O => \N__12088\,
            I => \N__12078\
        );

    \I__2942\ : Span4Mux_v
    port map (
            O => \N__12083\,
            I => \N__12078\
        );

    \I__2941\ : Span4Mux_v
    port map (
            O => \N__12078\,
            I => \N__12075\
        );

    \I__2940\ : Sp12to4
    port map (
            O => \N__12075\,
            I => \N__12072\
        );

    \I__2939\ : Odrv12
    port map (
            O => \N__12072\,
            I => \DRA_c_4\
        );

    \I__2938\ : InMux
    port map (
            O => \N__12069\,
            I => \N__12066\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__12066\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2936\ : InMux
    port map (
            O => \N__12063\,
            I => \N__12060\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__12060\,
            I => \N__12057\
        );

    \I__2934\ : Span4Mux_h
    port map (
            O => \N__12057\,
            I => \N__12054\
        );

    \I__2933\ : Odrv4
    port map (
            O => \N__12054\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2932\ : InMux
    port map (
            O => \N__12051\,
            I => \N__12048\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__12048\,
            I => \N__12045\
        );

    \I__2930\ : Odrv12
    port map (
            O => \N__12045\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\
        );

    \I__2929\ : InMux
    port map (
            O => \N__12042\,
            I => \N__12039\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__12039\,
            I => \N__12036\
        );

    \I__2927\ : Span4Mux_v
    port map (
            O => \N__12036\,
            I => \N__12032\
        );

    \I__2926\ : InMux
    port map (
            O => \N__12035\,
            I => \N__12029\
        );

    \I__2925\ : Span4Mux_h
    port map (
            O => \N__12032\,
            I => \N__12026\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__12029\,
            I => \N__12023\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__12026\,
            I => \RAS0n_c\
        );

    \I__2922\ : Odrv12
    port map (
            O => \N__12023\,
            I => \RAS0n_c\
        );

    \I__2921\ : InMux
    port map (
            O => \N__12018\,
            I => \N__12015\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__12015\,
            I => \N__12012\
        );

    \I__2919\ : Span12Mux_v
    port map (
            O => \N__12012\,
            I => \N__12009\
        );

    \I__2918\ : Odrv12
    port map (
            O => \N__12009\,
            I => \RAS1n_c\
        );

    \I__2917\ : CascadeMux
    port map (
            O => \N__12006\,
            I => \N__11996\
        );

    \I__2916\ : InMux
    port map (
            O => \N__12005\,
            I => \N__11977\
        );

    \I__2915\ : InMux
    port map (
            O => \N__12004\,
            I => \N__11977\
        );

    \I__2914\ : InMux
    port map (
            O => \N__12003\,
            I => \N__11977\
        );

    \I__2913\ : InMux
    port map (
            O => \N__12002\,
            I => \N__11977\
        );

    \I__2912\ : InMux
    port map (
            O => \N__12001\,
            I => \N__11970\
        );

    \I__2911\ : InMux
    port map (
            O => \N__12000\,
            I => \N__11965\
        );

    \I__2910\ : InMux
    port map (
            O => \N__11999\,
            I => \N__11965\
        );

    \I__2909\ : InMux
    port map (
            O => \N__11996\,
            I => \N__11960\
        );

    \I__2908\ : InMux
    port map (
            O => \N__11995\,
            I => \N__11960\
        );

    \I__2907\ : InMux
    port map (
            O => \N__11994\,
            I => \N__11953\
        );

    \I__2906\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11953\
        );

    \I__2905\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11953\
        );

    \I__2904\ : InMux
    port map (
            O => \N__11991\,
            I => \N__11950\
        );

    \I__2903\ : InMux
    port map (
            O => \N__11990\,
            I => \N__11943\
        );

    \I__2902\ : InMux
    port map (
            O => \N__11989\,
            I => \N__11943\
        );

    \I__2901\ : InMux
    port map (
            O => \N__11988\,
            I => \N__11943\
        );

    \I__2900\ : InMux
    port map (
            O => \N__11987\,
            I => \N__11938\
        );

    \I__2899\ : InMux
    port map (
            O => \N__11986\,
            I => \N__11938\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__11977\,
            I => \N__11935\
        );

    \I__2897\ : InMux
    port map (
            O => \N__11976\,
            I => \N__11932\
        );

    \I__2896\ : InMux
    port map (
            O => \N__11975\,
            I => \N__11927\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__11974\,
            I => \N__11916\
        );

    \I__2894\ : CascadeMux
    port map (
            O => \N__11973\,
            I => \N__11913\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__11970\,
            I => \N__11906\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__11965\,
            I => \N__11906\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__11960\,
            I => \N__11903\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__11953\,
            I => \N__11894\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__11950\,
            I => \N__11894\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__11943\,
            I => \N__11894\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__11938\,
            I => \N__11894\
        );

    \I__2886\ : Span4Mux_v
    port map (
            O => \N__11935\,
            I => \N__11889\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__11932\,
            I => \N__11889\
        );

    \I__2884\ : InMux
    port map (
            O => \N__11931\,
            I => \N__11886\
        );

    \I__2883\ : InMux
    port map (
            O => \N__11930\,
            I => \N__11883\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__11927\,
            I => \N__11880\
        );

    \I__2881\ : InMux
    port map (
            O => \N__11926\,
            I => \N__11873\
        );

    \I__2880\ : InMux
    port map (
            O => \N__11925\,
            I => \N__11873\
        );

    \I__2879\ : InMux
    port map (
            O => \N__11924\,
            I => \N__11873\
        );

    \I__2878\ : InMux
    port map (
            O => \N__11923\,
            I => \N__11870\
        );

    \I__2877\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11865\
        );

    \I__2876\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11865\
        );

    \I__2875\ : InMux
    port map (
            O => \N__11920\,
            I => \N__11862\
        );

    \I__2874\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11853\
        );

    \I__2873\ : InMux
    port map (
            O => \N__11916\,
            I => \N__11853\
        );

    \I__2872\ : InMux
    port map (
            O => \N__11913\,
            I => \N__11853\
        );

    \I__2871\ : InMux
    port map (
            O => \N__11912\,
            I => \N__11853\
        );

    \I__2870\ : InMux
    port map (
            O => \N__11911\,
            I => \N__11850\
        );

    \I__2869\ : Span4Mux_v
    port map (
            O => \N__11906\,
            I => \N__11847\
        );

    \I__2868\ : Span4Mux_v
    port map (
            O => \N__11903\,
            I => \N__11835\
        );

    \I__2867\ : Span4Mux_v
    port map (
            O => \N__11894\,
            I => \N__11835\
        );

    \I__2866\ : Span4Mux_h
    port map (
            O => \N__11889\,
            I => \N__11835\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__11886\,
            I => \N__11835\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__11883\,
            I => \N__11835\
        );

    \I__2863\ : Span12Mux_v
    port map (
            O => \N__11880\,
            I => \N__11829\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__11873\,
            I => \N__11820\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__11870\,
            I => \N__11820\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__11865\,
            I => \N__11820\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__11862\,
            I => \N__11820\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__11853\,
            I => \N__11815\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__11850\,
            I => \N__11815\
        );

    \I__2856\ : Span4Mux_v
    port map (
            O => \N__11847\,
            I => \N__11812\
        );

    \I__2855\ : InMux
    port map (
            O => \N__11846\,
            I => \N__11809\
        );

    \I__2854\ : Span4Mux_v
    port map (
            O => \N__11835\,
            I => \N__11806\
        );

    \I__2853\ : InMux
    port map (
            O => \N__11834\,
            I => \N__11803\
        );

    \I__2852\ : InMux
    port map (
            O => \N__11833\,
            I => \N__11798\
        );

    \I__2851\ : InMux
    port map (
            O => \N__11832\,
            I => \N__11798\
        );

    \I__2850\ : Span12Mux_h
    port map (
            O => \N__11829\,
            I => \N__11795\
        );

    \I__2849\ : Span12Mux_v
    port map (
            O => \N__11820\,
            I => \N__11792\
        );

    \I__2848\ : Span12Mux_v
    port map (
            O => \N__11815\,
            I => \N__11789\
        );

    \I__2847\ : Sp12to4
    port map (
            O => \N__11812\,
            I => \N__11784\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__11809\,
            I => \N__11784\
        );

    \I__2845\ : Span4Mux_h
    port map (
            O => \N__11806\,
            I => \N__11781\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__11803\,
            I => \N__11776\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__11798\,
            I => \N__11776\
        );

    \I__2842\ : Span12Mux_v
    port map (
            O => \N__11795\,
            I => \N__11771\
        );

    \I__2841\ : Span12Mux_h
    port map (
            O => \N__11792\,
            I => \N__11771\
        );

    \I__2840\ : Span12Mux_h
    port map (
            O => \N__11789\,
            I => \N__11768\
        );

    \I__2839\ : Span12Mux_h
    port map (
            O => \N__11784\,
            I => \N__11761\
        );

    \I__2838\ : Sp12to4
    port map (
            O => \N__11781\,
            I => \N__11761\
        );

    \I__2837\ : Span12Mux_v
    port map (
            O => \N__11776\,
            I => \N__11761\
        );

    \I__2836\ : Odrv12
    port map (
            O => \N__11771\,
            I => \RESETn_c\
        );

    \I__2835\ : Odrv12
    port map (
            O => \N__11768\,
            I => \RESETn_c\
        );

    \I__2834\ : Odrv12
    port map (
            O => \N__11761\,
            I => \RESETn_c\
        );

    \I__2833\ : InMux
    port map (
            O => \N__11754\,
            I => \N__11751\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__11751\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2831\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11745\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__11745\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__2829\ : InMux
    port map (
            O => \N__11742\,
            I => \N__11739\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__11739\,
            I => \N__11690\
        );

    \I__2827\ : ClkMux
    port map (
            O => \N__11738\,
            I => \N__11592\
        );

    \I__2826\ : ClkMux
    port map (
            O => \N__11737\,
            I => \N__11592\
        );

    \I__2825\ : ClkMux
    port map (
            O => \N__11736\,
            I => \N__11592\
        );

    \I__2824\ : ClkMux
    port map (
            O => \N__11735\,
            I => \N__11592\
        );

    \I__2823\ : ClkMux
    port map (
            O => \N__11734\,
            I => \N__11592\
        );

    \I__2822\ : ClkMux
    port map (
            O => \N__11733\,
            I => \N__11592\
        );

    \I__2821\ : ClkMux
    port map (
            O => \N__11732\,
            I => \N__11592\
        );

    \I__2820\ : ClkMux
    port map (
            O => \N__11731\,
            I => \N__11592\
        );

    \I__2819\ : ClkMux
    port map (
            O => \N__11730\,
            I => \N__11592\
        );

    \I__2818\ : ClkMux
    port map (
            O => \N__11729\,
            I => \N__11592\
        );

    \I__2817\ : ClkMux
    port map (
            O => \N__11728\,
            I => \N__11592\
        );

    \I__2816\ : ClkMux
    port map (
            O => \N__11727\,
            I => \N__11592\
        );

    \I__2815\ : ClkMux
    port map (
            O => \N__11726\,
            I => \N__11592\
        );

    \I__2814\ : ClkMux
    port map (
            O => \N__11725\,
            I => \N__11592\
        );

    \I__2813\ : ClkMux
    port map (
            O => \N__11724\,
            I => \N__11592\
        );

    \I__2812\ : ClkMux
    port map (
            O => \N__11723\,
            I => \N__11592\
        );

    \I__2811\ : ClkMux
    port map (
            O => \N__11722\,
            I => \N__11592\
        );

    \I__2810\ : ClkMux
    port map (
            O => \N__11721\,
            I => \N__11592\
        );

    \I__2809\ : ClkMux
    port map (
            O => \N__11720\,
            I => \N__11592\
        );

    \I__2808\ : ClkMux
    port map (
            O => \N__11719\,
            I => \N__11592\
        );

    \I__2807\ : ClkMux
    port map (
            O => \N__11718\,
            I => \N__11592\
        );

    \I__2806\ : ClkMux
    port map (
            O => \N__11717\,
            I => \N__11592\
        );

    \I__2805\ : ClkMux
    port map (
            O => \N__11716\,
            I => \N__11592\
        );

    \I__2804\ : ClkMux
    port map (
            O => \N__11715\,
            I => \N__11592\
        );

    \I__2803\ : ClkMux
    port map (
            O => \N__11714\,
            I => \N__11592\
        );

    \I__2802\ : ClkMux
    port map (
            O => \N__11713\,
            I => \N__11592\
        );

    \I__2801\ : ClkMux
    port map (
            O => \N__11712\,
            I => \N__11592\
        );

    \I__2800\ : ClkMux
    port map (
            O => \N__11711\,
            I => \N__11592\
        );

    \I__2799\ : ClkMux
    port map (
            O => \N__11710\,
            I => \N__11592\
        );

    \I__2798\ : ClkMux
    port map (
            O => \N__11709\,
            I => \N__11592\
        );

    \I__2797\ : ClkMux
    port map (
            O => \N__11708\,
            I => \N__11592\
        );

    \I__2796\ : ClkMux
    port map (
            O => \N__11707\,
            I => \N__11592\
        );

    \I__2795\ : ClkMux
    port map (
            O => \N__11706\,
            I => \N__11592\
        );

    \I__2794\ : ClkMux
    port map (
            O => \N__11705\,
            I => \N__11592\
        );

    \I__2793\ : ClkMux
    port map (
            O => \N__11704\,
            I => \N__11592\
        );

    \I__2792\ : ClkMux
    port map (
            O => \N__11703\,
            I => \N__11592\
        );

    \I__2791\ : ClkMux
    port map (
            O => \N__11702\,
            I => \N__11592\
        );

    \I__2790\ : ClkMux
    port map (
            O => \N__11701\,
            I => \N__11592\
        );

    \I__2789\ : ClkMux
    port map (
            O => \N__11700\,
            I => \N__11592\
        );

    \I__2788\ : ClkMux
    port map (
            O => \N__11699\,
            I => \N__11592\
        );

    \I__2787\ : ClkMux
    port map (
            O => \N__11698\,
            I => \N__11592\
        );

    \I__2786\ : ClkMux
    port map (
            O => \N__11697\,
            I => \N__11592\
        );

    \I__2785\ : ClkMux
    port map (
            O => \N__11696\,
            I => \N__11592\
        );

    \I__2784\ : ClkMux
    port map (
            O => \N__11695\,
            I => \N__11592\
        );

    \I__2783\ : ClkMux
    port map (
            O => \N__11694\,
            I => \N__11592\
        );

    \I__2782\ : ClkMux
    port map (
            O => \N__11693\,
            I => \N__11592\
        );

    \I__2781\ : Glb2LocalMux
    port map (
            O => \N__11690\,
            I => \N__11592\
        );

    \I__2780\ : ClkMux
    port map (
            O => \N__11689\,
            I => \N__11592\
        );

    \I__2779\ : GlobalMux
    port map (
            O => \N__11592\,
            I => \CLK80_PLL\
        );

    \I__2778\ : InMux
    port map (
            O => \N__11589\,
            I => \N__11586\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__11586\,
            I => \N__11580\
        );

    \I__2776\ : InMux
    port map (
            O => \N__11585\,
            I => \N__11577\
        );

    \I__2775\ : InMux
    port map (
            O => \N__11584\,
            I => \N__11572\
        );

    \I__2774\ : InMux
    port map (
            O => \N__11583\,
            I => \N__11572\
        );

    \I__2773\ : Span4Mux_v
    port map (
            O => \N__11580\,
            I => \N__11569\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__11577\,
            I => \N__11564\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__11572\,
            I => \N__11564\
        );

    \I__2770\ : Span4Mux_v
    port map (
            O => \N__11569\,
            I => \N__11561\
        );

    \I__2769\ : Span12Mux_v
    port map (
            O => \N__11564\,
            I => \N__11558\
        );

    \I__2768\ : Span4Mux_h
    port map (
            O => \N__11561\,
            I => \N__11555\
        );

    \I__2767\ : Odrv12
    port map (
            O => \N__11558\,
            I => \DRA_c_3\
        );

    \I__2766\ : Odrv4
    port map (
            O => \N__11555\,
            I => \DRA_c_3\
        );

    \I__2765\ : InMux
    port map (
            O => \N__11550\,
            I => \N__11547\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__11547\,
            I => \N__11544\
        );

    \I__2763\ : Span4Mux_v
    port map (
            O => \N__11544\,
            I => \N__11538\
        );

    \I__2762\ : InMux
    port map (
            O => \N__11543\,
            I => \N__11535\
        );

    \I__2761\ : InMux
    port map (
            O => \N__11542\,
            I => \N__11530\
        );

    \I__2760\ : InMux
    port map (
            O => \N__11541\,
            I => \N__11530\
        );

    \I__2759\ : Span4Mux_v
    port map (
            O => \N__11538\,
            I => \N__11527\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__11535\,
            I => \N__11522\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__11530\,
            I => \N__11522\
        );

    \I__2756\ : Span4Mux_h
    port map (
            O => \N__11527\,
            I => \N__11519\
        );

    \I__2755\ : Span12Mux_v
    port map (
            O => \N__11522\,
            I => \N__11516\
        );

    \I__2754\ : IoSpan4Mux
    port map (
            O => \N__11519\,
            I => \N__11513\
        );

    \I__2753\ : Odrv12
    port map (
            O => \N__11516\,
            I => \DRA_c_2\
        );

    \I__2752\ : Odrv4
    port map (
            O => \N__11513\,
            I => \DRA_c_2\
        );

    \I__2751\ : InMux
    port map (
            O => \N__11508\,
            I => \N__11505\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__11505\,
            I => \N__11502\
        );

    \I__2749\ : Span12Mux_h
    port map (
            O => \N__11502\,
            I => \N__11499\
        );

    \I__2748\ : Odrv12
    port map (
            O => \N__11499\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2747\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11490\
        );

    \I__2746\ : InMux
    port map (
            O => \N__11495\,
            I => \N__11487\
        );

    \I__2745\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11484\
        );

    \I__2744\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11481\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__11490\,
            I => \N__11474\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__11487\,
            I => \N__11474\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__11484\,
            I => \N__11474\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__11481\,
            I => \N__11471\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__11474\,
            I => \N__11468\
        );

    \I__2738\ : Span4Mux_v
    port map (
            O => \N__11471\,
            I => \N__11465\
        );

    \I__2737\ : Span4Mux_v
    port map (
            O => \N__11468\,
            I => \N__11462\
        );

    \I__2736\ : Span4Mux_h
    port map (
            O => \N__11465\,
            I => \N__11459\
        );

    \I__2735\ : Sp12to4
    port map (
            O => \N__11462\,
            I => \N__11456\
        );

    \I__2734\ : IoSpan4Mux
    port map (
            O => \N__11459\,
            I => \N__11453\
        );

    \I__2733\ : Odrv12
    port map (
            O => \N__11456\,
            I => \DRA_c_5\
        );

    \I__2732\ : Odrv4
    port map (
            O => \N__11453\,
            I => \DRA_c_5\
        );

    \I__2731\ : InMux
    port map (
            O => \N__11448\,
            I => \N__11444\
        );

    \I__2730\ : InMux
    port map (
            O => \N__11447\,
            I => \N__11441\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__11444\,
            I => \N__11434\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__11441\,
            I => \N__11434\
        );

    \I__2727\ : InMux
    port map (
            O => \N__11440\,
            I => \N__11431\
        );

    \I__2726\ : InMux
    port map (
            O => \N__11439\,
            I => \N__11428\
        );

    \I__2725\ : Span4Mux_h
    port map (
            O => \N__11434\,
            I => \N__11423\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__11431\,
            I => \N__11423\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__11428\,
            I => \N__11420\
        );

    \I__2722\ : Span4Mux_h
    port map (
            O => \N__11423\,
            I => \N__11417\
        );

    \I__2721\ : Span4Mux_v
    port map (
            O => \N__11420\,
            I => \N__11414\
        );

    \I__2720\ : Span4Mux_v
    port map (
            O => \N__11417\,
            I => \N__11411\
        );

    \I__2719\ : Sp12to4
    port map (
            O => \N__11414\,
            I => \N__11408\
        );

    \I__2718\ : Span4Mux_h
    port map (
            O => \N__11411\,
            I => \N__11405\
        );

    \I__2717\ : Odrv12
    port map (
            O => \N__11408\,
            I => \DRA_c_6\
        );

    \I__2716\ : Odrv4
    port map (
            O => \N__11405\,
            I => \DRA_c_6\
        );

    \I__2715\ : InMux
    port map (
            O => \N__11400\,
            I => \N__11397\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__11397\,
            I => \N__11390\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__11396\,
            I => \N__11387\
        );

    \I__2712\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11380\
        );

    \I__2711\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11370\
        );

    \I__2710\ : InMux
    port map (
            O => \N__11393\,
            I => \N__11370\
        );

    \I__2709\ : Span4Mux_v
    port map (
            O => \N__11390\,
            I => \N__11367\
        );

    \I__2708\ : InMux
    port map (
            O => \N__11387\,
            I => \N__11360\
        );

    \I__2707\ : InMux
    port map (
            O => \N__11386\,
            I => \N__11360\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11385\,
            I => \N__11360\
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__11384\,
            I => \N__11357\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__11383\,
            I => \N__11353\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__11380\,
            I => \N__11347\
        );

    \I__2702\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11344\
        );

    \I__2701\ : InMux
    port map (
            O => \N__11378\,
            I => \N__11339\
        );

    \I__2700\ : InMux
    port map (
            O => \N__11377\,
            I => \N__11339\
        );

    \I__2699\ : InMux
    port map (
            O => \N__11376\,
            I => \N__11334\
        );

    \I__2698\ : InMux
    port map (
            O => \N__11375\,
            I => \N__11334\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__11370\,
            I => \N__11331\
        );

    \I__2696\ : Span4Mux_h
    port map (
            O => \N__11367\,
            I => \N__11326\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__11360\,
            I => \N__11326\
        );

    \I__2694\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11317\
        );

    \I__2693\ : InMux
    port map (
            O => \N__11356\,
            I => \N__11317\
        );

    \I__2692\ : InMux
    port map (
            O => \N__11353\,
            I => \N__11317\
        );

    \I__2691\ : InMux
    port map (
            O => \N__11352\,
            I => \N__11317\
        );

    \I__2690\ : InMux
    port map (
            O => \N__11351\,
            I => \N__11314\
        );

    \I__2689\ : InMux
    port map (
            O => \N__11350\,
            I => \N__11311\
        );

    \I__2688\ : Span4Mux_v
    port map (
            O => \N__11347\,
            I => \N__11308\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__11344\,
            I => \N__11305\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__11339\,
            I => \N__11299\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__11334\,
            I => \N__11299\
        );

    \I__2684\ : Span4Mux_h
    port map (
            O => \N__11331\,
            I => \N__11286\
        );

    \I__2683\ : Span4Mux_v
    port map (
            O => \N__11326\,
            I => \N__11286\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__11317\,
            I => \N__11286\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__11314\,
            I => \N__11286\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__11311\,
            I => \N__11286\
        );

    \I__2679\ : Span4Mux_h
    port map (
            O => \N__11308\,
            I => \N__11281\
        );

    \I__2678\ : Span4Mux_v
    port map (
            O => \N__11305\,
            I => \N__11281\
        );

    \I__2677\ : InMux
    port map (
            O => \N__11304\,
            I => \N__11278\
        );

    \I__2676\ : Span4Mux_v
    port map (
            O => \N__11299\,
            I => \N__11275\
        );

    \I__2675\ : InMux
    port map (
            O => \N__11298\,
            I => \N__11272\
        );

    \I__2674\ : InMux
    port map (
            O => \N__11297\,
            I => \N__11269\
        );

    \I__2673\ : Span4Mux_h
    port map (
            O => \N__11286\,
            I => \N__11266\
        );

    \I__2672\ : Sp12to4
    port map (
            O => \N__11281\,
            I => \N__11263\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__11278\,
            I => \N__11254\
        );

    \I__2670\ : Sp12to4
    port map (
            O => \N__11275\,
            I => \N__11254\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__11272\,
            I => \N__11254\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__11269\,
            I => \N__11254\
        );

    \I__2667\ : Span4Mux_h
    port map (
            O => \N__11266\,
            I => \N__11251\
        );

    \I__2666\ : Span12Mux_h
    port map (
            O => \N__11263\,
            I => \N__11248\
        );

    \I__2665\ : Span12Mux_h
    port map (
            O => \N__11254\,
            I => \N__11243\
        );

    \I__2664\ : Sp12to4
    port map (
            O => \N__11251\,
            I => \N__11243\
        );

    \I__2663\ : Span12Mux_v
    port map (
            O => \N__11248\,
            I => \N__11240\
        );

    \I__2662\ : Span12Mux_v
    port map (
            O => \N__11243\,
            I => \N__11237\
        );

    \I__2661\ : Odrv12
    port map (
            O => \N__11240\,
            I => \AGNUS_REV_c\
        );

    \I__2660\ : Odrv12
    port map (
            O => \N__11237\,
            I => \AGNUS_REV_c\
        );

    \I__2659\ : InMux
    port map (
            O => \N__11232\,
            I => \N__11228\
        );

    \I__2658\ : InMux
    port map (
            O => \N__11231\,
            I => \N__11225\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__11228\,
            I => \N__11222\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__11225\,
            I => \N__11219\
        );

    \I__2655\ : Span4Mux_h
    port map (
            O => \N__11222\,
            I => \N__11216\
        );

    \I__2654\ : Span4Mux_h
    port map (
            O => \N__11219\,
            I => \N__11213\
        );

    \I__2653\ : Odrv4
    port map (
            O => \N__11216\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__11213\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2651\ : ClkMux
    port map (
            O => \N__11208\,
            I => \N__11190\
        );

    \I__2650\ : ClkMux
    port map (
            O => \N__11207\,
            I => \N__11190\
        );

    \I__2649\ : ClkMux
    port map (
            O => \N__11206\,
            I => \N__11190\
        );

    \I__2648\ : ClkMux
    port map (
            O => \N__11205\,
            I => \N__11190\
        );

    \I__2647\ : ClkMux
    port map (
            O => \N__11204\,
            I => \N__11190\
        );

    \I__2646\ : ClkMux
    port map (
            O => \N__11203\,
            I => \N__11190\
        );

    \I__2645\ : GlobalMux
    port map (
            O => \N__11190\,
            I => \N__11187\
        );

    \I__2644\ : gio2CtrlBuf
    port map (
            O => \N__11187\,
            I => \C3_c_g\
        );

    \I__2643\ : CEMux
    port map (
            O => \N__11184\,
            I => \N__11151\
        );

    \I__2642\ : CEMux
    port map (
            O => \N__11183\,
            I => \N__11151\
        );

    \I__2641\ : CEMux
    port map (
            O => \N__11182\,
            I => \N__11151\
        );

    \I__2640\ : CEMux
    port map (
            O => \N__11181\,
            I => \N__11151\
        );

    \I__2639\ : CEMux
    port map (
            O => \N__11180\,
            I => \N__11151\
        );

    \I__2638\ : CEMux
    port map (
            O => \N__11179\,
            I => \N__11151\
        );

    \I__2637\ : CEMux
    port map (
            O => \N__11178\,
            I => \N__11151\
        );

    \I__2636\ : CEMux
    port map (
            O => \N__11177\,
            I => \N__11151\
        );

    \I__2635\ : CEMux
    port map (
            O => \N__11176\,
            I => \N__11151\
        );

    \I__2634\ : CEMux
    port map (
            O => \N__11175\,
            I => \N__11151\
        );

    \I__2633\ : CEMux
    port map (
            O => \N__11174\,
            I => \N__11151\
        );

    \I__2632\ : GlobalMux
    port map (
            O => \N__11151\,
            I => \N__11148\
        );

    \I__2631\ : gio2CtrlBuf
    port map (
            O => \N__11148\,
            I => \DBRn_c_i_0_g\
        );

    \I__2630\ : InMux
    port map (
            O => \N__11145\,
            I => \N__11136\
        );

    \I__2629\ : InMux
    port map (
            O => \N__11144\,
            I => \N__11131\
        );

    \I__2628\ : InMux
    port map (
            O => \N__11143\,
            I => \N__11131\
        );

    \I__2627\ : InMux
    port map (
            O => \N__11142\,
            I => \N__11128\
        );

    \I__2626\ : InMux
    port map (
            O => \N__11141\,
            I => \N__11125\
        );

    \I__2625\ : InMux
    port map (
            O => \N__11140\,
            I => \N__11122\
        );

    \I__2624\ : InMux
    port map (
            O => \N__11139\,
            I => \N__11119\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__11136\,
            I => \N__11099\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__11131\,
            I => \N__11093\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__11128\,
            I => \N__11089\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__11125\,
            I => \N__11086\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__11122\,
            I => \N__11070\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__11119\,
            I => \N__11064\
        );

    \I__2617\ : SRMux
    port map (
            O => \N__11118\,
            I => \N__10971\
        );

    \I__2616\ : SRMux
    port map (
            O => \N__11117\,
            I => \N__10971\
        );

    \I__2615\ : SRMux
    port map (
            O => \N__11116\,
            I => \N__10971\
        );

    \I__2614\ : SRMux
    port map (
            O => \N__11115\,
            I => \N__10971\
        );

    \I__2613\ : SRMux
    port map (
            O => \N__11114\,
            I => \N__10971\
        );

    \I__2612\ : SRMux
    port map (
            O => \N__11113\,
            I => \N__10971\
        );

    \I__2611\ : SRMux
    port map (
            O => \N__11112\,
            I => \N__10971\
        );

    \I__2610\ : SRMux
    port map (
            O => \N__11111\,
            I => \N__10971\
        );

    \I__2609\ : SRMux
    port map (
            O => \N__11110\,
            I => \N__10971\
        );

    \I__2608\ : SRMux
    port map (
            O => \N__11109\,
            I => \N__10971\
        );

    \I__2607\ : SRMux
    port map (
            O => \N__11108\,
            I => \N__10971\
        );

    \I__2606\ : SRMux
    port map (
            O => \N__11107\,
            I => \N__10971\
        );

    \I__2605\ : SRMux
    port map (
            O => \N__11106\,
            I => \N__10971\
        );

    \I__2604\ : SRMux
    port map (
            O => \N__11105\,
            I => \N__10971\
        );

    \I__2603\ : SRMux
    port map (
            O => \N__11104\,
            I => \N__10971\
        );

    \I__2602\ : SRMux
    port map (
            O => \N__11103\,
            I => \N__10971\
        );

    \I__2601\ : SRMux
    port map (
            O => \N__11102\,
            I => \N__10971\
        );

    \I__2600\ : Glb2LocalMux
    port map (
            O => \N__11099\,
            I => \N__10971\
        );

    \I__2599\ : SRMux
    port map (
            O => \N__11098\,
            I => \N__10971\
        );

    \I__2598\ : SRMux
    port map (
            O => \N__11097\,
            I => \N__10971\
        );

    \I__2597\ : SRMux
    port map (
            O => \N__11096\,
            I => \N__10971\
        );

    \I__2596\ : Glb2LocalMux
    port map (
            O => \N__11093\,
            I => \N__10971\
        );

    \I__2595\ : SRMux
    port map (
            O => \N__11092\,
            I => \N__10971\
        );

    \I__2594\ : Glb2LocalMux
    port map (
            O => \N__11089\,
            I => \N__10971\
        );

    \I__2593\ : Glb2LocalMux
    port map (
            O => \N__11086\,
            I => \N__10971\
        );

    \I__2592\ : SRMux
    port map (
            O => \N__11085\,
            I => \N__10971\
        );

    \I__2591\ : SRMux
    port map (
            O => \N__11084\,
            I => \N__10971\
        );

    \I__2590\ : SRMux
    port map (
            O => \N__11083\,
            I => \N__10971\
        );

    \I__2589\ : SRMux
    port map (
            O => \N__11082\,
            I => \N__10971\
        );

    \I__2588\ : SRMux
    port map (
            O => \N__11081\,
            I => \N__10971\
        );

    \I__2587\ : SRMux
    port map (
            O => \N__11080\,
            I => \N__10971\
        );

    \I__2586\ : SRMux
    port map (
            O => \N__11079\,
            I => \N__10971\
        );

    \I__2585\ : SRMux
    port map (
            O => \N__11078\,
            I => \N__10971\
        );

    \I__2584\ : SRMux
    port map (
            O => \N__11077\,
            I => \N__10971\
        );

    \I__2583\ : SRMux
    port map (
            O => \N__11076\,
            I => \N__10971\
        );

    \I__2582\ : SRMux
    port map (
            O => \N__11075\,
            I => \N__10971\
        );

    \I__2581\ : SRMux
    port map (
            O => \N__11074\,
            I => \N__10971\
        );

    \I__2580\ : SRMux
    port map (
            O => \N__11073\,
            I => \N__10971\
        );

    \I__2579\ : Glb2LocalMux
    port map (
            O => \N__11070\,
            I => \N__10971\
        );

    \I__2578\ : SRMux
    port map (
            O => \N__11069\,
            I => \N__10971\
        );

    \I__2577\ : SRMux
    port map (
            O => \N__11068\,
            I => \N__10971\
        );

    \I__2576\ : SRMux
    port map (
            O => \N__11067\,
            I => \N__10971\
        );

    \I__2575\ : Glb2LocalMux
    port map (
            O => \N__11064\,
            I => \N__10971\
        );

    \I__2574\ : SRMux
    port map (
            O => \N__11063\,
            I => \N__10971\
        );

    \I__2573\ : SRMux
    port map (
            O => \N__11062\,
            I => \N__10971\
        );

    \I__2572\ : GlobalMux
    port map (
            O => \N__10971\,
            I => \N__10968\
        );

    \I__2571\ : gio2CtrlBuf
    port map (
            O => \N__10968\,
            I => \RESETn_c_i_g\
        );

    \I__2570\ : InMux
    port map (
            O => \N__10965\,
            I => \N__10960\
        );

    \I__2569\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10956\
        );

    \I__2568\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10952\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__10960\,
            I => \N__10949\
        );

    \I__2566\ : InMux
    port map (
            O => \N__10959\,
            I => \N__10946\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__10956\,
            I => \N__10943\
        );

    \I__2564\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10940\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__10952\,
            I => \N__10935\
        );

    \I__2562\ : Span4Mux_v
    port map (
            O => \N__10949\,
            I => \N__10935\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__10946\,
            I => \N__10932\
        );

    \I__2560\ : Span4Mux_v
    port map (
            O => \N__10943\,
            I => \N__10929\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__10940\,
            I => \N__10926\
        );

    \I__2558\ : Span4Mux_h
    port map (
            O => \N__10935\,
            I => \N__10923\
        );

    \I__2557\ : Span4Mux_v
    port map (
            O => \N__10932\,
            I => \N__10920\
        );

    \I__2556\ : Sp12to4
    port map (
            O => \N__10929\,
            I => \N__10917\
        );

    \I__2555\ : Sp12to4
    port map (
            O => \N__10926\,
            I => \N__10914\
        );

    \I__2554\ : Sp12to4
    port map (
            O => \N__10923\,
            I => \N__10909\
        );

    \I__2553\ : Sp12to4
    port map (
            O => \N__10920\,
            I => \N__10909\
        );

    \I__2552\ : Span12Mux_h
    port map (
            O => \N__10917\,
            I => \N__10904\
        );

    \I__2551\ : Span12Mux_v
    port map (
            O => \N__10914\,
            I => \N__10904\
        );

    \I__2550\ : Span12Mux_h
    port map (
            O => \N__10909\,
            I => \N__10901\
        );

    \I__2549\ : Span12Mux_h
    port map (
            O => \N__10904\,
            I => \N__10896\
        );

    \I__2548\ : Span12Mux_v
    port map (
            O => \N__10901\,
            I => \N__10896\
        );

    \I__2547\ : Odrv12
    port map (
            O => \N__10896\,
            I => \RnW_c\
        );

    \I__2546\ : InMux
    port map (
            O => \N__10893\,
            I => \N__10890\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__10890\,
            I => \N__10886\
        );

    \I__2544\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10883\
        );

    \I__2543\ : Span4Mux_v
    port map (
            O => \N__10886\,
            I => \N__10878\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__10883\,
            I => \N__10875\
        );

    \I__2541\ : InMux
    port map (
            O => \N__10882\,
            I => \N__10870\
        );

    \I__2540\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10870\
        );

    \I__2539\ : Span4Mux_v
    port map (
            O => \N__10878\,
            I => \N__10864\
        );

    \I__2538\ : Span4Mux_v
    port map (
            O => \N__10875\,
            I => \N__10864\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__10870\,
            I => \N__10861\
        );

    \I__2536\ : InMux
    port map (
            O => \N__10869\,
            I => \N__10858\
        );

    \I__2535\ : Span4Mux_h
    port map (
            O => \N__10864\,
            I => \N__10852\
        );

    \I__2534\ : Span4Mux_h
    port map (
            O => \N__10861\,
            I => \N__10852\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10858\,
            I => \N__10849\
        );

    \I__2532\ : InMux
    port map (
            O => \N__10857\,
            I => \N__10846\
        );

    \I__2531\ : Sp12to4
    port map (
            O => \N__10852\,
            I => \N__10843\
        );

    \I__2530\ : Span12Mux_v
    port map (
            O => \N__10849\,
            I => \N__10840\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10846\,
            I => \N__10837\
        );

    \I__2528\ : Span12Mux_v
    port map (
            O => \N__10843\,
            I => \N__10834\
        );

    \I__2527\ : Span12Mux_h
    port map (
            O => \N__10840\,
            I => \N__10831\
        );

    \I__2526\ : Span4Mux_v
    port map (
            O => \N__10837\,
            I => \N__10828\
        );

    \I__2525\ : Odrv12
    port map (
            O => \N__10834\,
            I => \CASUn_c\
        );

    \I__2524\ : Odrv12
    port map (
            O => \N__10831\,
            I => \CASUn_c\
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__10828\,
            I => \CASUn_c\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__10821\,
            I => \N__10818\
        );

    \I__2521\ : InMux
    port map (
            O => \N__10818\,
            I => \N__10815\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__10815\,
            I => \N__10811\
        );

    \I__2519\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10808\
        );

    \I__2518\ : Span12Mux_s7_v
    port map (
            O => \N__10811\,
            I => \N__10804\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__10808\,
            I => \N__10801\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__10807\,
            I => \N__10798\
        );

    \I__2515\ : Span12Mux_v
    port map (
            O => \N__10804\,
            I => \N__10795\
        );

    \I__2514\ : Span12Mux_v
    port map (
            O => \N__10801\,
            I => \N__10792\
        );

    \I__2513\ : InMux
    port map (
            O => \N__10798\,
            I => \N__10789\
        );

    \I__2512\ : Odrv12
    port map (
            O => \N__10795\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2511\ : Odrv12
    port map (
            O => \N__10792\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10789\,
            I => \DMA_WRITE_CYCLE\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__10782\,
            I => \N__10779\
        );

    \I__2508\ : InMux
    port map (
            O => \N__10779\,
            I => \N__10772\
        );

    \I__2507\ : InMux
    port map (
            O => \N__10778\,
            I => \N__10772\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10777\,
            I => \N__10767\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__10772\,
            I => \N__10764\
        );

    \I__2504\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10759\
        );

    \I__2503\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10759\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10767\,
            I => \N__10756\
        );

    \I__2501\ : Span4Mux_h
    port map (
            O => \N__10764\,
            I => \N__10753\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__10759\,
            I => \N__10750\
        );

    \I__2499\ : Span4Mux_h
    port map (
            O => \N__10756\,
            I => \N__10747\
        );

    \I__2498\ : Sp12to4
    port map (
            O => \N__10753\,
            I => \N__10743\
        );

    \I__2497\ : Span12Mux_v
    port map (
            O => \N__10750\,
            I => \N__10740\
        );

    \I__2496\ : Span4Mux_v
    port map (
            O => \N__10747\,
            I => \N__10737\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10746\,
            I => \N__10734\
        );

    \I__2494\ : Span12Mux_v
    port map (
            O => \N__10743\,
            I => \N__10731\
        );

    \I__2493\ : Span12Mux_h
    port map (
            O => \N__10740\,
            I => \N__10728\
        );

    \I__2492\ : Sp12to4
    port map (
            O => \N__10737\,
            I => \N__10725\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__10734\,
            I => \N__10722\
        );

    \I__2490\ : Span12Mux_h
    port map (
            O => \N__10731\,
            I => \N__10717\
        );

    \I__2489\ : Span12Mux_v
    port map (
            O => \N__10728\,
            I => \N__10717\
        );

    \I__2488\ : Span12Mux_h
    port map (
            O => \N__10725\,
            I => \N__10712\
        );

    \I__2487\ : Span12Mux_v
    port map (
            O => \N__10722\,
            I => \N__10712\
        );

    \I__2486\ : Odrv12
    port map (
            O => \N__10717\,
            I => \CASLn_c\
        );

    \I__2485\ : Odrv12
    port map (
            O => \N__10712\,
            I => \CASLn_c\
        );

    \I__2484\ : IoInMux
    port map (
            O => \N__10707\,
            I => \N__10704\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10704\,
            I => \N__10701\
        );

    \I__2482\ : IoSpan4Mux
    port map (
            O => \N__10701\,
            I => \N__10698\
        );

    \I__2481\ : IoSpan4Mux
    port map (
            O => \N__10698\,
            I => \N__10695\
        );

    \I__2480\ : Span4Mux_s3_v
    port map (
            O => \N__10695\,
            I => \N__10692\
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__10692\,
            I => \N_409\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10686\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__10686\,
            I => \N__10683\
        );

    \I__2476\ : Odrv12
    port map (
            O => \N__10683\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2475\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10677\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__10677\,
            I => \N__10674\
        );

    \I__2473\ : Span4Mux_h
    port map (
            O => \N__10674\,
            I => \N__10671\
        );

    \I__2472\ : Span4Mux_v
    port map (
            O => \N__10671\,
            I => \N__10668\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__10668\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10662\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__10662\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2468\ : InMux
    port map (
            O => \N__10659\,
            I => \N__10655\
        );

    \I__2467\ : InMux
    port map (
            O => \N__10658\,
            I => \N__10650\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10655\,
            I => \N__10647\
        );

    \I__2465\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10644\
        );

    \I__2464\ : InMux
    port map (
            O => \N__10653\,
            I => \N__10641\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__10650\,
            I => \N__10638\
        );

    \I__2462\ : Span4Mux_v
    port map (
            O => \N__10647\,
            I => \N__10631\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__10644\,
            I => \N__10631\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__10641\,
            I => \N__10631\
        );

    \I__2459\ : Span12Mux_h
    port map (
            O => \N__10638\,
            I => \N__10628\
        );

    \I__2458\ : Sp12to4
    port map (
            O => \N__10631\,
            I => \N__10625\
        );

    \I__2457\ : Span12Mux_v
    port map (
            O => \N__10628\,
            I => \N__10622\
        );

    \I__2456\ : Span12Mux_v
    port map (
            O => \N__10625\,
            I => \N__10619\
        );

    \I__2455\ : Odrv12
    port map (
            O => \N__10622\,
            I => \DRA_c_1\
        );

    \I__2454\ : Odrv12
    port map (
            O => \N__10619\,
            I => \DRA_c_1\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10614\,
            I => \N__10611\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__10611\,
            I => \N__10608\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__10608\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2450\ : InMux
    port map (
            O => \N__10605\,
            I => \N__10602\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__10602\,
            I => \N__10596\
        );

    \I__2448\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10591\
        );

    \I__2447\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10591\
        );

    \I__2446\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10587\
        );

    \I__2445\ : Span4Mux_v
    port map (
            O => \N__10596\,
            I => \N__10582\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__10591\,
            I => \N__10582\
        );

    \I__2443\ : InMux
    port map (
            O => \N__10590\,
            I => \N__10579\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__10587\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__10582\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__10579\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2439\ : IoInMux
    port map (
            O => \N__10572\,
            I => \N__10569\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__10569\,
            I => \N__10566\
        );

    \I__2437\ : IoSpan4Mux
    port map (
            O => \N__10566\,
            I => \N__10563\
        );

    \I__2436\ : Sp12to4
    port map (
            O => \N__10563\,
            I => \N__10560\
        );

    \I__2435\ : Span12Mux_s9_v
    port map (
            O => \N__10560\,
            I => \N__10557\
        );

    \I__2434\ : Odrv12
    port map (
            O => \N__10557\,
            I => \WEn_c\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10554\,
            I => \N__10551\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__10551\,
            I => \U712_CHIP_RAM.CMA_5_i_0_9\
        );

    \I__2431\ : InMux
    port map (
            O => \N__10548\,
            I => \N__10545\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__10545\,
            I => \N__10542\
        );

    \I__2429\ : Sp12to4
    port map (
            O => \N__10542\,
            I => \N__10539\
        );

    \I__2428\ : Span12Mux_v
    port map (
            O => \N__10539\,
            I => \N__10536\
        );

    \I__2427\ : Span12Mux_h
    port map (
            O => \N__10536\,
            I => \N__10533\
        );

    \I__2426\ : Odrv12
    port map (
            O => \N__10533\,
            I => \A_c_19\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__10530\,
            I => \N__10525\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10529\,
            I => \N__10522\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__10528\,
            I => \N__10519\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10525\,
            I => \N__10511\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__10522\,
            I => \N__10507\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10519\,
            I => \N__10504\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__10518\,
            I => \N__10501\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__10517\,
            I => \N__10495\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10516\,
            I => \N__10489\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10515\,
            I => \N__10489\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10514\,
            I => \N__10486\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__10511\,
            I => \N__10480\
        );

    \I__2413\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10477\
        );

    \I__2412\ : Span4Mux_h
    port map (
            O => \N__10507\,
            I => \N__10469\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__10504\,
            I => \N__10469\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10501\,
            I => \N__10463\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10460\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10457\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10498\,
            I => \N__10454\
        );

    \I__2406\ : InMux
    port map (
            O => \N__10495\,
            I => \N__10449\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10494\,
            I => \N__10449\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10489\,
            I => \N__10445\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__10486\,
            I => \N__10442\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__10485\,
            I => \N__10439\
        );

    \I__2401\ : InMux
    port map (
            O => \N__10484\,
            I => \N__10436\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10483\,
            I => \N__10432\
        );

    \I__2399\ : Span4Mux_v
    port map (
            O => \N__10480\,
            I => \N__10429\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__10477\,
            I => \N__10426\
        );

    \I__2397\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10423\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10475\,
            I => \N__10418\
        );

    \I__2395\ : InMux
    port map (
            O => \N__10474\,
            I => \N__10418\
        );

    \I__2394\ : Span4Mux_v
    port map (
            O => \N__10469\,
            I => \N__10415\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10468\,
            I => \N__10412\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10467\,
            I => \N__10407\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10466\,
            I => \N__10407\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__10463\,
            I => \N__10402\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__10460\,
            I => \N__10402\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__10457\,
            I => \N__10399\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10454\,
            I => \N__10396\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__10449\,
            I => \N__10393\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10448\,
            I => \N__10390\
        );

    \I__2384\ : Span4Mux_v
    port map (
            O => \N__10445\,
            I => \N__10384\
        );

    \I__2383\ : Span4Mux_v
    port map (
            O => \N__10442\,
            I => \N__10384\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10381\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10436\,
            I => \N__10378\
        );

    \I__2380\ : InMux
    port map (
            O => \N__10435\,
            I => \N__10375\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10432\,
            I => \N__10368\
        );

    \I__2378\ : Span4Mux_h
    port map (
            O => \N__10429\,
            I => \N__10368\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__10426\,
            I => \N__10368\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__10423\,
            I => \N__10359\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__10418\,
            I => \N__10359\
        );

    \I__2374\ : Sp12to4
    port map (
            O => \N__10415\,
            I => \N__10359\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__10412\,
            I => \N__10359\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10407\,
            I => \N__10354\
        );

    \I__2371\ : Span12Mux_h
    port map (
            O => \N__10402\,
            I => \N__10354\
        );

    \I__2370\ : Span4Mux_v
    port map (
            O => \N__10399\,
            I => \N__10345\
        );

    \I__2369\ : Span4Mux_h
    port map (
            O => \N__10396\,
            I => \N__10345\
        );

    \I__2368\ : Span4Mux_h
    port map (
            O => \N__10393\,
            I => \N__10345\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10390\,
            I => \N__10345\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10342\
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__10384\,
            I => \CPU_CYCLEm\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__10381\,
            I => \CPU_CYCLEm\
        );

    \I__2363\ : Odrv4
    port map (
            O => \N__10378\,
            I => \CPU_CYCLEm\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10375\,
            I => \CPU_CYCLEm\
        );

    \I__2361\ : Odrv4
    port map (
            O => \N__10368\,
            I => \CPU_CYCLEm\
        );

    \I__2360\ : Odrv12
    port map (
            O => \N__10359\,
            I => \CPU_CYCLEm\
        );

    \I__2359\ : Odrv12
    port map (
            O => \N__10354\,
            I => \CPU_CYCLEm\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__10345\,
            I => \CPU_CYCLEm\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10342\,
            I => \CPU_CYCLEm\
        );

    \I__2356\ : IoInMux
    port map (
            O => \N__10323\,
            I => \N__10320\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__10320\,
            I => \N__10317\
        );

    \I__2354\ : IoSpan4Mux
    port map (
            O => \N__10317\,
            I => \N__10314\
        );

    \I__2353\ : Sp12to4
    port map (
            O => \N__10314\,
            I => \N__10311\
        );

    \I__2352\ : Span12Mux_s9_h
    port map (
            O => \N__10311\,
            I => \N__10308\
        );

    \I__2351\ : Odrv12
    port map (
            O => \N__10308\,
            I => \CMA_c_9\
        );

    \I__2350\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10302\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__10302\,
            I => \N__10298\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10301\,
            I => \N__10295\
        );

    \I__2347\ : Span4Mux_h
    port map (
            O => \N__10298\,
            I => \N__10286\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10295\,
            I => \N__10283\
        );

    \I__2345\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10276\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10293\,
            I => \N__10276\
        );

    \I__2343\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10276\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10291\,
            I => \N__10273\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10290\,
            I => \N__10270\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10289\,
            I => \N__10267\
        );

    \I__2339\ : Span4Mux_h
    port map (
            O => \N__10286\,
            I => \N__10260\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__10283\,
            I => \N__10260\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__10276\,
            I => \N__10257\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__10273\,
            I => \N__10254\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__10270\,
            I => \N__10249\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__10267\,
            I => \N__10249\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10266\,
            I => \N__10246\
        );

    \I__2332\ : InMux
    port map (
            O => \N__10265\,
            I => \N__10243\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__10260\,
            I => \U712_CHIP_RAM.N_354\
        );

    \I__2330\ : Odrv12
    port map (
            O => \N__10257\,
            I => \U712_CHIP_RAM.N_354\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__10254\,
            I => \U712_CHIP_RAM.N_354\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__10249\,
            I => \U712_CHIP_RAM.N_354\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__10246\,
            I => \U712_CHIP_RAM.N_354\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__10243\,
            I => \U712_CHIP_RAM.N_354\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__10230\,
            I => \N__10224\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__10229\,
            I => \N__10221\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__10228\,
            I => \N__10218\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__10227\,
            I => \N__10215\
        );

    \I__2321\ : InMux
    port map (
            O => \N__10224\,
            I => \N__10212\
        );

    \I__2320\ : InMux
    port map (
            O => \N__10221\,
            I => \N__10209\
        );

    \I__2319\ : InMux
    port map (
            O => \N__10218\,
            I => \N__10204\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10215\,
            I => \N__10201\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__10212\,
            I => \N__10198\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__10209\,
            I => \N__10195\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__10208\,
            I => \N__10191\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__10207\,
            I => \N__10188\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__10204\,
            I => \N__10185\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__10201\,
            I => \N__10182\
        );

    \I__2311\ : Span4Mux_v
    port map (
            O => \N__10198\,
            I => \N__10179\
        );

    \I__2310\ : Span4Mux_v
    port map (
            O => \N__10195\,
            I => \N__10176\
        );

    \I__2309\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10173\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10191\,
            I => \N__10168\
        );

    \I__2307\ : InMux
    port map (
            O => \N__10188\,
            I => \N__10168\
        );

    \I__2306\ : Span4Mux_v
    port map (
            O => \N__10185\,
            I => \N__10165\
        );

    \I__2305\ : Span12Mux_s11_v
    port map (
            O => \N__10182\,
            I => \N__10162\
        );

    \I__2304\ : Span4Mux_h
    port map (
            O => \N__10179\,
            I => \N__10157\
        );

    \I__2303\ : Span4Mux_h
    port map (
            O => \N__10176\,
            I => \N__10157\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__10173\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10168\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__10165\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__2299\ : Odrv12
    port map (
            O => \N__10162\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__10157\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__2297\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10143\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__10143\,
            I => \N__10140\
        );

    \I__2295\ : Span4Mux_h
    port map (
            O => \N__10140\,
            I => \N__10137\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__10137\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__2293\ : IoInMux
    port map (
            O => \N__10134\,
            I => \N__10131\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__10131\,
            I => \N__10128\
        );

    \I__2291\ : IoSpan4Mux
    port map (
            O => \N__10128\,
            I => \N__10125\
        );

    \I__2290\ : IoSpan4Mux
    port map (
            O => \N__10125\,
            I => \N__10122\
        );

    \I__2289\ : Sp12to4
    port map (
            O => \N__10122\,
            I => \N__10119\
        );

    \I__2288\ : Span12Mux_s9_h
    port map (
            O => \N__10119\,
            I => \N__10116\
        );

    \I__2287\ : Odrv12
    port map (
            O => \N__10116\,
            I => \CMA_c_4\
        );

    \I__2286\ : CEMux
    port map (
            O => \N__10113\,
            I => \N__10109\
        );

    \I__2285\ : CEMux
    port map (
            O => \N__10112\,
            I => \N__10105\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__10109\,
            I => \N__10102\
        );

    \I__2283\ : CEMux
    port map (
            O => \N__10108\,
            I => \N__10099\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__10105\,
            I => \N__10093\
        );

    \I__2281\ : Span4Mux_v
    port map (
            O => \N__10102\,
            I => \N__10088\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__10099\,
            I => \N__10088\
        );

    \I__2279\ : CEMux
    port map (
            O => \N__10098\,
            I => \N__10085\
        );

    \I__2278\ : CEMux
    port map (
            O => \N__10097\,
            I => \N__10081\
        );

    \I__2277\ : CEMux
    port map (
            O => \N__10096\,
            I => \N__10077\
        );

    \I__2276\ : Span4Mux_h
    port map (
            O => \N__10093\,
            I => \N__10070\
        );

    \I__2275\ : Span4Mux_h
    port map (
            O => \N__10088\,
            I => \N__10070\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__10085\,
            I => \N__10070\
        );

    \I__2273\ : CEMux
    port map (
            O => \N__10084\,
            I => \N__10067\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__10081\,
            I => \N__10064\
        );

    \I__2271\ : CEMux
    port map (
            O => \N__10080\,
            I => \N__10061\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__10077\,
            I => \N__10058\
        );

    \I__2269\ : Span4Mux_h
    port map (
            O => \N__10070\,
            I => \N__10053\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__10067\,
            I => \N__10053\
        );

    \I__2267\ : Span4Mux_h
    port map (
            O => \N__10064\,
            I => \N__10050\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__10061\,
            I => \N__10047\
        );

    \I__2265\ : Span4Mux_h
    port map (
            O => \N__10058\,
            I => \N__10042\
        );

    \I__2264\ : Span4Mux_h
    port map (
            O => \N__10053\,
            I => \N__10042\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__10050\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2262\ : Odrv4
    port map (
            O => \N__10047\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__10042\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_0\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__10035\,
            I => \N__10031\
        );

    \I__2259\ : InMux
    port map (
            O => \N__10034\,
            I => \N__10027\
        );

    \I__2258\ : InMux
    port map (
            O => \N__10031\,
            I => \N__10023\
        );

    \I__2257\ : InMux
    port map (
            O => \N__10030\,
            I => \N__10020\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__10027\,
            I => \N__10017\
        );

    \I__2255\ : InMux
    port map (
            O => \N__10026\,
            I => \N__10014\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__10023\,
            I => \N__10011\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__10020\,
            I => \N__10004\
        );

    \I__2252\ : Span4Mux_h
    port map (
            O => \N__10017\,
            I => \N__10004\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__10014\,
            I => \N__10004\
        );

    \I__2250\ : Span4Mux_v
    port map (
            O => \N__10011\,
            I => \N__10001\
        );

    \I__2249\ : Span4Mux_v
    port map (
            O => \N__10004\,
            I => \N__9998\
        );

    \I__2248\ : Sp12to4
    port map (
            O => \N__10001\,
            I => \N__9993\
        );

    \I__2247\ : Sp12to4
    port map (
            O => \N__9998\,
            I => \N__9993\
        );

    \I__2246\ : Span12Mux_h
    port map (
            O => \N__9993\,
            I => \N__9990\
        );

    \I__2245\ : Span12Mux_v
    port map (
            O => \N__9990\,
            I => \N__9987\
        );

    \I__2244\ : Odrv12
    port map (
            O => \N__9987\,
            I => \DRA_c_9\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9984\,
            I => \N__9981\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__9981\,
            I => \N__9978\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__9978\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9975\,
            I => \N__9972\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__9972\,
            I => \N__9966\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9971\,
            I => \N__9963\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9970\,
            I => \N__9960\
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__9969\,
            I => \N__9956\
        );

    \I__2235\ : Span4Mux_v
    port map (
            O => \N__9966\,
            I => \N__9951\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__9963\,
            I => \N__9951\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__9960\,
            I => \N__9948\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__9959\,
            I => \N__9945\
        );

    \I__2231\ : InMux
    port map (
            O => \N__9956\,
            I => \N__9942\
        );

    \I__2230\ : Span4Mux_h
    port map (
            O => \N__9951\,
            I => \N__9939\
        );

    \I__2229\ : Span4Mux_v
    port map (
            O => \N__9948\,
            I => \N__9936\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9933\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__9942\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2226\ : Odrv4
    port map (
            O => \N__9939\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2225\ : Odrv4
    port map (
            O => \N__9936\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__9933\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2223\ : IoInMux
    port map (
            O => \N__9924\,
            I => \N__9921\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__9921\,
            I => \N__9918\
        );

    \I__2221\ : Span4Mux_s1_v
    port map (
            O => \N__9918\,
            I => \N__9915\
        );

    \I__2220\ : Span4Mux_v
    port map (
            O => \N__9915\,
            I => \N__9912\
        );

    \I__2219\ : Span4Mux_v
    port map (
            O => \N__9912\,
            I => \N__9909\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__9909\,
            I => \CMA_c_10\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__9906\,
            I => \N__9902\
        );

    \I__2216\ : InMux
    port map (
            O => \N__9905\,
            I => \N__9899\
        );

    \I__2215\ : InMux
    port map (
            O => \N__9902\,
            I => \N__9894\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__9899\,
            I => \N__9890\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9898\,
            I => \N__9887\
        );

    \I__2212\ : InMux
    port map (
            O => \N__9897\,
            I => \N__9884\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__9894\,
            I => \N__9881\
        );

    \I__2210\ : InMux
    port map (
            O => \N__9893\,
            I => \N__9877\
        );

    \I__2209\ : Span4Mux_v
    port map (
            O => \N__9890\,
            I => \N__9870\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__9887\,
            I => \N__9870\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__9884\,
            I => \N__9870\
        );

    \I__2206\ : Span4Mux_h
    port map (
            O => \N__9881\,
            I => \N__9867\
        );

    \I__2205\ : InMux
    port map (
            O => \N__9880\,
            I => \N__9864\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__9877\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__9870\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__9867\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__9864\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__9855\,
            I => \U712_CHIP_RAM.N_354_cascade_\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__9852\,
            I => \N__9841\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__9851\,
            I => \N__9838\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__9850\,
            I => \N__9832\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__9849\,
            I => \N__9829\
        );

    \I__2195\ : CascadeMux
    port map (
            O => \N__9848\,
            I => \N__9826\
        );

    \I__2194\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9817\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9814\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9845\,
            I => \N__9809\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9844\,
            I => \N__9809\
        );

    \I__2190\ : InMux
    port map (
            O => \N__9841\,
            I => \N__9805\
        );

    \I__2189\ : InMux
    port map (
            O => \N__9838\,
            I => \N__9802\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9837\,
            I => \N__9799\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9794\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9835\,
            I => \N__9794\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9832\,
            I => \N__9789\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9829\,
            I => \N__9789\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9826\,
            I => \N__9784\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9825\,
            I => \N__9784\
        );

    \I__2181\ : InMux
    port map (
            O => \N__9824\,
            I => \N__9777\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9823\,
            I => \N__9777\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9822\,
            I => \N__9777\
        );

    \I__2178\ : InMux
    port map (
            O => \N__9821\,
            I => \N__9774\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9820\,
            I => \N__9771\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9817\,
            I => \N__9761\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__9814\,
            I => \N__9761\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__9809\,
            I => \N__9761\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9808\,
            I => \N__9758\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9805\,
            I => \N__9755\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9802\,
            I => \N__9752\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9799\,
            I => \N__9749\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9794\,
            I => \N__9746\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__9789\,
            I => \N__9739\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9784\,
            I => \N__9739\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__9777\,
            I => \N__9739\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9774\,
            I => \N__9731\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9771\,
            I => \N__9731\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9723\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9769\,
            I => \N__9723\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9768\,
            I => \N__9723\
        );

    \I__2160\ : Span4Mux_v
    port map (
            O => \N__9761\,
            I => \N__9720\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__9758\,
            I => \N__9707\
        );

    \I__2158\ : Span4Mux_v
    port map (
            O => \N__9755\,
            I => \N__9707\
        );

    \I__2157\ : Span4Mux_v
    port map (
            O => \N__9752\,
            I => \N__9707\
        );

    \I__2156\ : Span4Mux_h
    port map (
            O => \N__9749\,
            I => \N__9707\
        );

    \I__2155\ : Span4Mux_v
    port map (
            O => \N__9746\,
            I => \N__9707\
        );

    \I__2154\ : Span4Mux_v
    port map (
            O => \N__9739\,
            I => \N__9707\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9738\,
            I => \N__9700\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9737\,
            I => \N__9700\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9736\,
            I => \N__9700\
        );

    \I__2150\ : Span4Mux_v
    port map (
            O => \N__9731\,
            I => \N__9697\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9730\,
            I => \N__9694\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9723\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__9720\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__9707\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__9700\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2144\ : Odrv4
    port map (
            O => \N__9697\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9694\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9681\,
            I => \N__9678\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9678\,
            I => \N__9675\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__9675\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9672\,
            I => \N__9669\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__9669\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9663\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9663\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__2135\ : IoInMux
    port map (
            O => \N__9660\,
            I => \N__9657\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9657\,
            I => \N__9654\
        );

    \I__2133\ : IoSpan4Mux
    port map (
            O => \N__9654\,
            I => \N__9651\
        );

    \I__2132\ : Span4Mux_s2_h
    port map (
            O => \N__9651\,
            I => \N__9648\
        );

    \I__2131\ : Sp12to4
    port map (
            O => \N__9648\,
            I => \N__9645\
        );

    \I__2130\ : Span12Mux_s10_h
    port map (
            O => \N__9645\,
            I => \N__9642\
        );

    \I__2129\ : Odrv12
    port map (
            O => \N__9642\,
            I => \CMA_c_5\
        );

    \I__2128\ : InMux
    port map (
            O => \N__9639\,
            I => \N__9636\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__9636\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__2126\ : IoInMux
    port map (
            O => \N__9633\,
            I => \N__9630\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__9630\,
            I => \N__9627\
        );

    \I__2124\ : Span4Mux_s1_h
    port map (
            O => \N__9627\,
            I => \N__9624\
        );

    \I__2123\ : Sp12to4
    port map (
            O => \N__9624\,
            I => \N__9621\
        );

    \I__2122\ : Span12Mux_v
    port map (
            O => \N__9621\,
            I => \N__9618\
        );

    \I__2121\ : Odrv12
    port map (
            O => \N__9618\,
            I => \CMA_c_3\
        );

    \I__2120\ : InMux
    port map (
            O => \N__9615\,
            I => \N__9612\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__9612\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2118\ : InMux
    port map (
            O => \N__9609\,
            I => \N__9606\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__9606\,
            I => \N__9603\
        );

    \I__2116\ : Odrv12
    port map (
            O => \N__9603\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2115\ : InMux
    port map (
            O => \N__9600\,
            I => \N__9597\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__9597\,
            I => \N__9594\
        );

    \I__2113\ : Span4Mux_h
    port map (
            O => \N__9594\,
            I => \N__9591\
        );

    \I__2112\ : Odrv4
    port map (
            O => \N__9591\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2111\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9585\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9585\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2109\ : InMux
    port map (
            O => \N__9582\,
            I => \N__9579\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__9579\,
            I => \N__9576\
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__9576\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9573\,
            I => \N__9570\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__9570\,
            I => \N__9567\
        );

    \I__2104\ : Span4Mux_h
    port map (
            O => \N__9567\,
            I => \N__9564\
        );

    \I__2103\ : Span4Mux_v
    port map (
            O => \N__9564\,
            I => \N__9561\
        );

    \I__2102\ : Odrv4
    port map (
            O => \N__9561\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9558\,
            I => \N__9552\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9557\,
            I => \N__9552\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9552\,
            I => \N__9549\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__9549\,
            I => \N__9544\
        );

    \I__2097\ : InMux
    port map (
            O => \N__9548\,
            I => \N__9539\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9547\,
            I => \N__9539\
        );

    \I__2095\ : Sp12to4
    port map (
            O => \N__9544\,
            I => \N__9534\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__9539\,
            I => \N__9534\
        );

    \I__2093\ : Span12Mux_h
    port map (
            O => \N__9534\,
            I => \N__9531\
        );

    \I__2092\ : Odrv12
    port map (
            O => \N__9531\,
            I => \DRA_c_7\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9523\
        );

    \I__2090\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9520\
        );

    \I__2089\ : InMux
    port map (
            O => \N__9526\,
            I => \N__9517\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__9523\,
            I => \N__9509\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__9520\,
            I => \N__9509\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9517\,
            I => \N__9509\
        );

    \I__2085\ : InMux
    port map (
            O => \N__9516\,
            I => \N__9506\
        );

    \I__2084\ : Span4Mux_v
    port map (
            O => \N__9509\,
            I => \N__9503\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9506\,
            I => \N__9500\
        );

    \I__2082\ : Sp12to4
    port map (
            O => \N__9503\,
            I => \N__9497\
        );

    \I__2081\ : Span12Mux_h
    port map (
            O => \N__9500\,
            I => \N__9494\
        );

    \I__2080\ : Odrv12
    port map (
            O => \N__9497\,
            I => \DRA_c_8\
        );

    \I__2079\ : Odrv12
    port map (
            O => \N__9494\,
            I => \DRA_c_8\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__9489\,
            I => \N__9486\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9483\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9483\,
            I => \N__9480\
        );

    \I__2075\ : Span12Mux_v
    port map (
            O => \N__9480\,
            I => \N__9477\
        );

    \I__2074\ : Odrv12
    port map (
            O => \N__9477\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__9474\,
            I => \N__9470\
        );

    \I__2072\ : InMux
    port map (
            O => \N__9473\,
            I => \N__9467\
        );

    \I__2071\ : InMux
    port map (
            O => \N__9470\,
            I => \N__9464\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__9467\,
            I => \N__9461\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__9464\,
            I => \N__9456\
        );

    \I__2068\ : Span4Mux_v
    port map (
            O => \N__9461\,
            I => \N__9456\
        );

    \I__2067\ : Sp12to4
    port map (
            O => \N__9456\,
            I => \N__9453\
        );

    \I__2066\ : Span12Mux_h
    port map (
            O => \N__9453\,
            I => \N__9450\
        );

    \I__2065\ : Span12Mux_v
    port map (
            O => \N__9450\,
            I => \N__9447\
        );

    \I__2064\ : Odrv12
    port map (
            O => \N__9447\,
            I => \DRA_c_0\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9444\,
            I => \N__9441\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9441\,
            I => \N__9438\
        );

    \I__2061\ : Span4Mux_h
    port map (
            O => \N__9438\,
            I => \N__9435\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__9435\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2059\ : IoInMux
    port map (
            O => \N__9432\,
            I => \N__9429\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__9429\,
            I => \N__9426\
        );

    \I__2057\ : Span4Mux_s3_v
    port map (
            O => \N__9426\,
            I => \N__9423\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__9423\,
            I => \N__9420\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__9420\,
            I => \RASn_c\
        );

    \I__2054\ : IoInMux
    port map (
            O => \N__9417\,
            I => \N__9414\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9414\,
            I => \N__9411\
        );

    \I__2052\ : IoSpan4Mux
    port map (
            O => \N__9411\,
            I => \N__9408\
        );

    \I__2051\ : Span4Mux_s3_v
    port map (
            O => \N__9408\,
            I => \N__9405\
        );

    \I__2050\ : Span4Mux_v
    port map (
            O => \N__9405\,
            I => \N__9402\
        );

    \I__2049\ : Odrv4
    port map (
            O => \N__9402\,
            I => \CRCSn_c\
        );

    \I__2048\ : IoInMux
    port map (
            O => \N__9399\,
            I => \N__9396\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9396\,
            I => \N__9393\
        );

    \I__2046\ : Span4Mux_s1_v
    port map (
            O => \N__9393\,
            I => \N__9390\
        );

    \I__2045\ : Sp12to4
    port map (
            O => \N__9390\,
            I => \N__9387\
        );

    \I__2044\ : Span12Mux_s10_h
    port map (
            O => \N__9387\,
            I => \N__9384\
        );

    \I__2043\ : Odrv12
    port map (
            O => \N__9384\,
            I => \CASn_c\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9381\,
            I => \N__9376\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__9380\,
            I => \N__9373\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9379\,
            I => \N__9370\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__9376\,
            I => \N__9367\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9373\,
            I => \N__9364\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__9370\,
            I => \N__9361\
        );

    \I__2036\ : Span4Mux_v
    port map (
            O => \N__9367\,
            I => \N__9357\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9364\,
            I => \N__9354\
        );

    \I__2034\ : Span4Mux_h
    port map (
            O => \N__9361\,
            I => \N__9351\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9348\
        );

    \I__2032\ : Span4Mux_v
    port map (
            O => \N__9357\,
            I => \N__9343\
        );

    \I__2031\ : Span4Mux_h
    port map (
            O => \N__9354\,
            I => \N__9343\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__9351\,
            I => \REG_CYCLEm\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__9348\,
            I => \REG_CYCLEm\
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__9343\,
            I => \REG_CYCLEm\
        );

    \I__2027\ : IoInMux
    port map (
            O => \N__9336\,
            I => \N__9333\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__9333\,
            I => \N__9330\
        );

    \I__2025\ : Span4Mux_s1_v
    port map (
            O => \N__9330\,
            I => \N__9327\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__9327\,
            I => \N__9324\
        );

    \I__2023\ : Sp12to4
    port map (
            O => \N__9324\,
            I => \N__9321\
        );

    \I__2022\ : Span12Mux_h
    port map (
            O => \N__9321\,
            I => \N__9318\
        );

    \I__2021\ : Span12Mux_v
    port map (
            O => \N__9318\,
            I => \N__9315\
        );

    \I__2020\ : Odrv12
    port map (
            O => \N__9315\,
            I => \N_207_i\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9312\,
            I => \N__9309\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__9309\,
            I => \N__9306\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__9306\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9303\,
            I => \N__9300\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9300\,
            I => \N__9297\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__9297\,
            I => \N__9294\
        );

    \I__2013\ : Span4Mux_v
    port map (
            O => \N__9294\,
            I => \N__9291\
        );

    \I__2012\ : Span4Mux_v
    port map (
            O => \N__9291\,
            I => \N__9288\
        );

    \I__2011\ : Sp12to4
    port map (
            O => \N__9288\,
            I => \N__9285\
        );

    \I__2010\ : Span12Mux_h
    port map (
            O => \N__9285\,
            I => \N__9282\
        );

    \I__2009\ : Odrv12
    port map (
            O => \N__9282\,
            I => \A_c_14\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__9279\,
            I => \N__9276\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9276\,
            I => \N__9273\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__9273\,
            I => \N__9270\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__9270\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\
        );

    \I__2004\ : InMux
    port map (
            O => \N__9267\,
            I => \N__9264\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__9264\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__2002\ : InMux
    port map (
            O => \N__9261\,
            I => \N__9258\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9258\,
            I => \N__9255\
        );

    \I__2000\ : Span4Mux_h
    port map (
            O => \N__9255\,
            I => \N__9252\
        );

    \I__1999\ : Span4Mux_v
    port map (
            O => \N__9252\,
            I => \N__9249\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__9249\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9246\,
            I => \N__9243\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__9243\,
            I => \N__9240\
        );

    \I__1995\ : Span4Mux_h
    port map (
            O => \N__9240\,
            I => \N__9237\
        );

    \I__1994\ : Span4Mux_v
    port map (
            O => \N__9237\,
            I => \N__9234\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__9234\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1992\ : InMux
    port map (
            O => \N__9231\,
            I => \N__9228\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__9228\,
            I => \N__9225\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__9225\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1989\ : IoInMux
    port map (
            O => \N__9222\,
            I => \N__9219\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9219\,
            I => \N__9216\
        );

    \I__1987\ : Span12Mux_s0_v
    port map (
            O => \N__9216\,
            I => \N__9213\
        );

    \I__1986\ : Span12Mux_v
    port map (
            O => \N__9213\,
            I => \N__9210\
        );

    \I__1985\ : Odrv12
    port map (
            O => \N__9210\,
            I => \CMA_c_0\
        );

    \I__1984\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9204\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__9204\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\
        );

    \I__1982\ : InMux
    port map (
            O => \N__9201\,
            I => \N__9198\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__9198\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__9195\,
            I => \U712_CHIP_RAM.N_147_i_i_a2_0_cascade_\
        );

    \I__1979\ : CEMux
    port map (
            O => \N__9192\,
            I => \N__9189\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__9189\,
            I => \N__9185\
        );

    \I__1977\ : CEMux
    port map (
            O => \N__9188\,
            I => \N__9182\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__9185\,
            I => \N__9178\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__9182\,
            I => \N__9175\
        );

    \I__1974\ : CEMux
    port map (
            O => \N__9181\,
            I => \N__9172\
        );

    \I__1973\ : Span4Mux_h
    port map (
            O => \N__9178\,
            I => \N__9169\
        );

    \I__1972\ : Span4Mux_h
    port map (
            O => \N__9175\,
            I => \N__9166\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__9172\,
            I => \N__9163\
        );

    \I__1970\ : Odrv4
    port map (
            O => \N__9169\,
            I => \U712_CHIP_RAM.N_500_i\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__9166\,
            I => \U712_CHIP_RAM.N_500_i\
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__9163\,
            I => \U712_CHIP_RAM.N_500_i\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9156\,
            I => \N__9153\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__9153\,
            I => \N__9150\
        );

    \I__1965\ : Span4Mux_h
    port map (
            O => \N__9150\,
            I => \N__9146\
        );

    \I__1964\ : InMux
    port map (
            O => \N__9149\,
            I => \N__9143\
        );

    \I__1963\ : Span4Mux_h
    port map (
            O => \N__9146\,
            I => \N__9140\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__9143\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1961\ : Odrv4
    port map (
            O => \N__9140\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1960\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9132\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__9132\,
            I => \N__9129\
        );

    \I__1958\ : Span4Mux_h
    port map (
            O => \N__9129\,
            I => \N__9126\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__9126\,
            I => \U712_CHIP_RAM.REFRESH5lto7_0\
        );

    \I__1956\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9120\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__9120\,
            I => \N__9117\
        );

    \I__1954\ : Span4Mux_h
    port map (
            O => \N__9117\,
            I => \N__9114\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__9114\,
            I => \N__9111\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__9111\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__9108\,
            I => \N__9105\
        );

    \I__1950\ : InMux
    port map (
            O => \N__9105\,
            I => \N__9102\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__9102\,
            I => \N__9097\
        );

    \I__1948\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9093\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__9100\,
            I => \N__9089\
        );

    \I__1946\ : Span4Mux_h
    port map (
            O => \N__9097\,
            I => \N__9082\
        );

    \I__1945\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9079\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__9093\,
            I => \N__9076\
        );

    \I__1943\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9071\
        );

    \I__1942\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9071\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9068\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9087\,
            I => \N__9063\
        );

    \I__1939\ : InMux
    port map (
            O => \N__9086\,
            I => \N__9063\
        );

    \I__1938\ : InMux
    port map (
            O => \N__9085\,
            I => \N__9060\
        );

    \I__1937\ : Odrv4
    port map (
            O => \N__9082\,
            I => \U712_CHIP_RAM.N_509\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__9079\,
            I => \U712_CHIP_RAM.N_509\
        );

    \I__1935\ : Odrv12
    port map (
            O => \N__9076\,
            I => \U712_CHIP_RAM.N_509\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__9071\,
            I => \U712_CHIP_RAM.N_509\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__9068\,
            I => \U712_CHIP_RAM.N_509\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__9063\,
            I => \U712_CHIP_RAM.N_509\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__9060\,
            I => \U712_CHIP_RAM.N_509\
        );

    \I__1930\ : InMux
    port map (
            O => \N__9045\,
            I => \N__9037\
        );

    \I__1929\ : InMux
    port map (
            O => \N__9044\,
            I => \N__9037\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9043\,
            I => \N__9032\
        );

    \I__1927\ : InMux
    port map (
            O => \N__9042\,
            I => \N__9032\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__9037\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__9032\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1924\ : InMux
    port map (
            O => \N__9027\,
            I => \N__9022\
        );

    \I__1923\ : InMux
    port map (
            O => \N__9026\,
            I => \N__9019\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__9025\,
            I => \N__9012\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__9022\,
            I => \N__9007\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__9019\,
            I => \N__9004\
        );

    \I__1919\ : InMux
    port map (
            O => \N__9018\,
            I => \N__9001\
        );

    \I__1918\ : InMux
    port map (
            O => \N__9017\,
            I => \N__8998\
        );

    \I__1917\ : InMux
    port map (
            O => \N__9016\,
            I => \N__8991\
        );

    \I__1916\ : InMux
    port map (
            O => \N__9015\,
            I => \N__8991\
        );

    \I__1915\ : InMux
    port map (
            O => \N__9012\,
            I => \N__8991\
        );

    \I__1914\ : InMux
    port map (
            O => \N__9011\,
            I => \N__8986\
        );

    \I__1913\ : InMux
    port map (
            O => \N__9010\,
            I => \N__8986\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__9007\,
            I => \N__8979\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__9004\,
            I => \N__8979\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__9001\,
            I => \N__8979\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__8998\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8991\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8986\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__8979\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8966\
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__8969\,
            I => \N__8962\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__8966\,
            I => \N__8953\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8950\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8962\,
            I => \N__8947\
        );

    \I__1900\ : InMux
    port map (
            O => \N__8961\,
            I => \N__8944\
        );

    \I__1899\ : InMux
    port map (
            O => \N__8960\,
            I => \N__8939\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8959\,
            I => \N__8939\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8958\,
            I => \N__8932\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8957\,
            I => \N__8932\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8956\,
            I => \N__8932\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__8953\,
            I => \U712_CHIP_RAM.N_508\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__8950\,
            I => \U712_CHIP_RAM.N_508\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__8947\,
            I => \U712_CHIP_RAM.N_508\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__8944\,
            I => \U712_CHIP_RAM.N_508\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__8939\,
            I => \U712_CHIP_RAM.N_508\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8932\,
            I => \U712_CHIP_RAM.N_508\
        );

    \I__1888\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8916\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__8916\,
            I => \U712_CHIP_RAM.N_494\
        );

    \I__1886\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8910\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8910\,
            I => \N__8907\
        );

    \I__1884\ : Span4Mux_v
    port map (
            O => \N__8907\,
            I => \N__8904\
        );

    \I__1883\ : Sp12to4
    port map (
            O => \N__8904\,
            I => \N__8901\
        );

    \I__1882\ : Span12Mux_h
    port map (
            O => \N__8901\,
            I => \N__8898\
        );

    \I__1881\ : Span12Mux_h
    port map (
            O => \N__8898\,
            I => \N__8895\
        );

    \I__1880\ : Odrv12
    port map (
            O => \N__8895\,
            I => \A_c_12\
        );

    \I__1879\ : InMux
    port map (
            O => \N__8892\,
            I => \N__8889\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8889\,
            I => \N__8886\
        );

    \I__1877\ : Span12Mux_v
    port map (
            O => \N__8886\,
            I => \N__8883\
        );

    \I__1876\ : Span12Mux_h
    port map (
            O => \N__8883\,
            I => \N__8880\
        );

    \I__1875\ : Odrv12
    port map (
            O => \N__8880\,
            I => \A_c_13\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__8877\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8871\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8871\,
            I => \N__8868\
        );

    \I__1871\ : Span12Mux_v
    port map (
            O => \N__8868\,
            I => \N__8865\
        );

    \I__1870\ : Span12Mux_h
    port map (
            O => \N__8865\,
            I => \N__8862\
        );

    \I__1869\ : Odrv12
    port map (
            O => \N__8862\,
            I => \A_c_5\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8859\,
            I => \N__8856\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8856\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8853\,
            I => \N__8850\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8850\,
            I => \N__8847\
        );

    \I__1864\ : Span4Mux_h
    port map (
            O => \N__8847\,
            I => \N__8844\
        );

    \I__1863\ : Span4Mux_v
    port map (
            O => \N__8844\,
            I => \N__8841\
        );

    \I__1862\ : Sp12to4
    port map (
            O => \N__8841\,
            I => \N__8838\
        );

    \I__1861\ : Span12Mux_h
    port map (
            O => \N__8838\,
            I => \N__8835\
        );

    \I__1860\ : Odrv12
    port map (
            O => \N__8835\,
            I => \A_c_6\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8829\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8829\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\
        );

    \I__1857\ : CEMux
    port map (
            O => \N__8826\,
            I => \N__8821\
        );

    \I__1856\ : CEMux
    port map (
            O => \N__8825\,
            I => \N__8818\
        );

    \I__1855\ : CEMux
    port map (
            O => \N__8824\,
            I => \N__8815\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8821\,
            I => \N__8812\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8818\,
            I => \N__8809\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8815\,
            I => \N__8806\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__8812\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__1850\ : Odrv12
    port map (
            O => \N__8809\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__1849\ : Odrv4
    port map (
            O => \N__8806\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8799\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__8796\,
            I => \N__8793\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8793\,
            I => \N__8789\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8792\,
            I => \N__8786\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8789\,
            I => \N__8783\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__8786\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__8783\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8778\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8771\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8774\,
            I => \N__8768\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8771\,
            I => \N__8765\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8768\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1836\ : Odrv4
    port map (
            O => \N__8765\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8760\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8757\,
            I => \N__8751\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8746\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8755\,
            I => \N__8746\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8754\,
            I => \N__8739\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8751\,
            I => \N__8736\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__8746\,
            I => \N__8733\
        );

    \I__1828\ : InMux
    port map (
            O => \N__8745\,
            I => \N__8724\
        );

    \I__1827\ : InMux
    port map (
            O => \N__8744\,
            I => \N__8724\
        );

    \I__1826\ : InMux
    port map (
            O => \N__8743\,
            I => \N__8724\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8742\,
            I => \N__8724\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8739\,
            I => \N__8721\
        );

    \I__1823\ : Span4Mux_v
    port map (
            O => \N__8736\,
            I => \N__8718\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__8733\,
            I => \U712_CHIP_RAM.N_132_i\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8724\,
            I => \U712_CHIP_RAM.N_132_i\
        );

    \I__1820\ : Odrv4
    port map (
            O => \N__8721\,
            I => \U712_CHIP_RAM.N_132_i\
        );

    \I__1819\ : Odrv4
    port map (
            O => \N__8718\,
            I => \U712_CHIP_RAM.N_132_i\
        );

    \I__1818\ : InMux
    port map (
            O => \N__8709\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8702\
        );

    \I__1816\ : InMux
    port map (
            O => \N__8705\,
            I => \N__8699\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__8702\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8699\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8685\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8678\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8692\,
            I => \N__8678\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8691\,
            I => \N__8678\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8690\,
            I => \N__8671\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8689\,
            I => \N__8671\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8688\,
            I => \N__8671\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8685\,
            I => \N__8668\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__8678\,
            I => \N__8663\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8671\,
            I => \N__8663\
        );

    \I__1803\ : Span4Mux_v
    port map (
            O => \N__8668\,
            I => \N__8660\
        );

    \I__1802\ : Span4Mux_h
    port map (
            O => \N__8663\,
            I => \N__8657\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__8660\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1800\ : Odrv4
    port map (
            O => \N__8657\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__8652\,
            I => \N__8648\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8643\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8640\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8647\,
            I => \N__8637\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8646\,
            I => \N__8634\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__8643\,
            I => \N__8628\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8640\,
            I => \N__8628\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__8637\,
            I => \N__8617\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__8634\,
            I => \N__8617\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8612\
        );

    \I__1789\ : Span4Mux_v
    port map (
            O => \N__8628\,
            I => \N__8609\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8627\,
            I => \N__8606\
        );

    \I__1787\ : InMux
    port map (
            O => \N__8626\,
            I => \N__8603\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8596\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8596\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8623\,
            I => \N__8596\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8622\,
            I => \N__8593\
        );

    \I__1782\ : Span4Mux_h
    port map (
            O => \N__8617\,
            I => \N__8590\
        );

    \I__1781\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8585\
        );

    \I__1780\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8585\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8612\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__8609\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__8606\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8603\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8596\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__8593\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__8590\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8585\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8565\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8565\,
            I => \U712_CHIP_RAM.N_436\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8559\,
            I => \N__8556\
        );

    \I__1767\ : Span4Mux_v
    port map (
            O => \N__8556\,
            I => \N__8553\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__8553\,
            I => \U712_CHIP_RAM.N_499\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8542\
        );

    \I__1764\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8542\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8538\
        );

    \I__1762\ : InMux
    port map (
            O => \N__8547\,
            I => \N__8535\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__8542\,
            I => \N__8532\
        );

    \I__1760\ : InMux
    port map (
            O => \N__8541\,
            I => \N__8529\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__8538\,
            I => \N__8526\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__8535\,
            I => \N__8523\
        );

    \I__1757\ : Span4Mux_v
    port map (
            O => \N__8532\,
            I => \N__8516\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8529\,
            I => \N__8516\
        );

    \I__1755\ : Span4Mux_h
    port map (
            O => \N__8526\,
            I => \N__8511\
        );

    \I__1754\ : Span4Mux_h
    port map (
            O => \N__8523\,
            I => \N__8511\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8508\
        );

    \I__1752\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8505\
        );

    \I__1751\ : Span4Mux_h
    port map (
            O => \N__8516\,
            I => \N__8502\
        );

    \I__1750\ : Span4Mux_v
    port map (
            O => \N__8511\,
            I => \N__8499\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__8508\,
            I => \N__8494\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8505\,
            I => \N__8494\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__8502\,
            I => \DMA_CYCLEm\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__8499\,
            I => \DMA_CYCLEm\
        );

    \I__1745\ : Odrv12
    port map (
            O => \N__8494\,
            I => \DMA_CYCLEm\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8487\,
            I => \N__8477\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8477\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8485\,
            I => \N__8477\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8484\,
            I => \N__8474\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8477\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8474\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__8469\,
            I => \N__8464\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__8468\,
            I => \N__8461\
        );

    \I__1736\ : InMux
    port map (
            O => \N__8467\,
            I => \N__8458\
        );

    \I__1735\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8453\
        );

    \I__1734\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8453\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8458\,
            I => \N__8450\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8453\,
            I => \N__8447\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__8450\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__1730\ : Odrv12
    port map (
            O => \N__8447\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\
        );

    \I__1729\ : InMux
    port map (
            O => \N__8442\,
            I => \N__8431\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8441\,
            I => \N__8427\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8440\,
            I => \N__8418\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8439\,
            I => \N__8418\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8410\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8410\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8436\,
            I => \N__8410\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__8435\,
            I => \N__8406\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__8434\,
            I => \N__8397\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8431\,
            I => \N__8394\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8391\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__8427\,
            I => \N__8388\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__8426\,
            I => \N__8385\
        );

    \I__1716\ : InMux
    port map (
            O => \N__8425\,
            I => \N__8379\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8379\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8423\,
            I => \N__8376\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__8418\,
            I => \N__8373\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__8417\,
            I => \N__8368\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__8410\,
            I => \N__8365\
        );

    \I__1710\ : InMux
    port map (
            O => \N__8409\,
            I => \N__8358\
        );

    \I__1709\ : InMux
    port map (
            O => \N__8406\,
            I => \N__8358\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8405\,
            I => \N__8358\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8351\
        );

    \I__1706\ : InMux
    port map (
            O => \N__8403\,
            I => \N__8351\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8402\,
            I => \N__8351\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__8401\,
            I => \N__8348\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8400\,
            I => \N__8343\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8397\,
            I => \N__8340\
        );

    \I__1701\ : Span4Mux_v
    port map (
            O => \N__8394\,
            I => \N__8333\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8391\,
            I => \N__8333\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__8388\,
            I => \N__8333\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8385\,
            I => \N__8328\
        );

    \I__1697\ : InMux
    port map (
            O => \N__8384\,
            I => \N__8328\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__8379\,
            I => \N__8321\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8376\,
            I => \N__8321\
        );

    \I__1694\ : Span4Mux_h
    port map (
            O => \N__8373\,
            I => \N__8321\
        );

    \I__1693\ : InMux
    port map (
            O => \N__8372\,
            I => \N__8314\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8314\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8368\,
            I => \N__8314\
        );

    \I__1690\ : Span4Mux_h
    port map (
            O => \N__8365\,
            I => \N__8307\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8358\,
            I => \N__8307\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8351\,
            I => \N__8307\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8300\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8300\
        );

    \I__1685\ : InMux
    port map (
            O => \N__8346\,
            I => \N__8300\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__8343\,
            I => \N__8297\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8340\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__8333\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__8328\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__8321\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8314\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__8307\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__8300\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__8297\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__8280\,
            I => \U712_CHIP_RAM.N_506_cascade_\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8274\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__8274\,
            I => \U712_CHIP_RAM.N_147_i_i_a2_0\
        );

    \I__1672\ : InMux
    port map (
            O => \N__8271\,
            I => \N__8268\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__8268\,
            I => \N__8265\
        );

    \I__1670\ : Span4Mux_h
    port map (
            O => \N__8265\,
            I => \N__8261\
        );

    \I__1669\ : InMux
    port map (
            O => \N__8264\,
            I => \N__8258\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__8261\,
            I => \U712_CHIP_RAM.N_359\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__8258\,
            I => \U712_CHIP_RAM.N_359\
        );

    \I__1666\ : InMux
    port map (
            O => \N__8253\,
            I => \N__8250\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8250\,
            I => \U712_CHIP_RAM.N_595\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__8247\,
            I => \N__8244\
        );

    \I__1663\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8240\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8243\,
            I => \N__8236\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__8240\,
            I => \N__8232\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8239\,
            I => \N__8229\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__8236\,
            I => \N__8226\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__8235\,
            I => \N__8223\
        );

    \I__1657\ : Span4Mux_h
    port map (
            O => \N__8232\,
            I => \N__8218\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__8229\,
            I => \N__8218\
        );

    \I__1655\ : Span4Mux_h
    port map (
            O => \N__8226\,
            I => \N__8215\
        );

    \I__1654\ : InMux
    port map (
            O => \N__8223\,
            I => \N__8212\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__8218\,
            I => \U712_CHIP_RAM.N_348\
        );

    \I__1652\ : Odrv4
    port map (
            O => \N__8215\,
            I => \U712_CHIP_RAM.N_348\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8212\,
            I => \U712_CHIP_RAM.N_348\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__8205\,
            I => \U712_CHIP_RAM.N_595_cascade_\
        );

    \I__1649\ : InMux
    port map (
            O => \N__8202\,
            I => \N__8196\
        );

    \I__1648\ : InMux
    port map (
            O => \N__8201\,
            I => \N__8191\
        );

    \I__1647\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8191\
        );

    \I__1646\ : InMux
    port map (
            O => \N__8199\,
            I => \N__8188\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__8196\,
            I => \U712_CHIP_RAM.N_577\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__8191\,
            I => \U712_CHIP_RAM.N_577\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__8188\,
            I => \U712_CHIP_RAM.N_577\
        );

    \I__1642\ : InMux
    port map (
            O => \N__8181\,
            I => \N__8178\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__8178\,
            I => \N__8175\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__8175\,
            I => \U712_CHIP_RAM.N_279\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__8172\,
            I => \N__8168\
        );

    \I__1638\ : InMux
    port map (
            O => \N__8171\,
            I => \N__8158\
        );

    \I__1637\ : InMux
    port map (
            O => \N__8168\,
            I => \N__8153\
        );

    \I__1636\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8153\
        );

    \I__1635\ : InMux
    port map (
            O => \N__8166\,
            I => \N__8150\
        );

    \I__1634\ : InMux
    port map (
            O => \N__8165\,
            I => \N__8147\
        );

    \I__1633\ : InMux
    port map (
            O => \N__8164\,
            I => \N__8142\
        );

    \I__1632\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8142\
        );

    \I__1631\ : InMux
    port map (
            O => \N__8162\,
            I => \N__8137\
        );

    \I__1630\ : InMux
    port map (
            O => \N__8161\,
            I => \N__8137\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__8158\,
            I => \N__8130\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__8153\,
            I => \N__8130\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__8150\,
            I => \N__8130\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__8147\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__8142\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__8137\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__8130\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1622\ : InMux
    port map (
            O => \N__8121\,
            I => \N__8118\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__8118\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_i_a2_0_1\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__8115\,
            I => \N__8107\
        );

    \I__1619\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8100\
        );

    \I__1618\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8100\
        );

    \I__1617\ : CascadeMux
    port map (
            O => \N__8112\,
            I => \N__8095\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8111\,
            I => \N__8085\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8110\,
            I => \N__8085\
        );

    \I__1614\ : InMux
    port map (
            O => \N__8107\,
            I => \N__8085\
        );

    \I__1613\ : InMux
    port map (
            O => \N__8106\,
            I => \N__8085\
        );

    \I__1612\ : InMux
    port map (
            O => \N__8105\,
            I => \N__8076\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__8100\,
            I => \N__8073\
        );

    \I__1610\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8064\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8098\,
            I => \N__8064\
        );

    \I__1608\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8064\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8094\,
            I => \N__8064\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__8085\,
            I => \N__8061\
        );

    \I__1605\ : InMux
    port map (
            O => \N__8084\,
            I => \N__8056\
        );

    \I__1604\ : InMux
    port map (
            O => \N__8083\,
            I => \N__8056\
        );

    \I__1603\ : InMux
    port map (
            O => \N__8082\,
            I => \N__8051\
        );

    \I__1602\ : InMux
    port map (
            O => \N__8081\,
            I => \N__8051\
        );

    \I__1601\ : InMux
    port map (
            O => \N__8080\,
            I => \N__8048\
        );

    \I__1600\ : InMux
    port map (
            O => \N__8079\,
            I => \N__8045\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__8076\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1598\ : Odrv4
    port map (
            O => \N__8073\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__8064\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__8061\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__8056\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__8051\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__8048\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__8045\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1591\ : InMux
    port map (
            O => \N__8028\,
            I => \N__8024\
        );

    \I__1590\ : InMux
    port map (
            O => \N__8027\,
            I => \N__8021\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__8024\,
            I => \N__8018\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__8021\,
            I => \N__8015\
        );

    \I__1587\ : Span4Mux_v
    port map (
            O => \N__8018\,
            I => \N__8010\
        );

    \I__1586\ : Span4Mux_h
    port map (
            O => \N__8015\,
            I => \N__8010\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__8010\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0\
        );

    \I__1584\ : InMux
    port map (
            O => \N__8007\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__1583\ : InMux
    port map (
            O => \N__8004\,
            I => \N__8001\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__8001\,
            I => \N__7998\
        );

    \I__1581\ : Span12Mux_h
    port map (
            O => \N__7998\,
            I => \N__7995\
        );

    \I__1580\ : Odrv12
    port map (
            O => \N__7995\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7992\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__7989\,
            I => \N__7985\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__7988\,
            I => \N__7981\
        );

    \I__1576\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7978\
        );

    \I__1575\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7975\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7971\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7978\,
            I => \N__7966\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__7975\,
            I => \N__7963\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__7974\,
            I => \N__7958\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__7971\,
            I => \N__7954\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7951\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7947\
        );

    \I__1567\ : Span4Mux_h
    port map (
            O => \N__7966\,
            I => \N__7942\
        );

    \I__1566\ : Span4Mux_v
    port map (
            O => \N__7963\,
            I => \N__7942\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7937\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7937\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7932\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7957\,
            I => \N__7932\
        );

    \I__1561\ : Span4Mux_v
    port map (
            O => \N__7954\,
            I => \N__7927\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__7951\,
            I => \N__7927\
        );

    \I__1559\ : InMux
    port map (
            O => \N__7950\,
            I => \N__7924\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7947\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1557\ : Odrv4
    port map (
            O => \N__7942\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7937\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7932\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__7927\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__7924\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7911\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7904\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7907\,
            I => \N__7901\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7904\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__7901\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__7896\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_\
        );

    \I__1546\ : IoInMux
    port map (
            O => \N__7893\,
            I => \N__7890\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7890\,
            I => \N__7887\
        );

    \I__1544\ : Span12Mux_s9_v
    port map (
            O => \N__7887\,
            I => \N__7884\
        );

    \I__1543\ : Span12Mux_h
    port map (
            O => \N__7884\,
            I => \N__7880\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7877\
        );

    \I__1541\ : Odrv12
    port map (
            O => \N__7880\,
            I => \LATCH_CLK_c\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7877\,
            I => \LATCH_CLK_c\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7872\,
            I => \N__7869\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7869\,
            I => \N__7866\
        );

    \I__1537\ : Span12Mux_h
    port map (
            O => \N__7866\,
            I => \N__7863\
        );

    \I__1536\ : Odrv12
    port map (
            O => \N__7863\,
            I => \DBRn_c_i\
        );

    \I__1535\ : InMux
    port map (
            O => \N__7860\,
            I => \N__7857\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7857\,
            I => \N__7854\
        );

    \I__1533\ : Span4Mux_h
    port map (
            O => \N__7854\,
            I => \N__7850\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7853\,
            I => \N__7847\
        );

    \I__1531\ : Span4Mux_v
    port map (
            O => \N__7850\,
            I => \N__7844\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__7847\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1529\ : Odrv4
    port map (
            O => \N__7844\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1528\ : IoInMux
    port map (
            O => \N__7839\,
            I => \N__7836\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7836\,
            I => \N__7833\
        );

    \I__1526\ : Span12Mux_s6_v
    port map (
            O => \N__7833\,
            I => \N__7830\
        );

    \I__1525\ : Odrv12
    port map (
            O => \N__7830\,
            I => \N_119_i\
        );

    \I__1524\ : InMux
    port map (
            O => \N__7827\,
            I => \N__7821\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7826\,
            I => \N__7818\
        );

    \I__1522\ : InMux
    port map (
            O => \N__7825\,
            I => \N__7813\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7824\,
            I => \N__7813\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7821\,
            I => \N__7810\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7818\,
            I => \N__7807\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7813\,
            I => \N__7804\
        );

    \I__1517\ : Span4Mux_v
    port map (
            O => \N__7810\,
            I => \N__7797\
        );

    \I__1516\ : Span4Mux_h
    port map (
            O => \N__7807\,
            I => \N__7792\
        );

    \I__1515\ : Span4Mux_v
    port map (
            O => \N__7804\,
            I => \N__7792\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7803\,
            I => \N__7787\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7802\,
            I => \N__7787\
        );

    \I__1512\ : InMux
    port map (
            O => \N__7801\,
            I => \N__7782\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7782\
        );

    \I__1510\ : Span4Mux_v
    port map (
            O => \N__7797\,
            I => \N__7779\
        );

    \I__1509\ : Span4Mux_v
    port map (
            O => \N__7792\,
            I => \N__7776\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__7787\,
            I => \N__7771\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__7782\,
            I => \N__7771\
        );

    \I__1506\ : Span4Mux_v
    port map (
            O => \N__7779\,
            I => \N__7768\
        );

    \I__1505\ : Span4Mux_v
    port map (
            O => \N__7776\,
            I => \N__7763\
        );

    \I__1504\ : Span4Mux_v
    port map (
            O => \N__7771\,
            I => \N__7763\
        );

    \I__1503\ : Sp12to4
    port map (
            O => \N__7768\,
            I => \N__7758\
        );

    \I__1502\ : Sp12to4
    port map (
            O => \N__7763\,
            I => \N__7758\
        );

    \I__1501\ : Span12Mux_h
    port map (
            O => \N__7758\,
            I => \N__7755\
        );

    \I__1500\ : Odrv12
    port map (
            O => \N__7755\,
            I => \A_c_1\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__7752\,
            I => \N__7745\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7751\,
            I => \N__7740\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7740\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__7749\,
            I => \N__7737\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7748\,
            I => \N__7733\
        );

    \I__1494\ : InMux
    port map (
            O => \N__7745\,
            I => \N__7727\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__7740\,
            I => \N__7724\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7737\,
            I => \N__7719\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7736\,
            I => \N__7719\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__7733\,
            I => \N__7716\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7732\,
            I => \N__7713\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7731\,
            I => \N__7710\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7730\,
            I => \N__7707\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7727\,
            I => \N__7704\
        );

    \I__1485\ : Span4Mux_v
    port map (
            O => \N__7724\,
            I => \N__7699\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__7719\,
            I => \N__7699\
        );

    \I__1483\ : Span4Mux_v
    port map (
            O => \N__7716\,
            I => \N__7692\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__7713\,
            I => \N__7692\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7710\,
            I => \N__7692\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7707\,
            I => \N__7689\
        );

    \I__1479\ : Span4Mux_v
    port map (
            O => \N__7704\,
            I => \N__7686\
        );

    \I__1478\ : Span4Mux_h
    port map (
            O => \N__7699\,
            I => \N__7683\
        );

    \I__1477\ : Span4Mux_h
    port map (
            O => \N__7692\,
            I => \N__7678\
        );

    \I__1476\ : Span4Mux_v
    port map (
            O => \N__7689\,
            I => \N__7678\
        );

    \I__1475\ : Span4Mux_v
    port map (
            O => \N__7686\,
            I => \N__7675\
        );

    \I__1474\ : Span4Mux_v
    port map (
            O => \N__7683\,
            I => \N__7670\
        );

    \I__1473\ : Span4Mux_v
    port map (
            O => \N__7678\,
            I => \N__7670\
        );

    \I__1472\ : Sp12to4
    port map (
            O => \N__7675\,
            I => \N__7665\
        );

    \I__1471\ : Sp12to4
    port map (
            O => \N__7670\,
            I => \N__7665\
        );

    \I__1470\ : Span12Mux_h
    port map (
            O => \N__7665\,
            I => \N__7662\
        );

    \I__1469\ : Odrv12
    port map (
            O => \N__7662\,
            I => \A_c_0\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__7659\,
            I => \N__7655\
        );

    \I__1467\ : CascadeMux
    port map (
            O => \N__7658\,
            I => \N__7652\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7655\,
            I => \N__7647\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7652\,
            I => \N__7642\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7651\,
            I => \N__7642\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__7650\,
            I => \N__7638\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__7647\,
            I => \N__7635\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__7642\,
            I => \N__7630\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7641\,
            I => \N__7625\
        );

    \I__1459\ : InMux
    port map (
            O => \N__7638\,
            I => \N__7625\
        );

    \I__1458\ : Span4Mux_v
    port map (
            O => \N__7635\,
            I => \N__7622\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7634\,
            I => \N__7619\
        );

    \I__1456\ : InMux
    port map (
            O => \N__7633\,
            I => \N__7616\
        );

    \I__1455\ : Span4Mux_h
    port map (
            O => \N__7630\,
            I => \N__7610\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7625\,
            I => \N__7610\
        );

    \I__1453\ : Span4Mux_h
    port map (
            O => \N__7622\,
            I => \N__7607\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7619\,
            I => \N__7604\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7616\,
            I => \N__7601\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7615\,
            I => \N__7598\
        );

    \I__1449\ : Span4Mux_h
    port map (
            O => \N__7610\,
            I => \N__7595\
        );

    \I__1448\ : Sp12to4
    port map (
            O => \N__7607\,
            I => \N__7586\
        );

    \I__1447\ : Span12Mux_h
    port map (
            O => \N__7604\,
            I => \N__7586\
        );

    \I__1446\ : Sp12to4
    port map (
            O => \N__7601\,
            I => \N__7586\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7598\,
            I => \N__7586\
        );

    \I__1444\ : Span4Mux_v
    port map (
            O => \N__7595\,
            I => \N__7583\
        );

    \I__1443\ : Span12Mux_h
    port map (
            O => \N__7586\,
            I => \N__7580\
        );

    \I__1442\ : Span4Mux_h
    port map (
            O => \N__7583\,
            I => \N__7577\
        );

    \I__1441\ : Span12Mux_v
    port map (
            O => \N__7580\,
            I => \N__7574\
        );

    \I__1440\ : Sp12to4
    port map (
            O => \N__7577\,
            I => \N__7571\
        );

    \I__1439\ : Odrv12
    port map (
            O => \N__7574\,
            I => \SIZ_c_0\
        );

    \I__1438\ : Odrv12
    port map (
            O => \N__7571\,
            I => \SIZ_c_0\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__7566\,
            I => \N__7562\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7554\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7562\,
            I => \N__7554\
        );

    \I__1434\ : InMux
    port map (
            O => \N__7561\,
            I => \N__7550\
        );

    \I__1433\ : CascadeMux
    port map (
            O => \N__7560\,
            I => \N__7547\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__7559\,
            I => \N__7544\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__7554\,
            I => \N__7540\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7553\,
            I => \N__7537\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7550\,
            I => \N__7532\
        );

    \I__1428\ : InMux
    port map (
            O => \N__7547\,
            I => \N__7529\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7544\,
            I => \N__7526\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7543\,
            I => \N__7523\
        );

    \I__1425\ : Span4Mux_h
    port map (
            O => \N__7540\,
            I => \N__7520\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__7537\,
            I => \N__7517\
        );

    \I__1423\ : InMux
    port map (
            O => \N__7536\,
            I => \N__7512\
        );

    \I__1422\ : InMux
    port map (
            O => \N__7535\,
            I => \N__7512\
        );

    \I__1421\ : Sp12to4
    port map (
            O => \N__7532\,
            I => \N__7509\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7529\,
            I => \N__7502\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__7526\,
            I => \N__7502\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__7523\,
            I => \N__7502\
        );

    \I__1417\ : Span4Mux_v
    port map (
            O => \N__7520\,
            I => \N__7499\
        );

    \I__1416\ : Span12Mux_v
    port map (
            O => \N__7517\,
            I => \N__7494\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__7512\,
            I => \N__7494\
        );

    \I__1414\ : Span12Mux_v
    port map (
            O => \N__7509\,
            I => \N__7491\
        );

    \I__1413\ : Span12Mux_h
    port map (
            O => \N__7502\,
            I => \N__7488\
        );

    \I__1412\ : Sp12to4
    port map (
            O => \N__7499\,
            I => \N__7483\
        );

    \I__1411\ : Span12Mux_v
    port map (
            O => \N__7494\,
            I => \N__7483\
        );

    \I__1410\ : Span12Mux_h
    port map (
            O => \N__7491\,
            I => \N__7480\
        );

    \I__1409\ : Span12Mux_v
    port map (
            O => \N__7488\,
            I => \N__7477\
        );

    \I__1408\ : Span12Mux_h
    port map (
            O => \N__7483\,
            I => \N__7474\
        );

    \I__1407\ : Odrv12
    port map (
            O => \N__7480\,
            I => \SIZ_c_1\
        );

    \I__1406\ : Odrv12
    port map (
            O => \N__7477\,
            I => \SIZ_c_1\
        );

    \I__1405\ : Odrv12
    port map (
            O => \N__7474\,
            I => \SIZ_c_1\
        );

    \I__1404\ : IoInMux
    port map (
            O => \N__7467\,
            I => \N__7464\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7464\,
            I => \N__7461\
        );

    \I__1402\ : Span4Mux_s3_v
    port map (
            O => \N__7461\,
            I => \N__7458\
        );

    \I__1401\ : Odrv4
    port map (
            O => \N__7458\,
            I => \N_61_i\
        );

    \I__1400\ : IoInMux
    port map (
            O => \N__7455\,
            I => \N__7452\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7452\,
            I => \N__7449\
        );

    \I__1398\ : Span4Mux_s0_v
    port map (
            O => \N__7449\,
            I => \N__7446\
        );

    \I__1397\ : Span4Mux_v
    port map (
            O => \N__7446\,
            I => \N__7443\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__7443\,
            I => \N__7440\
        );

    \I__1395\ : Span4Mux_h
    port map (
            O => \N__7440\,
            I => \N__7437\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__7437\,
            I => \CMA_c_2\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7434\,
            I => \N__7431\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7431\,
            I => \N__7428\
        );

    \I__1391\ : Span4Mux_v
    port map (
            O => \N__7428\,
            I => \N__7425\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__7425\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1389\ : InMux
    port map (
            O => \N__7422\,
            I => \N__7419\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__7419\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1387\ : IoInMux
    port map (
            O => \N__7416\,
            I => \N__7412\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7415\,
            I => \N__7409\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7412\,
            I => \N__7406\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__7409\,
            I => \N__7403\
        );

    \I__1383\ : Span4Mux_s3_v
    port map (
            O => \N__7406\,
            I => \N__7400\
        );

    \I__1382\ : Span4Mux_v
    port map (
            O => \N__7403\,
            I => \N__7397\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__7400\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__7397\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__7392\,
            I => \N__7389\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7389\,
            I => \N__7386\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7386\,
            I => \N__7383\
        );

    \I__1376\ : Span4Mux_h
    port map (
            O => \N__7383\,
            I => \N__7380\
        );

    \I__1375\ : Odrv4
    port map (
            O => \N__7380\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7377\,
            I => \N__7374\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7374\,
            I => \U712_CHIP_RAM.N_431\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7371\,
            I => \N__7368\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7368\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7365\,
            I => \N__7362\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__7362\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\
        );

    \I__1368\ : IoInMux
    port map (
            O => \N__7359\,
            I => \N__7356\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7356\,
            I => \N__7353\
        );

    \I__1366\ : IoSpan4Mux
    port map (
            O => \N__7353\,
            I => \N__7350\
        );

    \I__1365\ : Span4Mux_s2_v
    port map (
            O => \N__7350\,
            I => \N__7346\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7349\,
            I => \N__7343\
        );

    \I__1363\ : Sp12to4
    port map (
            O => \N__7346\,
            I => \N__7340\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__7343\,
            I => \N__7337\
        );

    \I__1361\ : Span12Mux_s8_v
    port map (
            O => \N__7340\,
            I => \N__7334\
        );

    \I__1360\ : Sp12to4
    port map (
            O => \N__7337\,
            I => \N__7331\
        );

    \I__1359\ : Span12Mux_h
    port map (
            O => \N__7334\,
            I => \N__7328\
        );

    \I__1358\ : Span12Mux_v
    port map (
            O => \N__7331\,
            I => \N__7325\
        );

    \I__1357\ : Span12Mux_v
    port map (
            O => \N__7328\,
            I => \N__7322\
        );

    \I__1356\ : Span12Mux_h
    port map (
            O => \N__7325\,
            I => \N__7319\
        );

    \I__1355\ : Odrv12
    port map (
            O => \N__7322\,
            I => \A_c_11\
        );

    \I__1354\ : Odrv12
    port map (
            O => \N__7319\,
            I => \A_c_11\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7314\,
            I => \N__7310\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7313\,
            I => \N__7307\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7310\,
            I => \U712_CHIP_RAM.N_350\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__7307\,
            I => \U712_CHIP_RAM.N_350\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7302\,
            I => \N__7299\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__7299\,
            I => \U712_CHIP_RAM.N_452\
        );

    \I__1347\ : IoInMux
    port map (
            O => \N__7296\,
            I => \N__7292\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7295\,
            I => \N__7289\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__7292\,
            I => \N__7286\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7289\,
            I => \N__7283\
        );

    \I__1343\ : Span12Mux_s4_v
    port map (
            O => \N__7286\,
            I => \N__7280\
        );

    \I__1342\ : Span4Mux_v
    port map (
            O => \N__7283\,
            I => \N__7277\
        );

    \I__1341\ : Span12Mux_v
    port map (
            O => \N__7280\,
            I => \N__7274\
        );

    \I__1340\ : Sp12to4
    port map (
            O => \N__7277\,
            I => \N__7271\
        );

    \I__1339\ : Span12Mux_h
    port map (
            O => \N__7274\,
            I => \N__7268\
        );

    \I__1338\ : Span12Mux_h
    port map (
            O => \N__7271\,
            I => \N__7265\
        );

    \I__1337\ : Odrv12
    port map (
            O => \N__7268\,
            I => \A_c_9\
        );

    \I__1336\ : Odrv12
    port map (
            O => \N__7265\,
            I => \A_c_9\
        );

    \I__1335\ : InMux
    port map (
            O => \N__7260\,
            I => \N__7257\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7257\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__7254\,
            I => \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a2_1_cascade_\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7251\,
            I => \N__7245\
        );

    \I__1331\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7242\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__7249\,
            I => \N__7239\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__7248\,
            I => \N__7235\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__7245\,
            I => \N__7230\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__7242\,
            I => \N__7227\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7239\,
            I => \N__7222\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7222\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7217\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7234\,
            I => \N__7217\
        );

    \I__1322\ : InMux
    port map (
            O => \N__7233\,
            I => \N__7214\
        );

    \I__1321\ : Odrv12
    port map (
            O => \N__7230\,
            I => \U712_CHIP_RAM.N_344\
        );

    \I__1320\ : Odrv4
    port map (
            O => \N__7227\,
            I => \U712_CHIP_RAM.N_344\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__7222\,
            I => \U712_CHIP_RAM.N_344\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__7217\,
            I => \U712_CHIP_RAM.N_344\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__7214\,
            I => \U712_CHIP_RAM.N_344\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7203\,
            I => \N__7200\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__7200\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_0\
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__7197\,
            I => \U712_CHIP_RAM.N_72_cascade_\
        );

    \I__1313\ : InMux
    port map (
            O => \N__7194\,
            I => \N__7191\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__7191\,
            I => \N__7188\
        );

    \I__1311\ : Span4Mux_h
    port map (
            O => \N__7188\,
            I => \N__7184\
        );

    \I__1310\ : InMux
    port map (
            O => \N__7187\,
            I => \N__7181\
        );

    \I__1309\ : Odrv4
    port map (
            O => \N__7184\,
            I => \CPU_TACKm\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__7181\,
            I => \CPU_TACKm\
        );

    \I__1307\ : InMux
    port map (
            O => \N__7176\,
            I => \N__7173\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__7173\,
            I => \U712_CHIP_RAM.N_462\
        );

    \I__1305\ : InMux
    port map (
            O => \N__7170\,
            I => \N__7164\
        );

    \I__1304\ : InMux
    port map (
            O => \N__7169\,
            I => \N__7159\
        );

    \I__1303\ : InMux
    port map (
            O => \N__7168\,
            I => \N__7159\
        );

    \I__1302\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7155\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__7164\,
            I => \N__7152\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7159\,
            I => \N__7149\
        );

    \I__1299\ : InMux
    port map (
            O => \N__7158\,
            I => \N__7146\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__7155\,
            I => \N__7142\
        );

    \I__1297\ : Span4Mux_v
    port map (
            O => \N__7152\,
            I => \N__7134\
        );

    \I__1296\ : Span4Mux_v
    port map (
            O => \N__7149\,
            I => \N__7134\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__7146\,
            I => \N__7131\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7128\
        );

    \I__1293\ : Span4Mux_h
    port map (
            O => \N__7142\,
            I => \N__7125\
        );

    \I__1292\ : InMux
    port map (
            O => \N__7141\,
            I => \N__7118\
        );

    \I__1291\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7118\
        );

    \I__1290\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7118\
        );

    \I__1289\ : Odrv4
    port map (
            O => \N__7134\,
            I => \U712_CHIP_RAM.N_503\
        );

    \I__1288\ : Odrv12
    port map (
            O => \N__7131\,
            I => \U712_CHIP_RAM.N_503\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__7128\,
            I => \U712_CHIP_RAM.N_503\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__7125\,
            I => \U712_CHIP_RAM.N_503\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__7118\,
            I => \U712_CHIP_RAM.N_503\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__7107\,
            I => \U712_CHIP_RAM.N_462_cascade_\
        );

    \I__1283\ : InMux
    port map (
            O => \N__7104\,
            I => \N__7095\
        );

    \I__1282\ : InMux
    port map (
            O => \N__7103\,
            I => \N__7095\
        );

    \I__1281\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7090\
        );

    \I__1280\ : InMux
    port map (
            O => \N__7101\,
            I => \N__7090\
        );

    \I__1279\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7085\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__7095\,
            I => \N__7082\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__7090\,
            I => \N__7079\
        );

    \I__1276\ : InMux
    port map (
            O => \N__7089\,
            I => \N__7074\
        );

    \I__1275\ : InMux
    port map (
            O => \N__7088\,
            I => \N__7074\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__7085\,
            I => \U712_CHIP_RAM.N_510\
        );

    \I__1273\ : Odrv12
    port map (
            O => \N__7082\,
            I => \U712_CHIP_RAM.N_510\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__7079\,
            I => \U712_CHIP_RAM.N_510\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__7074\,
            I => \U712_CHIP_RAM.N_510\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__7065\,
            I => \U712_CHIP_RAM.N_347_cascade_\
        );

    \I__1269\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7059\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__7059\,
            I => \U712_CHIP_RAM.N_590\
        );

    \I__1267\ : CascadeMux
    port map (
            O => \N__7056\,
            I => \U712_CHIP_RAM.N_590_cascade_\
        );

    \I__1266\ : InMux
    port map (
            O => \N__7053\,
            I => \N__7050\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__7050\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0\
        );

    \I__1264\ : InMux
    port map (
            O => \N__7047\,
            I => \N__7043\
        );

    \I__1263\ : InMux
    port map (
            O => \N__7046\,
            I => \N__7040\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__7043\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__7040\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__7035\,
            I => \U712_CHIP_RAM.N_509_cascade_\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__7032\,
            I => \N__7029\
        );

    \I__1258\ : InMux
    port map (
            O => \N__7029\,
            I => \N__7026\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__7026\,
            I => \N__7023\
        );

    \I__1256\ : Span4Mux_h
    port map (
            O => \N__7023\,
            I => \N__7020\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__7020\,
            I => \U712_CHIP_RAM.DBENn_8_0_0\
        );

    \I__1254\ : InMux
    port map (
            O => \N__7017\,
            I => \N__7014\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__7014\,
            I => \N__7010\
        );

    \I__1252\ : InMux
    port map (
            O => \N__7013\,
            I => \N__7007\
        );

    \I__1251\ : Span4Mux_v
    port map (
            O => \N__7010\,
            I => \N__7004\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__7007\,
            I => \N__7001\
        );

    \I__1249\ : Sp12to4
    port map (
            O => \N__7004\,
            I => \N__6998\
        );

    \I__1248\ : Span12Mux_v
    port map (
            O => \N__7001\,
            I => \N__6995\
        );

    \I__1247\ : Span12Mux_h
    port map (
            O => \N__6998\,
            I => \N__6992\
        );

    \I__1246\ : Span12Mux_h
    port map (
            O => \N__6995\,
            I => \N__6989\
        );

    \I__1245\ : Span12Mux_v
    port map (
            O => \N__6992\,
            I => \N__6986\
        );

    \I__1244\ : Odrv12
    port map (
            O => \N__6989\,
            I => \TSn_c\
        );

    \I__1243\ : Odrv12
    port map (
            O => \N__6986\,
            I => \TSn_c\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__6981\,
            I => \U712_CHIP_RAM.N_458_cascade_\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6978\,
            I => \N__6975\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__6975\,
            I => \N__6972\
        );

    \I__1239\ : Span4Mux_v
    port map (
            O => \N__6972\,
            I => \N__6969\
        );

    \I__1238\ : Sp12to4
    port map (
            O => \N__6969\,
            I => \N__6965\
        );

    \I__1237\ : IoInMux
    port map (
            O => \N__6968\,
            I => \N__6962\
        );

    \I__1236\ : Span12Mux_h
    port map (
            O => \N__6965\,
            I => \N__6959\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6962\,
            I => \N__6956\
        );

    \I__1234\ : Span12Mux_v
    port map (
            O => \N__6959\,
            I => \N__6953\
        );

    \I__1233\ : IoSpan4Mux
    port map (
            O => \N__6956\,
            I => \N__6950\
        );

    \I__1232\ : Odrv12
    port map (
            O => \N__6953\,
            I => \RAMENn_c\
        );

    \I__1231\ : Odrv4
    port map (
            O => \N__6950\,
            I => \RAMENn_c\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__6945\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_1_cascade_\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__6942\,
            I => \N__6936\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6933\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6926\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6939\,
            I => \N__6926\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6936\,
            I => \N__6926\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6933\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6926\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__6921\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_0_cascade_\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6918\,
            I => \N__6915\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6915\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0\
        );

    \I__1219\ : IoInMux
    port map (
            O => \N__6912\,
            I => \N__6909\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6909\,
            I => \N__6906\
        );

    \I__1217\ : Span4Mux_s1_h
    port map (
            O => \N__6906\,
            I => \N__6903\
        );

    \I__1216\ : Sp12to4
    port map (
            O => \N__6903\,
            I => \N__6900\
        );

    \I__1215\ : Span12Mux_s11_v
    port map (
            O => \N__6900\,
            I => \N__6897\
        );

    \I__1214\ : Odrv12
    port map (
            O => \N__6897\,
            I => \CLK_EN_c\
        );

    \I__1213\ : CEMux
    port map (
            O => \N__6894\,
            I => \N__6891\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__6891\,
            I => \N__6888\
        );

    \I__1211\ : Odrv12
    port map (
            O => \N__6888\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__6885\,
            I => \U712_CHIP_RAM.N_344_cascade_\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6882\,
            I => \N__6879\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6879\,
            I => \U712_CHIP_RAM.N_435\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6876\,
            I => \N__6870\
        );

    \I__1206\ : InMux
    port map (
            O => \N__6875\,
            I => \N__6870\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6870\,
            I => \N__6867\
        );

    \I__1204\ : Odrv4
    port map (
            O => \N__6867\,
            I => \U712_CHIP_RAM.N_430\
        );

    \I__1203\ : InMux
    port map (
            O => \N__6864\,
            I => \N__6861\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6861\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\
        );

    \I__1201\ : CascadeMux
    port map (
            O => \N__6858\,
            I => \N__6855\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6855\,
            I => \N__6840\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6854\,
            I => \N__6840\
        );

    \I__1198\ : InMux
    port map (
            O => \N__6853\,
            I => \N__6840\
        );

    \I__1197\ : InMux
    port map (
            O => \N__6852\,
            I => \N__6840\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6851\,
            I => \N__6836\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6850\,
            I => \N__6831\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6831\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6840\,
            I => \N__6828\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6839\,
            I => \N__6825\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N__6822\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__6831\,
            I => \N__6818\
        );

    \I__1189\ : Span4Mux_h
    port map (
            O => \N__6828\,
            I => \N__6813\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__6825\,
            I => \N__6813\
        );

    \I__1187\ : Span12Mux_h
    port map (
            O => \N__6822\,
            I => \N__6810\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6821\,
            I => \N__6807\
        );

    \I__1185\ : Span4Mux_h
    port map (
            O => \N__6818\,
            I => \N__6802\
        );

    \I__1184\ : Span4Mux_h
    port map (
            O => \N__6813\,
            I => \N__6802\
        );

    \I__1183\ : Odrv12
    port map (
            O => \N__6810\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6807\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__6802\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6795\,
            I => \N__6789\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6794\,
            I => \N__6789\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6789\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_1\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__6786\,
            I => \N__6783\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6783\,
            I => \N__6780\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6780\,
            I => \U712_CHIP_RAM.N_362\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__6777\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_165_i_i_0_cascade_\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6770\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6767\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6770\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6767\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6759\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6759\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_a2_1_0\
        );

    \I__1167\ : InMux
    port map (
            O => \N__6756\,
            I => \N__6753\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6753\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER19\
        );

    \I__1165\ : CascadeMux
    port map (
            O => \N__6750\,
            I => \N__6747\
        );

    \I__1164\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6743\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6746\,
            I => \N__6740\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6743\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__6740\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__6735\,
            I => \N__6731\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6734\,
            I => \N__6728\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6725\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6728\,
            I => \DBR_SYNC_i_1\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6725\,
            I => \DBR_SYNC_i_1\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__6720\,
            I => \N__6717\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6717\,
            I => \N__6714\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6714\,
            I => \N__6711\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__6711\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6708\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6705\,
            I => \N__6701\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6704\,
            I => \N__6698\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6701\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6698\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6693\,
            I => \N__6690\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__6690\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6687\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6684\,
            I => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__6681\,
            I => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3_cascade_\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6674\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6677\,
            I => \N__6671\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__6674\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6671\,
            I => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6666\,
            I => \N__6663\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6663\,
            I => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__6660\,
            I => \U712_CHIP_RAM.N_451_cascade_\
        );

    \I__1134\ : CEMux
    port map (
            O => \N__6657\,
            I => \N__6654\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6654\,
            I => \U712_CHIP_RAM.N_452_0\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6648\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6648\,
            I => \N__6644\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6647\,
            I => \N__6641\
        );

    \I__1129\ : Odrv4
    port map (
            O => \N__6644\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_2\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6641\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_2\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__6636\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_cascade_\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6633\,
            I => \N__6630\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6630\,
            I => \N__6626\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6623\
        );

    \I__1123\ : Span4Mux_h
    port map (
            O => \N__6626\,
            I => \N__6620\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6623\,
            I => \U712_REG_SM.N_406\
        );

    \I__1121\ : Odrv4
    port map (
            O => \N__6620\,
            I => \U712_REG_SM.N_406\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6612\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6612\,
            I => \N__6609\
        );

    \I__1118\ : Span4Mux_h
    port map (
            O => \N__6609\,
            I => \N__6602\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6608\,
            I => \N__6597\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6597\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6606\,
            I => \N__6592\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6605\,
            I => \N__6592\
        );

    \I__1113\ : Odrv4
    port map (
            O => \N__6602\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6597\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__6592\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_8\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6585\,
            I => \N__6578\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__6584\,
            I => \N__6574\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6571\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6568\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6565\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6578\,
            I => \N__6562\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6553\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6574\,
            I => \N__6553\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6571\,
            I => \N__6550\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__6568\,
            I => \N__6545\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6565\,
            I => \N__6545\
        );

    \I__1099\ : Span4Mux_h
    port map (
            O => \N__6562\,
            I => \N__6542\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6561\,
            I => \N__6535\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6560\,
            I => \N__6535\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6559\,
            I => \N__6535\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6558\,
            I => \N__6532\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6553\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1093\ : Odrv12
    port map (
            O => \N__6550\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__6545\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__6542\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__6535\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__6532\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__6519\,
            I => \U712_REG_SM.N_445_cascade_\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6516\,
            I => \N__6513\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6513\,
            I => \N__6510\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__6510\,
            I => \U712_REG_SM.REG_CYCLE_5_iv_0_0\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6507\,
            I => \N__6504\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__6504\,
            I => \U712_BYTE_ENABLE.LMBE_0_i_o3_0_oZ0Z2\
        );

    \I__1082\ : IoInMux
    port map (
            O => \N__6501\,
            I => \N__6498\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__6498\,
            I => \N__6495\
        );

    \I__1080\ : Span4Mux_s2_v
    port map (
            O => \N__6495\,
            I => \N__6492\
        );

    \I__1079\ : Span4Mux_h
    port map (
            O => \N__6492\,
            I => \N__6489\
        );

    \I__1078\ : Span4Mux_h
    port map (
            O => \N__6489\,
            I => \N__6486\
        );

    \I__1077\ : Span4Mux_v
    port map (
            O => \N__6486\,
            I => \N__6483\
        );

    \I__1076\ : Odrv4
    port map (
            O => \N__6483\,
            I => \N_282_i\
        );

    \I__1075\ : IoInMux
    port map (
            O => \N__6480\,
            I => \N__6477\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6477\,
            I => \N__6474\
        );

    \I__1073\ : Span4Mux_s2_v
    port map (
            O => \N__6474\,
            I => \N__6471\
        );

    \I__1072\ : Span4Mux_v
    port map (
            O => \N__6471\,
            I => \N__6468\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__6468\,
            I => \N_219\
        );

    \I__1070\ : IoInMux
    port map (
            O => \N__6465\,
            I => \N__6462\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6462\,
            I => \N__6459\
        );

    \I__1068\ : Span4Mux_s3_v
    port map (
            O => \N__6459\,
            I => \N__6456\
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__6456\,
            I => \N_60_i\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__6453\,
            I => \U712_CHIP_RAM.N_365_cascade_\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__6450\,
            I => \N__6446\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6449\,
            I => \N__6441\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6441\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__6441\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__6438\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6435\,
            I => \N__6432\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6432\,
            I => \N__6429\
        );

    \I__1058\ : Span12Mux_h
    port map (
            O => \N__6429\,
            I => \N__6426\
        );

    \I__1057\ : Span12Mux_v
    port map (
            O => \N__6426\,
            I => \N__6423\
        );

    \I__1056\ : Odrv12
    port map (
            O => \N__6423\,
            I => \A_c_2\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6420\,
            I => \N__6417\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__6417\,
            I => \N__6414\
        );

    \I__1053\ : Span12Mux_v
    port map (
            O => \N__6414\,
            I => \N__6411\
        );

    \I__1052\ : Span12Mux_h
    port map (
            O => \N__6411\,
            I => \N__6408\
        );

    \I__1051\ : Odrv12
    port map (
            O => \N__6408\,
            I => \A_c_3\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6405\,
            I => \N__6402\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6402\,
            I => \N__6399\
        );

    \I__1048\ : Odrv4
    port map (
            O => \N__6399\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6396\,
            I => \N__6393\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6393\,
            I => \N__6390\
        );

    \I__1045\ : Span12Mux_v
    port map (
            O => \N__6390\,
            I => \N__6387\
        );

    \I__1044\ : Span12Mux_h
    port map (
            O => \N__6387\,
            I => \N__6384\
        );

    \I__1043\ : Odrv12
    port map (
            O => \N__6384\,
            I => \A_c_4\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6381\,
            I => \N__6378\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__6378\,
            I => \N__6375\
        );

    \I__1040\ : Span4Mux_v
    port map (
            O => \N__6375\,
            I => \N__6372\
        );

    \I__1039\ : Sp12to4
    port map (
            O => \N__6372\,
            I => \N__6369\
        );

    \I__1038\ : Span12Mux_h
    port map (
            O => \N__6369\,
            I => \N__6366\
        );

    \I__1037\ : Odrv12
    port map (
            O => \N__6366\,
            I => \A_c_7\
        );

    \I__1036\ : IoInMux
    port map (
            O => \N__6363\,
            I => \N__6360\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6360\,
            I => \N__6357\
        );

    \I__1034\ : IoSpan4Mux
    port map (
            O => \N__6357\,
            I => \N__6354\
        );

    \I__1033\ : Span4Mux_s0_v
    port map (
            O => \N__6354\,
            I => \N__6350\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__6353\,
            I => \N__6345\
        );

    \I__1031\ : Sp12to4
    port map (
            O => \N__6350\,
            I => \N__6342\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6339\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6334\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6345\,
            I => \N__6334\
        );

    \I__1027\ : Span12Mux_v
    port map (
            O => \N__6342\,
            I => \N__6330\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__6339\,
            I => \N__6327\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6334\,
            I => \N__6324\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6333\,
            I => \N__6321\
        );

    \I__1023\ : Odrv12
    port map (
            O => \N__6330\,
            I => \DBENn_c\
        );

    \I__1022\ : Odrv4
    port map (
            O => \N__6327\,
            I => \DBENn_c\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__6324\,
            I => \DBENn_c\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6321\,
            I => \DBENn_c\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6309\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__6309\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1Z0Z_0\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__6306\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1Z0Z_0_cascade_\
        );

    \I__1016\ : IoInMux
    port map (
            O => \N__6303\,
            I => \N__6300\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6300\,
            I => \N__6297\
        );

    \I__1014\ : Span4Mux_s2_h
    port map (
            O => \N__6297\,
            I => \N__6294\
        );

    \I__1013\ : Sp12to4
    port map (
            O => \N__6294\,
            I => \N__6291\
        );

    \I__1012\ : Span12Mux_v
    port map (
            O => \N__6291\,
            I => \N__6288\
        );

    \I__1011\ : Span12Mux_h
    port map (
            O => \N__6288\,
            I => \N__6285\
        );

    \I__1010\ : Odrv12
    port map (
            O => \N__6285\,
            I => \N_62_i\
        );

    \I__1009\ : CascadeMux
    port map (
            O => \N__6282\,
            I => \U712_CHIP_RAM.N_596_cascade_\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6279\,
            I => \N__6276\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6276\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__6273\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6266\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6263\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6266\,
            I => \U712_CHIP_RAM.N_596\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6263\,
            I => \U712_CHIP_RAM.N_596\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__6258\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_0_cascade_\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6255\,
            I => \N__6251\
        );

    \I__999\ : InMux
    port map (
            O => \N__6254\,
            I => \N__6248\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__6251\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__6248\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\
        );

    \I__996\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6240\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__6240\,
            I => \N__6236\
        );

    \I__994\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6233\
        );

    \I__993\ : Span4Mux_v
    port map (
            O => \N__6236\,
            I => \N__6229\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__6233\,
            I => \N__6226\
        );

    \I__991\ : InMux
    port map (
            O => \N__6232\,
            I => \N__6223\
        );

    \I__990\ : Sp12to4
    port map (
            O => \N__6229\,
            I => \N__6220\
        );

    \I__989\ : Sp12to4
    port map (
            O => \N__6226\,
            I => \N__6215\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__6223\,
            I => \N__6215\
        );

    \I__987\ : Span12Mux_h
    port map (
            O => \N__6220\,
            I => \N__6212\
        );

    \I__986\ : Span12Mux_h
    port map (
            O => \N__6215\,
            I => \N__6209\
        );

    \I__985\ : Span12Mux_v
    port map (
            O => \N__6212\,
            I => \N__6206\
        );

    \I__984\ : Span12Mux_v
    port map (
            O => \N__6209\,
            I => \N__6203\
        );

    \I__983\ : Odrv12
    port map (
            O => \N__6206\,
            I => \AWEn_c\
        );

    \I__982\ : Odrv12
    port map (
            O => \N__6203\,
            I => \AWEn_c\
        );

    \I__981\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6194\
        );

    \I__980\ : InMux
    port map (
            O => \N__6197\,
            I => \N__6191\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__6194\,
            I => \N__6188\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6191\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__977\ : Odrv4
    port map (
            O => \N__6188\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__6183\,
            I => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_i_i_a2_0_cascade_\
        );

    \I__975\ : InMux
    port map (
            O => \N__6180\,
            I => \N__6173\
        );

    \I__974\ : InMux
    port map (
            O => \N__6179\,
            I => \N__6173\
        );

    \I__973\ : InMux
    port map (
            O => \N__6178\,
            I => \N__6170\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__6173\,
            I => \N__6167\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__6170\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__970\ : Odrv4
    port map (
            O => \N__6167\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__969\ : InMux
    port map (
            O => \N__6162\,
            I => \N__6159\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__6159\,
            I => \U712_CHIP_RAM.N_365\
        );

    \I__967\ : SRMux
    port map (
            O => \N__6156\,
            I => \N__6153\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__6153\,
            I => \N__6150\
        );

    \I__965\ : Span4Mux_h
    port map (
            O => \N__6150\,
            I => \N__6146\
        );

    \I__964\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6143\
        );

    \I__963\ : Span4Mux_h
    port map (
            O => \N__6146\,
            I => \N__6140\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__6143\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__961\ : Odrv4
    port map (
            O => \N__6140\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__6135\,
            I => \U712_CHIP_RAM.N_362_cascade_\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__6132\,
            I => \U712_CHIP_RAM.N_493_cascade_\
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__6129\,
            I => \U712_CHIP_RAM.N_503_cascade_\
        );

    \I__957\ : InMux
    port map (
            O => \N__6126\,
            I => \N__6123\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__6123\,
            I => \N__6120\
        );

    \I__955\ : Odrv12
    port map (
            O => \N__6120\,
            I => \U712_REG_SM.N_482\
        );

    \I__954\ : InMux
    port map (
            O => \N__6117\,
            I => \N__6113\
        );

    \I__953\ : IoInMux
    port map (
            O => \N__6116\,
            I => \N__6110\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__6113\,
            I => \N__6107\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__6110\,
            I => \N__6104\
        );

    \I__950\ : Span12Mux_h
    port map (
            O => \N__6107\,
            I => \N__6101\
        );

    \I__949\ : IoSpan4Mux
    port map (
            O => \N__6104\,
            I => \N__6098\
        );

    \I__948\ : Span12Mux_h
    port map (
            O => \N__6101\,
            I => \N__6095\
        );

    \I__947\ : IoSpan4Mux
    port map (
            O => \N__6098\,
            I => \N__6092\
        );

    \I__946\ : Span12Mux_v
    port map (
            O => \N__6095\,
            I => \N__6089\
        );

    \I__945\ : IoSpan4Mux
    port map (
            O => \N__6092\,
            I => \N__6086\
        );

    \I__944\ : Odrv12
    port map (
            O => \N__6089\,
            I => \C1_c\
        );

    \I__943\ : Odrv4
    port map (
            O => \N__6086\,
            I => \C1_c\
        );

    \I__942\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6078\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__6078\,
            I => \N__6075\
        );

    \I__940\ : Odrv12
    port map (
            O => \N__6075\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__939\ : InMux
    port map (
            O => \N__6072\,
            I => \N__6069\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__6069\,
            I => \N__6066\
        );

    \I__937\ : Odrv4
    port map (
            O => \N__6066\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__936\ : IoInMux
    port map (
            O => \N__6063\,
            I => \N__6060\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__6060\,
            I => \N__6057\
        );

    \I__934\ : Span4Mux_s2_h
    port map (
            O => \N__6057\,
            I => \N__6054\
        );

    \I__933\ : Span4Mux_v
    port map (
            O => \N__6054\,
            I => \N__6051\
        );

    \I__932\ : Sp12to4
    port map (
            O => \N__6051\,
            I => \N__6048\
        );

    \I__931\ : Span12Mux_h
    port map (
            O => \N__6048\,
            I => \N__6045\
        );

    \I__930\ : Odrv12
    port map (
            O => \N__6045\,
            I => \CMA_c_6\
        );

    \I__929\ : InMux
    port map (
            O => \N__6042\,
            I => \N__6039\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__6039\,
            I => \N__6036\
        );

    \I__927\ : Odrv4
    port map (
            O => \N__6036\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__926\ : IoInMux
    port map (
            O => \N__6033\,
            I => \N__6030\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__6030\,
            I => \N__6027\
        );

    \I__924\ : Span4Mux_s3_h
    port map (
            O => \N__6027\,
            I => \N__6024\
        );

    \I__923\ : Span4Mux_v
    port map (
            O => \N__6024\,
            I => \N__6021\
        );

    \I__922\ : Sp12to4
    port map (
            O => \N__6021\,
            I => \N__6018\
        );

    \I__921\ : Span12Mux_h
    port map (
            O => \N__6018\,
            I => \N__6015\
        );

    \I__920\ : Odrv12
    port map (
            O => \N__6015\,
            I => \CMA_c_7\
        );

    \I__919\ : InMux
    port map (
            O => \N__6012\,
            I => \N__6009\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__6009\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\
        );

    \I__917\ : IoInMux
    port map (
            O => \N__6006\,
            I => \N__6003\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__6003\,
            I => \N__6000\
        );

    \I__915\ : Span4Mux_s2_h
    port map (
            O => \N__6000\,
            I => \N__5997\
        );

    \I__914\ : Sp12to4
    port map (
            O => \N__5997\,
            I => \N__5994\
        );

    \I__913\ : Span12Mux_s9_v
    port map (
            O => \N__5994\,
            I => \N__5991\
        );

    \I__912\ : Span12Mux_h
    port map (
            O => \N__5991\,
            I => \N__5988\
        );

    \I__911\ : Odrv12
    port map (
            O => \N__5988\,
            I => \CMA_c_8\
        );

    \I__910\ : InMux
    port map (
            O => \N__5985\,
            I => \N__5982\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5982\,
            I => \N__5979\
        );

    \I__908\ : Span4Mux_v
    port map (
            O => \N__5979\,
            I => \N__5976\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__5976\,
            I => \U712_REG_SM.N_481\
        );

    \I__906\ : IoInMux
    port map (
            O => \N__5973\,
            I => \N__5970\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5970\,
            I => \N__5967\
        );

    \I__904\ : Span4Mux_s2_v
    port map (
            O => \N__5967\,
            I => \N__5964\
        );

    \I__903\ : Sp12to4
    port map (
            O => \N__5964\,
            I => \N__5961\
        );

    \I__902\ : Span12Mux_h
    port map (
            O => \N__5961\,
            I => \N__5958\
        );

    \I__901\ : Span12Mux_v
    port map (
            O => \N__5958\,
            I => \N__5954\
        );

    \I__900\ : InMux
    port map (
            O => \N__5957\,
            I => \N__5951\
        );

    \I__899\ : Odrv12
    port map (
            O => \N__5954\,
            I => \LDSn_c\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__5951\,
            I => \LDSn_c\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__5946\,
            I => \N__5942\
        );

    \I__896\ : InMux
    port map (
            O => \N__5945\,
            I => \N__5937\
        );

    \I__895\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5937\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__5937\,
            I => \U712_REG_SM.N_185\
        );

    \I__893\ : IoInMux
    port map (
            O => \N__5934\,
            I => \N__5931\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5931\,
            I => \N__5928\
        );

    \I__891\ : IoSpan4Mux
    port map (
            O => \N__5928\,
            I => \N__5925\
        );

    \I__890\ : Sp12to4
    port map (
            O => \N__5925\,
            I => \N__5922\
        );

    \I__889\ : Span12Mux_s6_v
    port map (
            O => \N__5922\,
            I => \N__5919\
        );

    \I__888\ : Span12Mux_v
    port map (
            O => \N__5919\,
            I => \N__5915\
        );

    \I__887\ : InMux
    port map (
            O => \N__5918\,
            I => \N__5912\
        );

    \I__886\ : Odrv12
    port map (
            O => \N__5915\,
            I => \UDSn_c\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5912\,
            I => \UDSn_c\
        );

    \I__884\ : CascadeMux
    port map (
            O => \N__5907\,
            I => \N__5904\
        );

    \I__883\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5901\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5901\,
            I => \N__5898\
        );

    \I__881\ : Odrv12
    port map (
            O => \N__5898\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0Z0Z_0\
        );

    \I__880\ : InMux
    port map (
            O => \N__5895\,
            I => \N__5892\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5892\,
            I => \N__5889\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__5889\,
            I => \U712_BYTE_ENABLE.N_468\
        );

    \I__877\ : IoInMux
    port map (
            O => \N__5886\,
            I => \N__5883\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5883\,
            I => \N__5880\
        );

    \I__875\ : IoSpan4Mux
    port map (
            O => \N__5880\,
            I => \N__5877\
        );

    \I__874\ : Span4Mux_s1_h
    port map (
            O => \N__5877\,
            I => \N__5874\
        );

    \I__873\ : Sp12to4
    port map (
            O => \N__5874\,
            I => \N__5871\
        );

    \I__872\ : Span12Mux_h
    port map (
            O => \N__5871\,
            I => \N__5868\
        );

    \I__871\ : Span12Mux_v
    port map (
            O => \N__5868\,
            I => \N__5865\
        );

    \I__870\ : Odrv12
    port map (
            O => \N__5865\,
            I => \N_65_i\
        );

    \I__869\ : InMux
    port map (
            O => \N__5862\,
            I => \N__5855\
        );

    \I__868\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5855\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__5860\,
            I => \N__5852\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__5855\,
            I => \N__5849\
        );

    \I__865\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5846\
        );

    \I__864\ : Span4Mux_v
    port map (
            O => \N__5849\,
            I => \N__5843\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5846\,
            I => \N__5840\
        );

    \I__862\ : Odrv4
    port map (
            O => \N__5843\,
            I => \U712_BYTE_ENABLE.N_343_i\
        );

    \I__861\ : Odrv4
    port map (
            O => \N__5840\,
            I => \U712_BYTE_ENABLE.N_343_i\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__5835\,
            I => \U712_BYTE_ENABLE.N_466_cascade_\
        );

    \I__859\ : IoInMux
    port map (
            O => \N__5832\,
            I => \N__5829\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5829\,
            I => \N__5826\
        );

    \I__857\ : Span12Mux_s3_h
    port map (
            O => \N__5826\,
            I => \N__5823\
        );

    \I__856\ : Span12Mux_h
    port map (
            O => \N__5823\,
            I => \N__5820\
        );

    \I__855\ : Odrv12
    port map (
            O => \N__5820\,
            I => \N_67_i\
        );

    \I__854\ : IoInMux
    port map (
            O => \N__5817\,
            I => \N__5814\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5814\,
            I => \N__5811\
        );

    \I__852\ : Span12Mux_s4_v
    port map (
            O => \N__5811\,
            I => \N__5808\
        );

    \I__851\ : Span12Mux_h
    port map (
            O => \N__5808\,
            I => \N__5805\
        );

    \I__850\ : Odrv12
    port map (
            O => \N__5805\,
            I => \ASn_c\
        );

    \I__849\ : CEMux
    port map (
            O => \N__5802\,
            I => \N__5799\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5799\,
            I => \N__5796\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__5796\,
            I => \U712_REG_SM.N_185_0\
        );

    \I__846\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5787\
        );

    \I__845\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5787\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__5787\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\
        );

    \I__843\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5781\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5781\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\
        );

    \I__841\ : InMux
    port map (
            O => \N__5778\,
            I => \N__5775\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5775\,
            I => \N__5772\
        );

    \I__839\ : Sp12to4
    port map (
            O => \N__5772\,
            I => \N__5769\
        );

    \I__838\ : Span12Mux_v
    port map (
            O => \N__5769\,
            I => \N__5766\
        );

    \I__837\ : Span12Mux_h
    port map (
            O => \N__5766\,
            I => \N__5763\
        );

    \I__836\ : Odrv12
    port map (
            O => \N__5763\,
            I => \A_c_8\
        );

    \I__835\ : InMux
    port map (
            O => \N__5760\,
            I => \N__5757\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5757\,
            I => \N__5754\
        );

    \I__833\ : Odrv4
    port map (
            O => \N__5754\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\
        );

    \I__832\ : InMux
    port map (
            O => \N__5751\,
            I => \N__5748\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5748\,
            I => \N__5745\
        );

    \I__830\ : Sp12to4
    port map (
            O => \N__5745\,
            I => \N__5742\
        );

    \I__829\ : Span12Mux_v
    port map (
            O => \N__5742\,
            I => \N__5739\
        );

    \I__828\ : Span12Mux_h
    port map (
            O => \N__5739\,
            I => \N__5736\
        );

    \I__827\ : Odrv12
    port map (
            O => \N__5736\,
            I => \A_c_18\
        );

    \I__826\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5730\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5730\,
            I => \N__5727\
        );

    \I__824\ : Odrv4
    port map (
            O => \N__5727\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\
        );

    \I__823\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5721\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__5721\,
            I => \N__5718\
        );

    \I__821\ : Sp12to4
    port map (
            O => \N__5718\,
            I => \N__5715\
        );

    \I__820\ : Span12Mux_v
    port map (
            O => \N__5715\,
            I => \N__5712\
        );

    \I__819\ : Span12Mux_h
    port map (
            O => \N__5712\,
            I => \N__5709\
        );

    \I__818\ : Odrv12
    port map (
            O => \N__5709\,
            I => \A_c_20\
        );

    \I__817\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5702\
        );

    \I__816\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5699\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5702\,
            I => \N__5696\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__5699\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__813\ : Odrv4
    port map (
            O => \N__5696\,
            I => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\
        );

    \I__812\ : InMux
    port map (
            O => \N__5691\,
            I => \N__5688\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5688\,
            I => \N__5685\
        );

    \I__810\ : Span4Mux_v
    port map (
            O => \N__5685\,
            I => \N__5682\
        );

    \I__809\ : Span4Mux_v
    port map (
            O => \N__5682\,
            I => \N__5679\
        );

    \I__808\ : Sp12to4
    port map (
            O => \N__5679\,
            I => \N__5676\
        );

    \I__807\ : Span12Mux_h
    port map (
            O => \N__5676\,
            I => \N__5673\
        );

    \I__806\ : Odrv12
    port map (
            O => \N__5673\,
            I => \A_c_15\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__5670\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\
        );

    \I__804\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5664\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__5664\,
            I => \N__5659\
        );

    \I__802\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5656\
        );

    \I__801\ : InMux
    port map (
            O => \N__5662\,
            I => \N__5653\
        );

    \I__800\ : Span4Mux_h
    port map (
            O => \N__5659\,
            I => \N__5645\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5656\,
            I => \N__5640\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5653\,
            I => \N__5640\
        );

    \I__797\ : InMux
    port map (
            O => \N__5652\,
            I => \N__5635\
        );

    \I__796\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5635\
        );

    \I__795\ : InMux
    port map (
            O => \N__5650\,
            I => \N__5628\
        );

    \I__794\ : InMux
    port map (
            O => \N__5649\,
            I => \N__5628\
        );

    \I__793\ : InMux
    port map (
            O => \N__5648\,
            I => \N__5628\
        );

    \I__792\ : Odrv4
    port map (
            O => \N__5645\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__5640\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5635\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5628\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__788\ : InMux
    port map (
            O => \N__5619\,
            I => \N__5616\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__5616\,
            I => \U712_REG_SM.N_407\
        );

    \I__786\ : CascadeMux
    port map (
            O => \N__5613\,
            I => \U712_REG_SM.N_369_cascade_\
        );

    \I__785\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5606\
        );

    \I__784\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5603\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5606\,
            I => \N__5600\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5603\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__781\ : Odrv4
    port map (
            O => \N__5600\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__780\ : CEMux
    port map (
            O => \N__5595\,
            I => \N__5592\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5592\,
            I => \N__5589\
        );

    \I__778\ : Span4Mux_v
    port map (
            O => \N__5589\,
            I => \N__5586\
        );

    \I__777\ : Odrv4
    port map (
            O => \N__5586\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0\
        );

    \I__776\ : InMux
    port map (
            O => \N__5583\,
            I => \N__5580\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5580\,
            I => \N__5577\
        );

    \I__774\ : Span4Mux_v
    port map (
            O => \N__5577\,
            I => \N__5574\
        );

    \I__773\ : Span4Mux_v
    port map (
            O => \N__5574\,
            I => \N__5571\
        );

    \I__772\ : Sp12to4
    port map (
            O => \N__5571\,
            I => \N__5568\
        );

    \I__771\ : Span12Mux_h
    port map (
            O => \N__5568\,
            I => \N__5565\
        );

    \I__770\ : Odrv12
    port map (
            O => \N__5565\,
            I => \A_c_17\
        );

    \I__769\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5559\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5559\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__5556\,
            I => \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__5553\,
            I => \U712_REG_SM.N_366_cascade_\
        );

    \I__765\ : InMux
    port map (
            O => \N__5550\,
            I => \N__5544\
        );

    \I__764\ : InMux
    port map (
            O => \N__5549\,
            I => \N__5544\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5544\,
            I => \U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0\
        );

    \I__762\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5538\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__5538\,
            I => \N__5534\
        );

    \I__760\ : ClkMux
    port map (
            O => \N__5537\,
            I => \N__5531\
        );

    \I__759\ : Span4Mux_v
    port map (
            O => \N__5534\,
            I => \N__5527\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5531\,
            I => \N__5524\
        );

    \I__757\ : ClkMux
    port map (
            O => \N__5530\,
            I => \N__5521\
        );

    \I__756\ : Span4Mux_v
    port map (
            O => \N__5527\,
            I => \N__5514\
        );

    \I__755\ : Span4Mux_h
    port map (
            O => \N__5524\,
            I => \N__5514\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5521\,
            I => \N__5514\
        );

    \I__753\ : Span4Mux_v
    port map (
            O => \N__5514\,
            I => \N__5511\
        );

    \I__752\ : Span4Mux_v
    port map (
            O => \N__5511\,
            I => \N__5508\
        );

    \I__751\ : Odrv4
    port map (
            O => \N__5508\,
            I => \CLK40_PLL\
        );

    \I__750\ : IoInMux
    port map (
            O => \N__5505\,
            I => \N__5501\
        );

    \I__749\ : IoInMux
    port map (
            O => \N__5504\,
            I => \N__5498\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5501\,
            I => \N__5495\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__5498\,
            I => \N__5492\
        );

    \I__746\ : Span4Mux_s0_v
    port map (
            O => \N__5495\,
            I => \N__5489\
        );

    \I__745\ : Span4Mux_s3_v
    port map (
            O => \N__5492\,
            I => \N__5486\
        );

    \I__744\ : Span4Mux_v
    port map (
            O => \N__5489\,
            I => \N__5483\
        );

    \I__743\ : Span4Mux_h
    port map (
            O => \N__5486\,
            I => \N__5480\
        );

    \I__742\ : Sp12to4
    port map (
            O => \N__5483\,
            I => \N__5476\
        );

    \I__741\ : Span4Mux_h
    port map (
            O => \N__5480\,
            I => \N__5473\
        );

    \I__740\ : IoInMux
    port map (
            O => \N__5479\,
            I => \N__5470\
        );

    \I__739\ : Span12Mux_s11_h
    port map (
            O => \N__5476\,
            I => \N__5465\
        );

    \I__738\ : Sp12to4
    port map (
            O => \N__5473\,
            I => \N__5465\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__5470\,
            I => \N__5462\
        );

    \I__736\ : Span12Mux_v
    port map (
            O => \N__5465\,
            I => \N__5457\
        );

    \I__735\ : Span12Mux_s8_h
    port map (
            O => \N__5462\,
            I => \N__5457\
        );

    \I__734\ : Odrv12
    port map (
            O => \N__5457\,
            I => \CLK40_PLL_iso_i\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__5454\,
            I => \N__5449\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__5453\,
            I => \N__5446\
        );

    \I__731\ : CascadeMux
    port map (
            O => \N__5452\,
            I => \N__5443\
        );

    \I__730\ : InMux
    port map (
            O => \N__5449\,
            I => \N__5437\
        );

    \I__729\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5437\
        );

    \I__728\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5432\
        );

    \I__727\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5432\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5437\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5432\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__5427\,
            I => \N__5424\
        );

    \I__723\ : InMux
    port map (
            O => \N__5424\,
            I => \N__5421\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__5421\,
            I => \U712_REG_SM.N_375\
        );

    \I__721\ : InMux
    port map (
            O => \N__5418\,
            I => \N__5412\
        );

    \I__720\ : InMux
    port map (
            O => \N__5417\,
            I => \N__5409\
        );

    \I__719\ : InMux
    port map (
            O => \N__5416\,
            I => \N__5404\
        );

    \I__718\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5404\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5412\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5409\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5404\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__714\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5390\
        );

    \I__713\ : InMux
    port map (
            O => \N__5396\,
            I => \N__5390\
        );

    \I__712\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5387\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5390\,
            I => \N__5384\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5387\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__709\ : Odrv4
    port map (
            O => \N__5384\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__708\ : InMux
    port map (
            O => \N__5379\,
            I => \N__5373\
        );

    \I__707\ : InMux
    port map (
            O => \N__5378\,
            I => \N__5373\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5373\,
            I => \U712_REG_SM.N_483\
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__5370\,
            I => \U712_REG_SM.N_483_cascade_\
        );

    \I__704\ : InMux
    port map (
            O => \N__5367\,
            I => \N__5363\
        );

    \I__703\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5360\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5363\,
            I => \N__5356\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5360\,
            I => \N__5353\
        );

    \I__700\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5350\
        );

    \I__699\ : Odrv12
    port map (
            O => \N__5356\,
            I => \U712_REG_SM.N_367\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__5353\,
            I => \U712_REG_SM.N_367\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5350\,
            I => \U712_REG_SM.N_367\
        );

    \I__696\ : InMux
    port map (
            O => \N__5343\,
            I => \N__5337\
        );

    \I__695\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5333\
        );

    \I__694\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5328\
        );

    \I__693\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5328\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5337\,
            I => \N__5325\
        );

    \I__691\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5322\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5333\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5328\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__688\ : Odrv12
    port map (
            O => \N__5325\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__5322\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__686\ : InMux
    port map (
            O => \N__5313\,
            I => \N__5307\
        );

    \I__685\ : InMux
    port map (
            O => \N__5312\,
            I => \N__5304\
        );

    \I__684\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5299\
        );

    \I__683\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5299\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5307\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5304\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5299\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__679\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5285\
        );

    \I__678\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5280\
        );

    \I__677\ : InMux
    port map (
            O => \N__5290\,
            I => \N__5280\
        );

    \I__676\ : InMux
    port map (
            O => \N__5289\,
            I => \N__5275\
        );

    \I__675\ : InMux
    port map (
            O => \N__5288\,
            I => \N__5275\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__5285\,
            I => \U712_REG_SM.N_358\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__5280\,
            I => \U712_REG_SM.N_358\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__5275\,
            I => \U712_REG_SM.N_358\
        );

    \I__671\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5265\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__5265\,
            I => \U712_REG_SM.N_592\
        );

    \I__669\ : IoInMux
    port map (
            O => \N__5262\,
            I => \N__5258\
        );

    \I__668\ : IoInMux
    port map (
            O => \N__5261\,
            I => \N__5254\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__5258\,
            I => \N__5251\
        );

    \I__666\ : IoInMux
    port map (
            O => \N__5257\,
            I => \N__5248\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5254\,
            I => \N__5245\
        );

    \I__664\ : IoSpan4Mux
    port map (
            O => \N__5251\,
            I => \N__5242\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__5248\,
            I => \N__5239\
        );

    \I__662\ : Span4Mux_s2_h
    port map (
            O => \N__5245\,
            I => \N__5236\
        );

    \I__661\ : Span4Mux_s2_v
    port map (
            O => \N__5242\,
            I => \N__5233\
        );

    \I__660\ : Span4Mux_s2_v
    port map (
            O => \N__5239\,
            I => \N__5230\
        );

    \I__659\ : Sp12to4
    port map (
            O => \N__5236\,
            I => \N__5226\
        );

    \I__658\ : Span4Mux_v
    port map (
            O => \N__5233\,
            I => \N__5223\
        );

    \I__657\ : Span4Mux_v
    port map (
            O => \N__5230\,
            I => \N__5220\
        );

    \I__656\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5216\
        );

    \I__655\ : Span12Mux_v
    port map (
            O => \N__5226\,
            I => \N__5213\
        );

    \I__654\ : Sp12to4
    port map (
            O => \N__5223\,
            I => \N__5210\
        );

    \I__653\ : Sp12to4
    port map (
            O => \N__5220\,
            I => \N__5207\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__5219\,
            I => \N__5204\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__5216\,
            I => \N__5201\
        );

    \I__650\ : Span12Mux_h
    port map (
            O => \N__5213\,
            I => \N__5194\
        );

    \I__649\ : Span12Mux_h
    port map (
            O => \N__5210\,
            I => \N__5194\
        );

    \I__648\ : Span12Mux_h
    port map (
            O => \N__5207\,
            I => \N__5194\
        );

    \I__647\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5191\
        );

    \I__646\ : Span4Mux_v
    port map (
            O => \N__5201\,
            I => \N__5188\
        );

    \I__645\ : Odrv12
    port map (
            O => \N__5194\,
            I => \TACK_EN\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__5191\,
            I => \TACK_EN\
        );

    \I__643\ : Odrv4
    port map (
            O => \N__5188\,
            I => \TACK_EN\
        );

    \I__642\ : SRMux
    port map (
            O => \N__5181\,
            I => \N__5178\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__5178\,
            I => \N__5175\
        );

    \I__640\ : Span4Mux_h
    port map (
            O => \N__5175\,
            I => \N__5172\
        );

    \I__639\ : Span4Mux_h
    port map (
            O => \N__5172\,
            I => \N__5169\
        );

    \I__638\ : Odrv4
    port map (
            O => \N__5169\,
            I => \U712_CYCLE_TERM.TACK_RST_0_i\
        );

    \I__637\ : IoInMux
    port map (
            O => \N__5166\,
            I => \N__5163\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__5163\,
            I => \N__5160\
        );

    \I__635\ : Span12Mux_s5_v
    port map (
            O => \N__5160\,
            I => \N__5157\
        );

    \I__634\ : Odrv12
    port map (
            O => \N__5157\,
            I => \RESETn_c_i\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__5154\,
            I => \U712_REG_SM.N_185_cascade_\
        );

    \I__632\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5148\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__5148\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_7\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__5145\,
            I => \U712_REG_SM.N_368_cascade_\
        );

    \I__629\ : InMux
    port map (
            O => \N__5142\,
            I => \N__5139\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__5139\,
            I => \N__5136\
        );

    \I__627\ : Odrv4
    port map (
            O => \N__5136\,
            I => \U712_CHIP_RAM.N_378\
        );

    \I__626\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5128\
        );

    \I__625\ : InMux
    port map (
            O => \N__5132\,
            I => \N__5125\
        );

    \I__624\ : InMux
    port map (
            O => \N__5131\,
            I => \N__5122\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__5128\,
            I => \U712_REG_SM.N_441\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__5125\,
            I => \U712_REG_SM.N_441\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__5122\,
            I => \U712_REG_SM.N_441\
        );

    \I__620\ : CascadeMux
    port map (
            O => \N__5115\,
            I => \U712_REG_SM.N_358_cascade_\
        );

    \I__619\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5109\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__5109\,
            I => \U712_REG_SM.N_368\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__5106\,
            I => \N__5103\
        );

    \I__616\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5100\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__5100\,
            I => \U712_REG_SM.N_366\
        );

    \I__614\ : IoInMux
    port map (
            O => \N__5097\,
            I => \N__5094\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__5094\,
            I => \N__5091\
        );

    \I__612\ : Span12Mux_s7_v
    port map (
            O => \N__5091\,
            I => \N__5088\
        );

    \I__611\ : Odrv12
    port map (
            O => \N__5088\,
            I => \CMA_c_1\
        );

    \I__610\ : InMux
    port map (
            O => \N__5085\,
            I => \N__5081\
        );

    \I__609\ : InMux
    port map (
            O => \N__5084\,
            I => \N__5078\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__5081\,
            I => \N__5075\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__5078\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__606\ : Odrv4
    port map (
            O => \N__5075\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__605\ : InMux
    port map (
            O => \N__5070\,
            I => \N__5067\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__5067\,
            I => \N__5064\
        );

    \I__603\ : Span4Mux_v
    port map (
            O => \N__5064\,
            I => \N__5061\
        );

    \I__602\ : Sp12to4
    port map (
            O => \N__5061\,
            I => \N__5058\
        );

    \I__601\ : Span12Mux_h
    port map (
            O => \N__5058\,
            I => \N__5055\
        );

    \I__600\ : Odrv12
    port map (
            O => \N__5055\,
            I => \REGSPACEn_c\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__5052\,
            I => \U712_REG_SM.N_455_cascade_\
        );

    \I__598\ : IoInMux
    port map (
            O => \N__5049\,
            I => \N__5046\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__5046\,
            I => \N__5043\
        );

    \I__596\ : Span4Mux_s0_v
    port map (
            O => \N__5043\,
            I => \N__5040\
        );

    \I__595\ : Span4Mux_v
    port map (
            O => \N__5040\,
            I => \N__5036\
        );

    \I__594\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5033\
        );

    \I__593\ : Span4Mux_v
    port map (
            O => \N__5036\,
            I => \N__5030\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__5033\,
            I => \N__5027\
        );

    \I__591\ : Sp12to4
    port map (
            O => \N__5030\,
            I => \N__5024\
        );

    \I__590\ : Span4Mux_v
    port map (
            O => \N__5027\,
            I => \N__5021\
        );

    \I__589\ : Span12Mux_h
    port map (
            O => \N__5024\,
            I => \N__5018\
        );

    \I__588\ : Sp12to4
    port map (
            O => \N__5021\,
            I => \N__5015\
        );

    \I__587\ : Span12Mux_v
    port map (
            O => \N__5018\,
            I => \N__5010\
        );

    \I__586\ : Span12Mux_h
    port map (
            O => \N__5015\,
            I => \N__5010\
        );

    \I__585\ : Odrv12
    port map (
            O => \N__5010\,
            I => \A_c_10\
        );

    \I__584\ : InMux
    port map (
            O => \N__5007\,
            I => \N__5004\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__5004\,
            I => \U712_CHIP_RAM.N_387\
        );

    \I__582\ : InMux
    port map (
            O => \N__5001\,
            I => \N__4997\
        );

    \I__581\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4994\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4997\,
            I => \REG_TACK\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__4994\,
            I => \REG_TACK\
        );

    \I__578\ : IoInMux
    port map (
            O => \N__4989\,
            I => \N__4986\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__4986\,
            I => \N__4983\
        );

    \I__576\ : Span4Mux_s2_v
    port map (
            O => \N__4983\,
            I => \N__4980\
        );

    \I__575\ : Span4Mux_v
    port map (
            O => \N__4980\,
            I => \N__4977\
        );

    \I__574\ : Span4Mux_h
    port map (
            O => \N__4977\,
            I => \N__4974\
        );

    \I__573\ : Odrv4
    port map (
            O => \N__4974\,
            I => \VBENn_c\
        );

    \I__572\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4966\
        );

    \I__571\ : InMux
    port map (
            O => \N__4970\,
            I => \N__4961\
        );

    \I__570\ : InMux
    port map (
            O => \N__4969\,
            I => \N__4961\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__4966\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4961\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__4956\,
            I => \N__4952\
        );

    \I__566\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4948\
        );

    \I__565\ : InMux
    port map (
            O => \N__4952\,
            I => \N__4943\
        );

    \I__564\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4943\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4948\,
            I => \N__4937\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4943\,
            I => \N__4937\
        );

    \I__561\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4934\
        );

    \I__560\ : Span4Mux_v
    port map (
            O => \N__4937\,
            I => \N__4931\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4934\,
            I => \U712_CYCLE_TERM.TACK_STARTZ0\
        );

    \I__558\ : Odrv4
    port map (
            O => \N__4931\,
            I => \U712_CYCLE_TERM.TACK_STARTZ0\
        );

    \I__557\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4919\
        );

    \I__556\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4910\
        );

    \I__555\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4910\
        );

    \I__554\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4910\
        );

    \I__553\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4910\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__4919\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4910\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__4905\,
            I => \U712_CYCLE_TERM.N_36_0_cascade_\
        );

    \I__549\ : IoInMux
    port map (
            O => \N__4902\,
            I => \N__4898\
        );

    \I__548\ : IoInMux
    port map (
            O => \N__4901\,
            I => \N__4895\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4898\,
            I => \N__4891\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__4895\,
            I => \N__4888\
        );

    \I__545\ : IoInMux
    port map (
            O => \N__4894\,
            I => \N__4885\
        );

    \I__544\ : Span4Mux_s3_h
    port map (
            O => \N__4891\,
            I => \N__4882\
        );

    \I__543\ : IoSpan4Mux
    port map (
            O => \N__4888\,
            I => \N__4879\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4885\,
            I => \N__4876\
        );

    \I__541\ : Sp12to4
    port map (
            O => \N__4882\,
            I => \N__4873\
        );

    \I__540\ : Span4Mux_s3_v
    port map (
            O => \N__4879\,
            I => \N__4870\
        );

    \I__539\ : Span4Mux_s3_v
    port map (
            O => \N__4876\,
            I => \N__4867\
        );

    \I__538\ : Span12Mux_v
    port map (
            O => \N__4873\,
            I => \N__4864\
        );

    \I__537\ : Sp12to4
    port map (
            O => \N__4870\,
            I => \N__4861\
        );

    \I__536\ : Sp12to4
    port map (
            O => \N__4867\,
            I => \N__4858\
        );

    \I__535\ : Span12Mux_h
    port map (
            O => \N__4864\,
            I => \N__4850\
        );

    \I__534\ : Span12Mux_h
    port map (
            O => \N__4861\,
            I => \N__4850\
        );

    \I__533\ : Span12Mux_h
    port map (
            O => \N__4858\,
            I => \N__4850\
        );

    \I__532\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4847\
        );

    \I__531\ : Odrv12
    port map (
            O => \N__4850\,
            I => \TACK_OUT\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4847\,
            I => \TACK_OUT\
        );

    \I__529\ : InMux
    port map (
            O => \N__4842\,
            I => \N__4839\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__4839\,
            I => \N__4836\
        );

    \I__527\ : Span4Mux_h
    port map (
            O => \N__4836\,
            I => \N__4833\
        );

    \I__526\ : Sp12to4
    port map (
            O => \N__4833\,
            I => \N__4830\
        );

    \I__525\ : Span12Mux_v
    port map (
            O => \N__4830\,
            I => \N__4827\
        );

    \I__524\ : Span12Mux_h
    port map (
            O => \N__4827\,
            I => \N__4824\
        );

    \I__523\ : Odrv12
    port map (
            O => \N__4824\,
            I => \A_c_16\
        );

    \I__522\ : CascadeMux
    port map (
            O => \N__4821\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\
        );

    \I__521\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4815\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__4815\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_4\
        );

    \I__519\ : InMux
    port map (
            O => \N__4812\,
            I => \N__4806\
        );

    \I__518\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4806\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4806\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_5\
        );

    \I__516\ : InMux
    port map (
            O => \N__4803\,
            I => \N__4800\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4800\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_6\
        );

    \I__514\ : IoInMux
    port map (
            O => \N__4797\,
            I => \N__4794\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4794\,
            I => \N__4791\
        );

    \I__512\ : IoSpan4Mux
    port map (
            O => \N__4791\,
            I => \N__4788\
        );

    \I__511\ : Span4Mux_s2_v
    port map (
            O => \N__4788\,
            I => \N__4785\
        );

    \I__510\ : Span4Mux_v
    port map (
            O => \N__4785\,
            I => \N__4782\
        );

    \I__509\ : Sp12to4
    port map (
            O => \N__4782\,
            I => \N__4779\
        );

    \I__508\ : Span12Mux_v
    port map (
            O => \N__4779\,
            I => \N__4775\
        );

    \I__507\ : InMux
    port map (
            O => \N__4778\,
            I => \N__4772\
        );

    \I__506\ : Odrv12
    port map (
            O => \N__4775\,
            I => \PRnW_c\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4772\,
            I => \PRnW_c\
        );

    \I__504\ : InMux
    port map (
            O => \N__4767\,
            I => \N__4764\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__4764\,
            I => \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\
        );

    \I__502\ : IoInMux
    port map (
            O => \N__4761\,
            I => \N__4757\
        );

    \I__501\ : IoInMux
    port map (
            O => \N__4760\,
            I => \N__4754\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4757\,
            I => \N__4751\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4754\,
            I => \N__4748\
        );

    \I__498\ : IoSpan4Mux
    port map (
            O => \N__4751\,
            I => \N__4745\
        );

    \I__497\ : Span12Mux_s4_v
    port map (
            O => \N__4748\,
            I => \N__4742\
        );

    \I__496\ : Span4Mux_s3_v
    port map (
            O => \N__4745\,
            I => \N__4739\
        );

    \I__495\ : Span12Mux_h
    port map (
            O => \N__4742\,
            I => \N__4736\
        );

    \I__494\ : Sp12to4
    port map (
            O => \N__4739\,
            I => \N__4733\
        );

    \I__493\ : Span12Mux_v
    port map (
            O => \N__4736\,
            I => \N__4727\
        );

    \I__492\ : Span12Mux_v
    port map (
            O => \N__4733\,
            I => \N__4727\
        );

    \I__491\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4724\
        );

    \I__490\ : Odrv12
    port map (
            O => \N__4727\,
            I => \BLSn_c\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4724\,
            I => \BLSn_c\
        );

    \I__488\ : IoInMux
    port map (
            O => \N__4719\,
            I => \N__4716\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4716\,
            I => \N__4713\
        );

    \I__486\ : IoSpan4Mux
    port map (
            O => \N__4713\,
            I => \N__4710\
        );

    \I__485\ : Span4Mux_s3_v
    port map (
            O => \N__4710\,
            I => \N__4707\
        );

    \I__484\ : Sp12to4
    port map (
            O => \N__4707\,
            I => \N__4704\
        );

    \I__483\ : Span12Mux_v
    port map (
            O => \N__4704\,
            I => \N__4701\
        );

    \I__482\ : Odrv12
    port map (
            O => \N__4701\,
            I => \N_58_i\
        );

    \I__481\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4692\
        );

    \I__480\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4692\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4692\,
            I => \U712_BYTE_ENABLE.N_352\
        );

    \I__478\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4685\
        );

    \I__477\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4682\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4685\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__4682\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__474\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4673\
        );

    \I__473\ : InMux
    port map (
            O => \N__4676\,
            I => \N__4670\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4673\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__4670\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__470\ : CascadeMux
    port map (
            O => \N__4665\,
            I => \N__4661\
        );

    \I__469\ : InMux
    port map (
            O => \N__4664\,
            I => \N__4658\
        );

    \I__468\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4655\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4658\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4655\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__465\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4646\
        );

    \I__464\ : InMux
    port map (
            O => \N__4649\,
            I => \N__4643\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4646\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4643\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__461\ : IoInMux
    port map (
            O => \N__4638\,
            I => \N__4635\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4635\,
            I => \N__4632\
        );

    \I__459\ : Span12Mux_s0_v
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__458\ : Span12Mux_v
    port map (
            O => \N__4629\,
            I => \N__4625\
        );

    \I__457\ : InMux
    port map (
            O => \N__4628\,
            I => \N__4622\
        );

    \I__456\ : Odrv12
    port map (
            O => \N__4625\,
            I => \DBDIR_c\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4622\,
            I => \DBDIR_c\
        );

    \I__454\ : InMux
    port map (
            O => \N__4617\,
            I => \N__4614\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4614\,
            I => \N__4611\
        );

    \I__452\ : Odrv4
    port map (
            O => \N__4611\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__451\ : InMux
    port map (
            O => \N__4608\,
            I => \N__4605\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4605\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__449\ : InMux
    port map (
            O => \N__4602\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__448\ : InMux
    port map (
            O => \N__4599\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__447\ : InMux
    port map (
            O => \N__4596\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__446\ : InMux
    port map (
            O => \N__4593\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__445\ : InMux
    port map (
            O => \N__4590\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__444\ : InMux
    port map (
            O => \N__4587\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__443\ : ClkMux
    port map (
            O => \N__4584\,
            I => \N__4563\
        );

    \I__442\ : ClkMux
    port map (
            O => \N__4583\,
            I => \N__4563\
        );

    \I__441\ : ClkMux
    port map (
            O => \N__4582\,
            I => \N__4563\
        );

    \I__440\ : ClkMux
    port map (
            O => \N__4581\,
            I => \N__4563\
        );

    \I__439\ : ClkMux
    port map (
            O => \N__4580\,
            I => \N__4563\
        );

    \I__438\ : ClkMux
    port map (
            O => \N__4579\,
            I => \N__4563\
        );

    \I__437\ : ClkMux
    port map (
            O => \N__4578\,
            I => \N__4563\
        );

    \I__436\ : GlobalMux
    port map (
            O => \N__4563\,
            I => \N__4560\
        );

    \I__435\ : gio2CtrlBuf
    port map (
            O => \N__4560\,
            I => \C1_c_g\
        );

    \I__434\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4553\
        );

    \I__433\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4550\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4553\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__4550\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__430\ : InMux
    port map (
            O => \N__4545\,
            I => \N__4541\
        );

    \I__429\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4538\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__4541\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__4538\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__426\ : IoInMux
    port map (
            O => \N__4533\,
            I => \N__4530\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__4530\,
            I => \N__4527\
        );

    \I__424\ : IoSpan4Mux
    port map (
            O => \N__4527\,
            I => \N__4524\
        );

    \I__423\ : Span4Mux_s3_h
    port map (
            O => \N__4524\,
            I => \N__4521\
        );

    \I__422\ : Span4Mux_h
    port map (
            O => \N__4521\,
            I => \N__4517\
        );

    \I__421\ : InMux
    port map (
            O => \N__4520\,
            I => \N__4514\
        );

    \I__420\ : Span4Mux_h
    port map (
            O => \N__4517\,
            I => \N__4511\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__4514\,
            I => \N__4508\
        );

    \I__418\ : Span4Mux_h
    port map (
            O => \N__4511\,
            I => \N__4505\
        );

    \I__417\ : Span4Mux_v
    port map (
            O => \N__4508\,
            I => \N__4502\
        );

    \I__416\ : Sp12to4
    port map (
            O => \N__4505\,
            I => \N__4497\
        );

    \I__415\ : Sp12to4
    port map (
            O => \N__4502\,
            I => \N__4497\
        );

    \I__414\ : Span12Mux_h
    port map (
            O => \N__4497\,
            I => \N__4494\
        );

    \I__413\ : Span12Mux_v
    port map (
            O => \N__4494\,
            I => \N__4491\
        );

    \I__412\ : Odrv12
    port map (
            O => \N__4491\,
            I => \C3_c\
        );

    \I__411\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4485\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__4485\,
            I => \N__4481\
        );

    \I__409\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4478\
        );

    \I__408\ : Span4Mux_v
    port map (
            O => \N__4481\,
            I => \N__4475\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__4478\,
            I => \N__4472\
        );

    \I__406\ : Sp12to4
    port map (
            O => \N__4475\,
            I => \N__4469\
        );

    \I__405\ : Span12Mux_h
    port map (
            O => \N__4472\,
            I => \N__4466\
        );

    \I__404\ : Span12Mux_h
    port map (
            O => \N__4469\,
            I => \N__4463\
        );

    \I__403\ : Span12Mux_v
    port map (
            O => \N__4466\,
            I => \N__4460\
        );

    \I__402\ : Span12Mux_v
    port map (
            O => \N__4463\,
            I => \N__4457\
        );

    \I__401\ : Odrv12
    port map (
            O => \N__4460\,
            I => \DBRn_c\
        );

    \I__400\ : Odrv12
    port map (
            O => \N__4457\,
            I => \DBRn_c\
        );

    \I__399\ : IoInMux
    port map (
            O => \N__4452\,
            I => \N__4449\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__4449\,
            I => \N__4446\
        );

    \I__397\ : Span12Mux_s6_v
    port map (
            O => \N__4446\,
            I => \N__4443\
        );

    \I__396\ : Odrv12
    port map (
            O => \N__4443\,
            I => \CLK80_PLL_i_i\
        );

    \I__395\ : CascadeMux
    port map (
            O => \N__4440\,
            I => \DBRn_c_i_cascade_\
        );

    \I__394\ : IoInMux
    port map (
            O => \N__4437\,
            I => \N__4434\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__4434\,
            I => \N__4431\
        );

    \I__392\ : Span12Mux_s3_h
    port map (
            O => \N__4431\,
            I => \N__4428\
        );

    \I__391\ : Odrv12
    port map (
            O => \N__4428\,
            I => \DBRn_c_i_0\
        );

    \I__390\ : InMux
    port map (
            O => \N__4425\,
            I => \N__4422\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__4422\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__388\ : InMux
    port map (
            O => \N__4419\,
            I => \bfn_10_6_0_\
        );

    \I__387\ : InMux
    port map (
            O => \N__4416\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__386\ : IoInMux
    port map (
            O => \N__4413\,
            I => \N__4410\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__4410\,
            I => \N__4407\
        );

    \I__384\ : IoSpan4Mux
    port map (
            O => \N__4407\,
            I => \N__4404\
        );

    \I__383\ : Span4Mux_s2_v
    port map (
            O => \N__4404\,
            I => \N__4401\
        );

    \I__382\ : Sp12to4
    port map (
            O => \N__4401\,
            I => \N__4398\
        );

    \I__381\ : Span12Mux_v
    port map (
            O => \N__4398\,
            I => \N__4395\
        );

    \I__380\ : Odrv12
    port map (
            O => \N__4395\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            I => \N__4584\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__4582\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__4580\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__4581\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__4579\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            I => \N__4578\
        );

    \INVU712_CYCLE_TERM.TACK_STATE_0C\ : INV
    port map (
            O => \INVU712_CYCLE_TERM.TACK_STATE_0C_net\,
            I => \N__5530\
        );

    \INVU712_CYCLE_TERM.TACK_ENC\ : INV
    port map (
            O => \INVU712_CYCLE_TERM.TACK_ENC_net\,
            I => \N__5537\
        );

    \IN_MUX_bfv_10_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_6_0_\
        );

    \IN_MUX_bfv_16_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_6_0_\
        );

    \IN_MUX_bfv_15_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_4_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6116\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5166\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4437\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4533\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11742\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4488\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DBRn_c_i\,
            ltout => \DBRn_c_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11141\,
            in1 => \_gnd_net_\,
            in2 => \N__4440\,
            in3 => \_gnd_net_\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4425\,
            in2 => \_gnd_net_\,
            in3 => \N__4419\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_10_6_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__4583\,
            ce => 'H',
            sr => \N__6156\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4677\,
            in2 => \_gnd_net_\,
            in3 => \N__4416\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__4583\,
            ce => 'H',
            sr => \N__6156\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4650\,
            in2 => \_gnd_net_\,
            in3 => \N__4602\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__4583\,
            ce => 'H',
            sr => \N__6156\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4689\,
            in2 => \_gnd_net_\,
            in3 => \N__4599\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__4583\,
            ce => 'H',
            sr => \N__6156\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4664\,
            in2 => \_gnd_net_\,
            in3 => \N__4596\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__4583\,
            ce => 'H',
            sr => \N__6156\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4545\,
            in2 => \_gnd_net_\,
            in3 => \N__4593\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__4583\,
            ce => 'H',
            sr => \N__6156\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4557\,
            in2 => \_gnd_net_\,
            in3 => \N__4590\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__4583\,
            ce => 'H',
            sr => \N__6156\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9149\,
            in2 => \_gnd_net_\,
            in3 => \N__4587\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4583\,
            ce => 'H',
            sr => \N__6156\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4556\,
            in2 => \_gnd_net_\,
            in3 => \N__4544\,
            lcout => \U712_CHIP_RAM.REFRESH5lto7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4520\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11713\,
            ce => 'H',
            sr => \N__11081\
        );

    \DBR_SYNC_0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4484\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11720\,
            ce => 'H',
            sr => \N__11074\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000000"
        )
    port map (
            in0 => \N__7825\,
            in1 => \N__4698\,
            in2 => \N__5860\,
            in3 => \N__10516\,
            lcout => \U712_BYTE_ENABLE.N_468\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_58_i_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__7824\,
            in1 => \N__4697\,
            in2 => \N__5907\,
            in3 => \N__10515\,
            lcout => \N_58_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_o2_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7730\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7561\,
            lcout => \U712_BYTE_ENABLE.N_352\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_x2_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__7543\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7615\,
            lcout => \U712_BYTE_ENABLE.N_343_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100110000"
        )
    port map (
            in0 => \N__4926\,
            in1 => \N__4971\,
            in2 => \N__5219\,
            in3 => \N__4955\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_ENC_net\,
            ce => 'H',
            sr => \N__11096\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__4688\,
            in1 => \N__4676\,
            in2 => \N__4665\,
            in3 => \N__4649\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__6232\,
            in1 => \N__4628\,
            in2 => \_gnd_net_\,
            in3 => \N__6198\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11701\,
            ce => 'H',
            sr => \N__11082\
        );

    \DBR_SYNC_1_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4617\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11701\,
            ce => 'H',
            sr => \N__11082\
        );

    \U712_REG_SM.C3_SYNC_1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4608\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11707\,
            ce => 'H',
            sr => \N__11075\
        );

    \U712_REG_SM.STATE_COUNT_7_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12005\,
            in2 => \_gnd_net_\,
            in3 => \N__4803\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12003\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4818\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__12002\,
            in1 => \N__5312\,
            in2 => \_gnd_net_\,
            in3 => \N__5292\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_2_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4811\,
            in1 => \N__5417\,
            in2 => \_gnd_net_\,
            in3 => \N__5132\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12004\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4812\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.PRnW_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111101000101"
        )
    port map (
            in0 => \N__5550\,
            in1 => \N__5663\,
            in2 => \N__5453\,
            in3 => \N__4778\,
            lcout => \PRnW_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11721\,
            ce => 'H',
            sr => \N__11067\
        );

    \U712_REG_SM.WRITE_CYCLE_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__10955\,
            in1 => \_gnd_net_\,
            in2 => \N__5454\,
            in3 => \N__5379\,
            lcout => \U712_REG_SM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11721\,
            ce => 'H',
            sr => \N__11067\
        );

    \U712_REG_SM.REG_TACK_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__5001\,
            in1 => \N__4767\,
            in2 => \N__5427\,
            in3 => \N__5268\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11721\,
            ce => 'H',
            sr => \N__11067\
        );

    \U712_REG_SM.START_RST_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__5084\,
            in1 => \N__5342\,
            in2 => \_gnd_net_\,
            in3 => \N__5378\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11721\,
            ce => 'H',
            sr => \N__11067\
        );

    \U712_REG_SM.REGENn_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__5291\,
            in1 => \N__4732\,
            in2 => \_gnd_net_\,
            in3 => \N__5549\,
            lcout => \BLSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11721\,
            ce => 'H',
            sr => \N__11067\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110001111"
        )
    port map (
            in0 => \N__5418\,
            in1 => \N__5290\,
            in2 => \N__5106\,
            in3 => \N__5133\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11721\,
            ce => 'H',
            sr => \N__11067\
        );

    \U712_CYCLE_TERM.TACK_START_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5000\,
            in1 => \N__7194\,
            in2 => \_gnd_net_\,
            in3 => \N__4942\,
            lcout => \U712_CYCLE_TERM.TACK_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11726\,
            ce => 'H',
            sr => \N__5181\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__10499\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9381\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4924\,
            in1 => \N__11925\,
            in2 => \N__4956\,
            in3 => \N__4970\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11926\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4923\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUT_RNO_0_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__4969\,
            in1 => \N__4922\,
            in2 => \_gnd_net_\,
            in3 => \N__4951\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_36_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUT_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110110011"
        )
    port map (
            in0 => \N__4925\,
            in1 => \N__11924\,
            in2 => \N__4905\,
            in3 => \N__4857\,
            lcout => \TACK_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CYCLE_TERM.TACK_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5733\,
            in1 => \N__4842\,
            in2 => \_gnd_net_\,
            in3 => \N__9835\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9836\,
            in1 => \N__10498\,
            in2 => \N__4821\,
            in3 => \N__9246\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9026\,
            in1 => \N__8442\,
            in2 => \N__9108\,
            in3 => \N__7170\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11689\,
            ce => \N__5595\,
            sr => \N__11080\
        );

    \U712_REG_SM.STATE_COUNT_RNO_1_2_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__5343\,
            in1 => \N__5609\,
            in2 => \_gnd_net_\,
            in3 => \N__5366\,
            lcout => \U712_REG_SM.N_407\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__10305\,
            in1 => \N__5007\,
            in2 => \N__9852\,
            in3 => \N__5142\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11695\,
            ce => \N__10084\,
            sr => \N__11073\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5085\,
            in2 => \_gnd_net_\,
            in3 => \N__5395\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_455_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__5070\,
            in1 => \N__7017\,
            in2 => \N__5052\,
            in3 => \N__11923\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11700\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5039\,
            in1 => \N__10476\,
            in2 => \_gnd_net_\,
            in3 => \N__9609\,
            lcout => \U712_CHIP_RAM.N_387\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNITI8N_2_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__5652\,
            in1 => \N__5610\,
            in2 => \_gnd_net_\,
            in3 => \N__6821\,
            lcout => \U712_REG_SM.N_406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5651\,
            in2 => \_gnd_net_\,
            in3 => \N__6558\,
            lcout => \U712_REG_SM.N_367\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI902R1_1_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__5336\,
            in1 => \N__5131\,
            in2 => \_gnd_net_\,
            in3 => \N__5359\,
            lcout => \U712_REG_SM.N_185\,
            ltout => \U712_REG_SM.N_185_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11139\,
            in1 => \_gnd_net_\,
            in2 => \N__5154\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.N_185_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_0_1_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__6560\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5649\,
            lcout => \U712_REG_SM.N_368\,
            ltout => \U712_REG_SM.N_368_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_8_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__11922\,
            in1 => \N__5151\,
            in2 => \N__5145\,
            in3 => \N__6606\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6405\,
            in1 => \N__10435\,
            in2 => \_gnd_net_\,
            in3 => \N__10689\,
            lcout => \U712_CHIP_RAM.N_378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIO3HT_8_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5648\,
            in1 => \N__6605\,
            in2 => \_gnd_net_\,
            in3 => \N__6559\,
            lcout => \U712_REG_SM.N_441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_1_1_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__6561\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5650\,
            lcout => \U712_REG_SM.N_358\,
            ltout => \U712_REG_SM.N_358_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010100000"
        )
    port map (
            in0 => \N__11921\,
            in1 => \N__5313\,
            in2 => \N__5115\,
            in3 => \N__6629\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11706\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_1_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__5442\,
            in1 => \N__5112\,
            in2 => \N__9380\,
            in3 => \N__6608\,
            lcout => \U712_REG_SM.REG_CYCLE_5_iv_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNIT80J_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__5415\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5396\,
            lcout => \U712_REG_SM.N_366\,
            ltout => \U712_REG_SM.N_366_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIE5HG1_1_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010001"
        )
    port map (
            in0 => \N__5340\,
            in1 => \N__5662\,
            in2 => \N__5553\,
            in3 => \N__6585\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_1_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40_PLL_derived_clock_RNIIOT_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5541\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_iso_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__5310\,
            in1 => \_gnd_net_\,
            in2 => \N__5452\,
            in3 => \N__6607\,
            lcout => \U712_REG_SM.N_375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNI3OIA1_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5416\,
            in1 => \N__5397\,
            in2 => \_gnd_net_\,
            in3 => \N__5288\,
            lcout => \U712_REG_SM.N_483\,
            ltout => \U712_REG_SM.N_483_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__5341\,
            in1 => \N__11920\,
            in2 => \N__5370\,
            in3 => \N__5367\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11712\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5311\,
            in2 => \_gnd_net_\,
            in3 => \N__5289\,
            lcout => \U712_REG_SM.N_592\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_START_RNO_0_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__11846\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5229\,
            lcout => \U712_CYCLE_TERM.TACK_RST_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__10959\,
            in1 => \N__7731\,
            in2 => \N__7559\,
            in3 => \N__7633\,
            lcout => \U712_REG_SM.N_481\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11975\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9770\,
            in1 => \N__5562\,
            in2 => \N__10518\,
            in3 => \N__7860\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5691\,
            in1 => \N__5760\,
            in2 => \_gnd_net_\,
            in3 => \N__9768\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__9769\,
            in1 => \N__10484\,
            in2 => \N__5670\,
            in3 => \N__9600\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5667\,
            in2 => \_gnd_net_\,
            in3 => \N__6851\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000100010"
        )
    port map (
            in0 => \N__12001\,
            in1 => \N__5619\,
            in2 => \N__5613\,
            in3 => \N__6583\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11693\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6254\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11143\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5583\,
            in1 => \N__5706\,
            in2 => \_gnd_net_\,
            in3 => \N__9738\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__9736\,
            in1 => \N__9970\,
            in2 => \N__9906\,
            in3 => \N__6149\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA25_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11144\,
            in1 => \_gnd_net_\,
            in2 => \N__5556\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA25_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__8694\,
            in1 => \N__5784\,
            in2 => \_gnd_net_\,
            in3 => \N__5792\,
            lcout => \U712_CHIP_RAM.N_499\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10448\,
            in2 => \_gnd_net_\,
            in3 => \N__9737\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_3_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__11999\,
            in1 => \N__12051\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_4_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5793\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12000\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11696\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5778\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11702\,
            ce => \N__8826\,
            sr => \N__11083\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5751\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11702\,
            ce => \N__8826\,
            sr => \N__11083\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__5724\,
            in1 => \N__11400\,
            in2 => \N__6450\,
            in3 => \N__5705\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11708\,
            ce => 'H',
            sr => \N__11076\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011111100"
        )
    port map (
            in0 => \N__6162\,
            in1 => \N__6449\,
            in2 => \N__10485\,
            in3 => \N__6270\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11708\,
            ce => 'H',
            sr => \N__11076\
        );

    \U712_CHIP_RAM.DBENn_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__6255\,
            in1 => \N__6333\,
            in2 => \N__7032\,
            in3 => \N__9444\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11708\,
            ce => 'H',
            sr => \N__11076\
        );

    \U712_REG_SM.LDSn_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__5985\,
            in1 => \N__5957\,
            in2 => \N__6584\,
            in3 => \N__5945\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11708\,
            ce => 'H',
            sr => \N__11076\
        );

    \U712_REG_SM.UDSn_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__5918\,
            in1 => \N__6577\,
            in2 => \N__5946\,
            in3 => \N__6126\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11708\,
            ce => 'H',
            sr => \N__11076\
        );

    \U712_REG_SM.C1_SYNC_1_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6081\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11708\,
            ce => 'H',
            sr => \N__11076\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__6243\,
            in1 => \N__10963\,
            in2 => \_gnd_net_\,
            in3 => \N__9027\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11715\,
            ce => \N__6657\,
            sr => \N__11068\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_0_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001010"
        )
    port map (
            in0 => \N__6312\,
            in1 => \N__5861\,
            in2 => \N__10782\,
            in3 => \N__10466\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_65_i_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100110011"
        )
    port map (
            in0 => \N__10778\,
            in1 => \N__5895\,
            in2 => \N__6353\,
            in3 => \N__8549\,
            lcout => \N_65_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__7827\,
            in1 => \N__5862\,
            in2 => \N__7752\,
            in3 => \N__10467\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_466_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_67_i_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__8550\,
            in1 => \N__6348\,
            in2 => \N__5835\,
            in3 => \N__10893\,
            lcout => \N_67_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6582\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11727\,
            ce => \N__5802\,
            sr => \N__11063\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__7732\,
            in1 => \N__7634\,
            in2 => \N__7560\,
            in3 => \N__10965\,
            lcout => \U712_REG_SM.N_482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_0_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6117\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11735\,
            ce => 'H',
            sr => \N__11062\
        );

    \U712_CHIP_RAM.CAS_COUNTER_0_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__6850\,
            in1 => \N__11995\,
            in2 => \N__6720\,
            in3 => \N__8689\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_RNITKK4_1_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6839\,
            lcout => \DBR_SYNC_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_2_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__8690\,
            in1 => \N__6849\,
            in2 => \N__12006\,
            in3 => \N__6693\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11694\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__8688\,
            in1 => \N__6704\,
            in2 => \N__6750\,
            in3 => \N__6677\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__10292\,
            in1 => \N__9573\,
            in2 => \N__10207\,
            in3 => \N__6072\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11697\,
            ce => \N__10080\,
            sr => \N__11102\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__10194\,
            in1 => \N__10293\,
            in2 => \N__9489\,
            in3 => \N__6042\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11697\,
            ce => \N__10080\,
            sr => \N__11102\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__10294\,
            in1 => \N__9261\,
            in2 => \N__10208\,
            in3 => \N__6012\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11697\,
            ce => \N__10080\,
            sr => \N__11102\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9730\,
            in1 => \N__10590\,
            in2 => \N__9959\,
            in3 => \N__9880\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMER12_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100110111"
        )
    port map (
            in0 => \N__8402\,
            in1 => \N__8163\,
            in2 => \N__8235\,
            in3 => \N__8094\,
            lcout => \U712_CHIP_RAM.N_362\,
            ltout => \U712_CHIP_RAM.N_362_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010100010"
        )
    port map (
            in0 => \N__11991\,
            in1 => \N__8271\,
            in2 => \N__6135\,
            in3 => \N__6774\,
            lcout => \U712_CHIP_RAM.N_435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__8404\,
            in1 => \N__8099\,
            in2 => \N__7989\,
            in3 => \N__8965\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_493_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__7053\,
            in1 => \N__6941\,
            in2 => \N__6132\,
            in3 => \N__9808\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11703\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11145\,
            in2 => \_gnd_net_\,
            in3 => \N__6279\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNIBERN2_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__8164\,
            in1 => \N__8522\,
            in2 => \N__8112\,
            in3 => \N__7238\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_o2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8403\,
            in1 => \N__7100\,
            in2 => \N__7249\,
            in3 => \N__8098\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5V372_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8166\,
            in2 => \_gnd_net_\,
            in3 => \N__7233\,
            lcout => \U712_CHIP_RAM.N_503\,
            ltout => \U712_CHIP_RAM.N_503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__7101\,
            in1 => \_gnd_net_\,
            in2 => \N__6129\,
            in3 => \N__8084\,
            lcout => \U712_CHIP_RAM.N_596\,
            ltout => \U712_CHIP_RAM.N_596_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__7141\,
            in1 => \N__8372\,
            in2 => \N__6282\,
            in3 => \N__6647\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__9085\,
            in1 => \N__9018\,
            in2 => \N__8417\,
            in3 => \N__7139\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNILJ788_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__7140\,
            in1 => \N__8027\,
            in2 => \N__6273\,
            in3 => \N__7102\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__8371\,
            in1 => \N__6269\,
            in2 => \N__6258\,
            in3 => \N__6180\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011000000"
        )
    port map (
            in0 => \N__6239\,
            in1 => \N__11976\,
            in2 => \N__10807\,
            in3 => \N__6197\,
            lcout => \DMA_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11709\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIVFJO_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6179\,
            in2 => \_gnd_net_\,
            in3 => \N__8083\,
            lcout => \U712_CHIP_RAM.N_348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__7314\,
            in1 => \_gnd_net_\,
            in2 => \N__8401\,
            in3 => \N__9092\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa_i_i_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__8757\,
            in1 => \N__8004\,
            in2 => \N__6183\,
            in3 => \N__8970\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11716\,
            ce => \N__9192\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__8346\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6178\,
            lcout => \U712_CHIP_RAM.N_365\,
            ltout => \U712_CHIP_RAM.N_365_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIIFS82_1_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__10389\,
            in1 => \N__8647\,
            in2 => \N__6453\,
            in3 => \N__7047\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIU7TF5_2_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7371\,
            in1 => \N__8347\,
            in2 => \N__9100\,
            in3 => \N__7145\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11142\,
            in1 => \_gnd_net_\,
            in2 => \N__6438\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6435\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11722\,
            ce => \N__8824\,
            sr => \N__11077\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6420\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11722\,
            ce => \N__8824\,
            sr => \N__11077\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6396\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11722\,
            ce => \N__8824\,
            sr => \N__11077\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6381\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11722\,
            ce => \N__8824\,
            sr => \N__11077\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1_0_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6349\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8548\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1Z0Z_0\,
            ltout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a2_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_62_i_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000111"
        )
    port map (
            in0 => \N__6507\,
            in1 => \N__10514\,
            in2 => \N__6306\,
            in3 => \N__10889\,
            lcout => \N_62_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__11140\,
            in1 => \N__7302\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_452_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8239\,
            in1 => \N__7984\,
            in2 => \N__8652\,
            in3 => \N__8423\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6651\,
            in2 => \N__6636\,
            in3 => \N__7158\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_6_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6633\,
            in1 => \N__6615\,
            in2 => \_gnd_net_\,
            in3 => \N__6581\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_445_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100100"
        )
    port map (
            in0 => \N__11930\,
            in1 => \N__9360\,
            in2 => \N__6519\,
            in3 => \N__6516\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11728\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LMBE_0_i_o3_0_o2_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000101111"
        )
    port map (
            in0 => \N__7826\,
            in1 => \N__7748\,
            in2 => \N__7659\,
            in3 => \N__7553\,
            lcout => \U712_BYTE_ENABLE.LMBE_0_i_o3_0_oZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.N_282_i_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__10814\,
            in1 => \N__10869\,
            in2 => \_gnd_net_\,
            in3 => \N__10777\,
            lcout => \N_282_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_0_i_o3_i_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101110000"
        )
    port map (
            in0 => \N__7800\,
            in1 => \N__7736\,
            in2 => \N__7650\,
            in3 => \N__7535\,
            lcout => \N_219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_60_i_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010010101000"
        )
    port map (
            in0 => \N__7536\,
            in1 => \N__7801\,
            in2 => \N__7749\,
            in3 => \N__7641\,
            lcout => \N_60_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_15_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6746\,
            in2 => \N__6735\,
            in3 => \N__6734\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_15_4_0_\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6794\,
            in2 => \_gnd_net_\,
            in3 => \N__6708\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6705\,
            in2 => \_gnd_net_\,
            in3 => \N__6687\,
            lcout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6678\,
            in2 => \_gnd_net_\,
            in3 => \N__6684\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_3_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__11993\,
            in1 => \N__6853\,
            in2 => \N__6681\,
            in3 => \N__8692\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6852\,
            in1 => \N__6666\,
            in2 => \_gnd_net_\,
            in3 => \N__6795\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__11994\,
            in1 => \N__6854\,
            in2 => \N__6660\,
            in3 => \N__8693\,
            lcout => \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_COUNTER_1_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__8691\,
            in1 => \N__6864\,
            in2 => \N__6858\,
            in3 => \N__11992\,
            lcout => \U712_CHIP_RAM.CAS_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11698\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4OVQ3_1_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__6762\,
            in1 => \N__8616\,
            in2 => \N__6786\,
            in3 => \N__11990\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_165_i_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0MGF8_1_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001101"
        )
    port map (
            in0 => \N__11989\,
            in1 => \N__8264\,
            in2 => \N__6777\,
            in3 => \N__6773\,
            lcout => \U712_CHIP_RAM.N_132_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__7377\,
            in1 => \N__6875\,
            in2 => \N__6942\,
            in3 => \N__9893\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__8181\,
            in1 => \N__6940\,
            in2 => \_gnd_net_\,
            in3 => \N__10599\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__6939\,
            in1 => \N__6876\,
            in2 => \N__9969\,
            in3 => \N__8253\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQ8AQ_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8400\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8161\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_i_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8615\,
            in2 => \_gnd_net_\,
            in3 => \N__7950\,
            lcout => \U712_CHIP_RAM.N_510\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__11988\,
            in1 => \N__6756\,
            in2 => \_gnd_net_\,
            in3 => \N__8162\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11704\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI36AQC_2_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__8957\,
            in1 => \N__9101\,
            in2 => \N__8435\,
            in3 => \N__6918\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNINN3QI_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__9017\,
            in1 => \N__8277\,
            in2 => \N__6945\,
            in3 => \N__8958\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__8405\,
            in1 => \N__8626\,
            in2 => \N__8172\,
            in3 => \N__7046\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIEVI78_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__7088\,
            in1 => \N__8956\,
            in2 => \N__6921\,
            in3 => \N__8199\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_ess_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8409\,
            in1 => \N__7089\,
            in2 => \N__7248\,
            in3 => \N__8105\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11710\,
            ce => \N__6894\,
            sr => \N__11103\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0OJB2_7_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__11987\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7234\,
            lcout => \U712_CHIP_RAM.N_577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__8775\,
            in1 => \N__7907\,
            in2 => \N__8796\,
            in3 => \N__8705\,
            lcout => \U712_CHIP_RAM.N_344\,
            ltout => \U712_CHIP_RAM.N_344_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIR80N2_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__11986\,
            in1 => \_gnd_net_\,
            in2 => \N__6885\,
            in3 => \N__8167\,
            lcout => \U712_CHIP_RAM.N_508\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__8568\,
            in1 => \N__6882\,
            in2 => \N__7392\,
            in3 => \N__8754\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11717\,
            ce => \N__9181\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIF4EE6_2_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111000000000"
        )
    port map (
            in0 => \N__7062\,
            in1 => \N__9096\,
            in2 => \N__8426\,
            in3 => \N__8200\,
            lcout => \U712_CHIP_RAM.N_430\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001000100"
        )
    port map (
            in0 => \N__8082\,
            in1 => \N__8622\,
            in2 => \N__7974\,
            in3 => \N__8384\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_0_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7065\,
            in3 => \N__8171\,
            lcout => \U712_CHIP_RAM.N_590\,
            ltout => \U712_CHIP_RAM.N_590_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__8201\,
            in1 => \_gnd_net_\,
            in2 => \N__7056\,
            in3 => \N__8919\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7957\,
            in2 => \_gnd_net_\,
            in3 => \N__8081\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000100"
        )
    port map (
            in0 => \N__9044\,
            in1 => \N__8485\,
            in2 => \N__8468\,
            in3 => \N__9010\,
            lcout => \U712_CHIP_RAM.N_350\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__8646\,
            in1 => \N__7970\,
            in2 => \_gnd_net_\,
            in3 => \N__8080\,
            lcout => \U712_CHIP_RAM.N_509\,
            ltout => \U712_CHIP_RAM.N_509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8430\,
            in2 => \N__7035\,
            in3 => \N__7250\,
            lcout => \U712_CHIP_RAM.DBENn_8_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8487\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10483\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_458_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__11931\,
            in1 => \N__7013\,
            in2 => \N__6981\,
            in3 => \N__6978\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11723\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_0_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9045\,
            in1 => \N__8486\,
            in2 => \N__8469\,
            in3 => \N__9011\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7365\,
            in1 => \N__7349\,
            in2 => \_gnd_net_\,
            in3 => \N__9820\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_1_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7313\,
            in1 => \N__9088\,
            in2 => \N__8434\,
            in3 => \N__7167\,
            lcout => \U712_CHIP_RAM.N_452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7295\,
            in1 => \N__7260\,
            in2 => \_gnd_net_\,
            in3 => \N__9821\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__8425\,
            in1 => \N__8113\,
            in2 => \N__7988\,
            in3 => \N__10510\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CPU_TACK_8_iv_i_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8651\,
            in2 => \N__7254\,
            in3 => \N__7251\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_72_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__7187\,
            in1 => \N__7203\,
            in2 => \N__7197\,
            in3 => \N__7176\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11731\,
            ce => 'H',
            sr => \N__11078\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI1NGC4_2_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7103\,
            in1 => \N__8424\,
            in2 => \N__8247\,
            in3 => \N__7168\,
            lcout => \U712_CHIP_RAM.N_462\,
            ltout => \U712_CHIP_RAM.N_462_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__7169\,
            in1 => \N__8028\,
            in2 => \N__7107\,
            in3 => \N__7104\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__8114\,
            in1 => \N__8547\,
            in2 => \N__7896\,
            in3 => \N__7883\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11731\,
            ce => 'H',
            sr => \N__11078\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__7872\,
            in1 => \N__11304\,
            in2 => \N__10035\,
            in3 => \N__7853\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net\,
            ce => 'H',
            sr => \N__11069\
        );

    \U712_BYTE_ENABLE.N_119_i_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111000000"
        )
    port map (
            in0 => \N__7750\,
            in1 => \N__7802\,
            in2 => \N__7566\,
            in3 => \N__7651\,
            lcout => \N_119_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_61_i_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111010000"
        )
    port map (
            in0 => \N__7803\,
            in1 => \N__7751\,
            in2 => \N__7658\,
            in3 => \N__7565\,
            lcout => \N_61_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_16_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__10301\,
            in1 => \N__11508\,
            in2 => \N__10227\,
            in3 => \N__7422\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11699\,
            ce => \N__10096\,
            sr => \N__11113\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_16_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10529\,
            in1 => \N__7434\,
            in2 => \N__9851\,
            in3 => \N__10680\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_2_0_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8110\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7415\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8625\,
            in1 => \N__8438\,
            in2 => \N__8969\,
            in3 => \N__8111\,
            lcout => \U712_CHIP_RAM.N_431\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000010001"
        )
    port map (
            in0 => \N__8106\,
            in1 => \N__8623\,
            in2 => \_gnd_net_\,
            in3 => \N__7961\,
            lcout => \U712_CHIP_RAM.N_359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIONRK3_1_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8624\,
            in1 => \N__8437\,
            in2 => \_gnd_net_\,
            in3 => \N__8961\,
            lcout => \U712_CHIP_RAM.N_595\,
            ltout => \U712_CHIP_RAM.N_595_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__8121\,
            in1 => \N__8243\,
            in2 => \N__8205\,
            in3 => \N__8202\,
            lcout => \U712_CHIP_RAM.N_279\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8436\,
            in1 => \N__8165\,
            in2 => \N__8115\,
            in3 => \N__7962\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_i_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI6FNG_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8079\,
            in2 => \_gnd_net_\,
            in3 => \N__8521\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0_a2_0\,
            ltout => OPEN,
            carryin => \bfn_16_6_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8742\,
            in1 => \N__8627\,
            in2 => \_gnd_net_\,
            in3 => \N__8007\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__11718\,
            ce => \N__9188\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_2_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8441\,
            in2 => \_gnd_net_\,
            in3 => \N__7992\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8743\,
            in1 => \N__7969\,
            in2 => \_gnd_net_\,
            in3 => \N__7911\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__11718\,
            ce => \N__9188\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8755\,
            in1 => \N__7908\,
            in2 => \_gnd_net_\,
            in3 => \N__8799\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__11718\,
            ce => \N__9188\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8744\,
            in1 => \N__8792\,
            in2 => \_gnd_net_\,
            in3 => \N__8778\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__11718\,
            ce => \N__9188\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8756\,
            in1 => \N__8774\,
            in2 => \_gnd_net_\,
            in3 => \N__8760\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__11718\,
            ce => \N__9188\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8745\,
            in1 => \N__8706\,
            in2 => \_gnd_net_\,
            in3 => \N__8709\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11718\,
            ce => \N__9188\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11912\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9312\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11724\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__8440\,
            in1 => \N__11919\,
            in2 => \_gnd_net_\,
            in3 => \N__8633\,
            lcout => \U712_CHIP_RAM.N_436\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100000"
        )
    port map (
            in0 => \N__8562\,
            in1 => \N__9016\,
            in2 => \N__11973\,
            in3 => \N__8541\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11724\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIHSKQ_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9042\,
            in2 => \_gnd_net_\,
            in3 => \N__8484\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNICG3P2_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__8467\,
            in1 => \N__8439\,
            in2 => \N__8280\,
            in3 => \N__9086\,
            lcout => \U712_CHIP_RAM.N_147_i_i_a2_0\,
            ltout => \U712_CHIP_RAM.N_147_i_i_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIKHPV5_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111111111"
        )
    port map (
            in0 => \N__9015\,
            in1 => \_gnd_net_\,
            in2 => \N__9195\,
            in3 => \N__8960\,
            lcout => \U712_CHIP_RAM.N_500_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__9156\,
            in1 => \N__9135\,
            in2 => \N__11974\,
            in3 => \N__9123\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11724\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__9087\,
            in1 => \N__9043\,
            in2 => \N__9025\,
            in3 => \N__8959\,
            lcout => \U712_CHIP_RAM.N_494\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8913\,
            in1 => \N__9823\,
            in2 => \_gnd_net_\,
            in3 => \N__8859\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9822\,
            in1 => \N__8892\,
            in2 => \_gnd_net_\,
            in3 => \N__8832\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__10468\,
            in1 => \N__9824\,
            in2 => \N__8877\,
            in3 => \N__12063\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8874\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11729\,
            ce => \N__8825\,
            sr => \N__11097\
        );

    \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8853\,
            lcout => \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11729\,
            ce => \N__8825\,
            sr => \N__11097\
        );

    \U712_BUFFERS.N_207_i_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__10881\,
            in1 => \N__10770\,
            in2 => \N__10517\,
            in3 => \N__9379\,
            lcout => \N_207_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__10882\,
            in1 => \N__11911\,
            in2 => \_gnd_net_\,
            in3 => \N__10771\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__9303\,
            in1 => \_gnd_net_\,
            in2 => \N__9279\,
            in3 => \N__9825\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__9267\,
            in1 => \N__10494\,
            in2 => \N__9848\,
            in3 => \N__10614\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9527\,
            in1 => \N__10030\,
            in2 => \_gnd_net_\,
            in3 => \N__11395\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11207\,
            ce => \N__11176\,
            sr => \N__11084\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10026\,
            in1 => \N__9528\,
            in2 => \_gnd_net_\,
            in3 => \N__11298\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__11174\,
            sr => \N__11079\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__10290\,
            in1 => \N__9582\,
            in2 => \N__10228\,
            in3 => \N__9231\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11730\,
            ce => \N__10098\,
            sr => \N__11105\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10474\,
            in1 => \N__9207\,
            in2 => \N__9849\,
            in3 => \N__9588\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10475\,
            in1 => \N__9201\,
            in2 => \N__9850\,
            in3 => \N__10665\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9558\,
            in1 => \N__11394\,
            in2 => \_gnd_net_\,
            in3 => \N__9516\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__11178\,
            sr => \N__11098\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9557\,
            in1 => \N__11393\,
            in2 => \_gnd_net_\,
            in3 => \N__11448\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__11178\,
            sr => \N__11098\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__10654\,
            in1 => \_gnd_net_\,
            in2 => \N__9474\,
            in3 => \N__11385\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11205\,
            ce => \N__11177\,
            sr => \N__11092\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11439\,
            in1 => \N__11386\,
            in2 => \_gnd_net_\,
            in3 => \N__9547\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11205\,
            ce => \N__11177\,
            sr => \N__11092\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9548\,
            in1 => \_gnd_net_\,
            in2 => \N__11396\,
            in3 => \N__9526\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11205\,
            ce => \N__11177\,
            sr => \N__11092\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11297\,
            in1 => \N__10653\,
            in2 => \_gnd_net_\,
            in3 => \N__9473\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__11175\,
            sr => \N__11085\
        );

    \U712_CHIP_RAM.RASn_LC_18_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9905\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11705\,
            ce => 'H',
            sr => \N__11118\
        );

    \U712_CHIP_RAM.CRCSn_LC_18_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9971\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11711\,
            ce => 'H',
            sr => \N__11116\
        );

    \U712_CHIP_RAM.CASn_LC_18_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9847\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11711\,
            ce => 'H',
            sr => \N__11116\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_18_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__10266\,
            in1 => \N__9975\,
            in2 => \_gnd_net_\,
            in3 => \N__9846\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11719\,
            ce => \N__10113\,
            sr => \N__11115\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_18_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__10601\,
            in1 => \N__9898\,
            in2 => \_gnd_net_\,
            in3 => \N__9845\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_18_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9897\,
            in2 => \_gnd_net_\,
            in3 => \N__10600\,
            lcout => \U712_CHIP_RAM.N_354\,
            ltout => \U712_CHIP_RAM.N_354_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_18_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__10500\,
            in1 => \N__11232\,
            in2 => \N__9855\,
            in3 => \N__9844\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_18_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001010101"
        )
    port map (
            in0 => \N__10265\,
            in1 => \N__11231\,
            in2 => \N__10528\,
            in3 => \N__9837\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9681\,
            in1 => \N__9672\,
            in2 => \_gnd_net_\,
            in3 => \N__9666\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11733\,
            ce => \N__10108\,
            sr => \N__11108\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__10289\,
            in1 => \N__9615\,
            in2 => \N__10230\,
            in3 => \N__9639\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11733\,
            ce => \N__10108\,
            sr => \N__11108\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12105\,
            in1 => \N__11378\,
            in2 => \_gnd_net_\,
            in3 => \N__11585\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11208\,
            ce => \N__11180\,
            sr => \N__11106\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10659\,
            in1 => \N__11377\,
            in2 => \_gnd_net_\,
            in3 => \N__11543\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11208\,
            ce => \N__11180\,
            sr => \N__11106\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__11542\,
            in1 => \_gnd_net_\,
            in2 => \N__11383\,
            in3 => \N__11583\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__11179\,
            sr => \N__11104\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11584\,
            in1 => \N__11356\,
            in2 => \_gnd_net_\,
            in3 => \N__12102\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__11179\,
            sr => \N__11104\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__12103\,
            in1 => \_gnd_net_\,
            in2 => \N__11384\,
            in3 => \N__11495\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__11179\,
            sr => \N__11104\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10658\,
            in1 => \N__11352\,
            in2 => \_gnd_net_\,
            in3 => \N__11541\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__11179\,
            sr => \N__11104\
        );

    \U712_CHIP_RAM.WEn_LC_19_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10605\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11725\,
            ce => 'H',
            sr => \N__11117\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_19_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__10554\,
            in1 => \N__10548\,
            in2 => \N__10530\,
            in3 => \N__9984\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11734\,
            ce => \N__10097\,
            sr => \N__11114\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__10291\,
            in1 => \N__12069\,
            in2 => \N__10229\,
            in3 => \N__10146\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11736\,
            ce => \N__10112\,
            sr => \N__11111\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_19_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11376\,
            in1 => \N__12035\,
            in2 => \_gnd_net_\,
            in3 => \N__10034\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11206\,
            ce => \N__11182\,
            sr => \N__11109\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11496\,
            in1 => \N__11375\,
            in2 => \_gnd_net_\,
            in3 => \N__12104\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11206\,
            ce => \N__11182\,
            sr => \N__11109\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11494\,
            in1 => \N__11351\,
            in2 => \_gnd_net_\,
            in3 => \N__11447\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4C_net\,
            ce => \N__11181\,
            sr => \N__11107\
        );

    \U712_CHIP_RAM.RAS_SYNC_2_LC_20_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11834\,
            in2 => \_gnd_net_\,
            in3 => \N__11748\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11737\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_20_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__12042\,
            in1 => \N__11832\,
            in2 => \_gnd_net_\,
            in3 => \N__12018\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_20_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11833\,
            in2 => \_gnd_net_\,
            in3 => \N__11754\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_20_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11589\,
            in1 => \N__11379\,
            in2 => \_gnd_net_\,
            in3 => \N__11550\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11204\,
            ce => \N__11184\,
            sr => \N__11112\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11493\,
            in1 => \N__11440\,
            in2 => \_gnd_net_\,
            in3 => \N__11350\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11203\,
            ce => \N__11183\,
            sr => \N__11110\
        );

    \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_24_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100001111"
        )
    port map (
            in0 => \N__10964\,
            in1 => \N__10857\,
            in2 => \N__10821\,
            in3 => \N__10746\,
            lcout => \N_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Apr 7 2025 15:46:56

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U409_TOP" view "INTERFACE"

module U409_TOP (
    TM,
    TT,
    D,
    A,
    TICK60,
    CIACS0n,
    CLK6,
    CLK_CIA,
    BUFENn,
    CIACS1n,
    TICK50,
    RAMSPACEn,
    CLK40_IN,
    CLK28_IN,
    REGSPACEn,
    TSn,
    RTC_ENn,
    RESETn,
    OVL,
    TACKn,
    ROMENn,
    PORTSIZE);

    input [1:0] TM;
    input [1:0] TT;
    output [7:0] D;
    input [31:1] A;
    output TICK60;
    output CIACS0n;
    input CLK6;
    output CLK_CIA;
    output BUFENn;
    output CIACS1n;
    output TICK50;
    output RAMSPACEn;
    input CLK40_IN;
    input CLK28_IN;
    output REGSPACEn;
    input TSn;
    output RTC_ENn;
    input RESETn;
    input OVL;
    inout TACKn;
    output ROMENn;
    output PORTSIZE;

    wire N__7375;
    wire N__7374;
    wire N__7373;
    wire N__7365;
    wire N__7364;
    wire N__7363;
    wire N__7354;
    wire N__7353;
    wire N__7352;
    wire N__7345;
    wire N__7344;
    wire N__7343;
    wire N__7336;
    wire N__7335;
    wire N__7334;
    wire N__7327;
    wire N__7326;
    wire N__7325;
    wire N__7318;
    wire N__7317;
    wire N__7316;
    wire N__7309;
    wire N__7308;
    wire N__7307;
    wire N__7300;
    wire N__7299;
    wire N__7298;
    wire N__7291;
    wire N__7290;
    wire N__7289;
    wire N__7282;
    wire N__7281;
    wire N__7280;
    wire N__7273;
    wire N__7272;
    wire N__7271;
    wire N__7264;
    wire N__7263;
    wire N__7262;
    wire N__7255;
    wire N__7254;
    wire N__7253;
    wire N__7246;
    wire N__7245;
    wire N__7244;
    wire N__7237;
    wire N__7236;
    wire N__7235;
    wire N__7228;
    wire N__7227;
    wire N__7226;
    wire N__7219;
    wire N__7218;
    wire N__7217;
    wire N__7210;
    wire N__7209;
    wire N__7208;
    wire N__7201;
    wire N__7200;
    wire N__7199;
    wire N__7192;
    wire N__7191;
    wire N__7190;
    wire N__7183;
    wire N__7182;
    wire N__7181;
    wire N__7174;
    wire N__7173;
    wire N__7172;
    wire N__7165;
    wire N__7164;
    wire N__7163;
    wire N__7156;
    wire N__7155;
    wire N__7154;
    wire N__7147;
    wire N__7146;
    wire N__7145;
    wire N__7138;
    wire N__7137;
    wire N__7136;
    wire N__7129;
    wire N__7128;
    wire N__7127;
    wire N__7120;
    wire N__7119;
    wire N__7118;
    wire N__7111;
    wire N__7110;
    wire N__7109;
    wire N__7102;
    wire N__7101;
    wire N__7100;
    wire N__7093;
    wire N__7092;
    wire N__7091;
    wire N__7084;
    wire N__7083;
    wire N__7082;
    wire N__7075;
    wire N__7074;
    wire N__7073;
    wire N__7066;
    wire N__7065;
    wire N__7064;
    wire N__7057;
    wire N__7056;
    wire N__7055;
    wire N__7048;
    wire N__7047;
    wire N__7046;
    wire N__7039;
    wire N__7038;
    wire N__7037;
    wire N__7030;
    wire N__7029;
    wire N__7028;
    wire N__7021;
    wire N__7020;
    wire N__7019;
    wire N__7012;
    wire N__7011;
    wire N__7010;
    wire N__7003;
    wire N__7002;
    wire N__7001;
    wire N__6994;
    wire N__6993;
    wire N__6992;
    wire N__6985;
    wire N__6984;
    wire N__6983;
    wire N__6976;
    wire N__6975;
    wire N__6974;
    wire N__6967;
    wire N__6966;
    wire N__6965;
    wire N__6958;
    wire N__6957;
    wire N__6956;
    wire N__6949;
    wire N__6948;
    wire N__6947;
    wire N__6930;
    wire N__6927;
    wire N__6924;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6912;
    wire N__6911;
    wire N__6910;
    wire N__6909;
    wire N__6908;
    wire N__6907;
    wire N__6906;
    wire N__6905;
    wire N__6894;
    wire N__6887;
    wire N__6882;
    wire N__6881;
    wire N__6880;
    wire N__6879;
    wire N__6878;
    wire N__6877;
    wire N__6876;
    wire N__6875;
    wire N__6866;
    wire N__6857;
    wire N__6852;
    wire N__6849;
    wire N__6846;
    wire N__6843;
    wire N__6840;
    wire N__6839;
    wire N__6838;
    wire N__6837;
    wire N__6836;
    wire N__6835;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6820;
    wire N__6819;
    wire N__6816;
    wire N__6813;
    wire N__6808;
    wire N__6799;
    wire N__6792;
    wire N__6789;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6777;
    wire N__6776;
    wire N__6775;
    wire N__6774;
    wire N__6773;
    wire N__6772;
    wire N__6771;
    wire N__6770;
    wire N__6769;
    wire N__6750;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6732;
    wire N__6729;
    wire N__6726;
    wire N__6723;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6708;
    wire N__6705;
    wire N__6702;
    wire N__6699;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6687;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6675;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6663;
    wire N__6662;
    wire N__6659;
    wire N__6656;
    wire N__6655;
    wire N__6650;
    wire N__6647;
    wire N__6642;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6615;
    wire N__6614;
    wire N__6611;
    wire N__6608;
    wire N__6603;
    wire N__6600;
    wire N__6597;
    wire N__6594;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6582;
    wire N__6579;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6567;
    wire N__6564;
    wire N__6561;
    wire N__6558;
    wire N__6557;
    wire N__6554;
    wire N__6551;
    wire N__6546;
    wire N__6545;
    wire N__6542;
    wire N__6539;
    wire N__6534;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6501;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6489;
    wire N__6486;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6465;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6441;
    wire N__6440;
    wire N__6437;
    wire N__6434;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6422;
    wire N__6419;
    wire N__6416;
    wire N__6411;
    wire N__6410;
    wire N__6409;
    wire N__6408;
    wire N__6405;
    wire N__6398;
    wire N__6395;
    wire N__6390;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6378;
    wire N__6375;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6363;
    wire N__6362;
    wire N__6359;
    wire N__6356;
    wire N__6351;
    wire N__6348;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6336;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6312;
    wire N__6309;
    wire N__6306;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6294;
    wire N__6291;
    wire N__6288;
    wire N__6285;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6273;
    wire N__6270;
    wire N__6267;
    wire N__6264;
    wire N__6261;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6249;
    wire N__6246;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6234;
    wire N__6231;
    wire N__6230;
    wire N__6227;
    wire N__6224;
    wire N__6219;
    wire N__6216;
    wire N__6213;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6193;
    wire N__6190;
    wire N__6187;
    wire N__6184;
    wire N__6177;
    wire N__6176;
    wire N__6175;
    wire N__6174;
    wire N__6171;
    wire N__6164;
    wire N__6161;
    wire N__6156;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6144;
    wire N__6141;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6129;
    wire N__6126;
    wire N__6125;
    wire N__6122;
    wire N__6119;
    wire N__6114;
    wire N__6111;
    wire N__6108;
    wire N__6105;
    wire N__6102;
    wire N__6099;
    wire N__6096;
    wire N__6093;
    wire N__6090;
    wire N__6087;
    wire N__6084;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6063;
    wire N__6060;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6038;
    wire N__6037;
    wire N__6036;
    wire N__6035;
    wire N__6034;
    wire N__6033;
    wire N__6030;
    wire N__6023;
    wire N__6016;
    wire N__6009;
    wire N__6008;
    wire N__6007;
    wire N__6006;
    wire N__6005;
    wire N__6002;
    wire N__6001;
    wire N__6000;
    wire N__5997;
    wire N__5990;
    wire N__5983;
    wire N__5976;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5968;
    wire N__5967;
    wire N__5966;
    wire N__5965;
    wire N__5964;
    wire N__5961;
    wire N__5956;
    wire N__5947;
    wire N__5944;
    wire N__5937;
    wire N__5934;
    wire N__5933;
    wire N__5932;
    wire N__5931;
    wire N__5930;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5912;
    wire N__5907;
    wire N__5906;
    wire N__5905;
    wire N__5904;
    wire N__5903;
    wire N__5900;
    wire N__5891;
    wire N__5886;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5878;
    wire N__5877;
    wire N__5874;
    wire N__5871;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5848;
    wire N__5847;
    wire N__5846;
    wire N__5839;
    wire N__5838;
    wire N__5837;
    wire N__5832;
    wire N__5829;
    wire N__5828;
    wire N__5827;
    wire N__5826;
    wire N__5823;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5794;
    wire N__5789;
    wire N__5788;
    wire N__5785;
    wire N__5780;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5727;
    wire N__5724;
    wire N__5723;
    wire N__5722;
    wire N__5721;
    wire N__5718;
    wire N__5711;
    wire N__5706;
    wire N__5703;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5690;
    wire N__5689;
    wire N__5686;
    wire N__5683;
    wire N__5682;
    wire N__5681;
    wire N__5678;
    wire N__5677;
    wire N__5672;
    wire N__5669;
    wire N__5662;
    wire N__5655;
    wire N__5654;
    wire N__5653;
    wire N__5652;
    wire N__5651;
    wire N__5650;
    wire N__5649;
    wire N__5646;
    wire N__5639;
    wire N__5632;
    wire N__5625;
    wire N__5624;
    wire N__5623;
    wire N__5622;
    wire N__5621;
    wire N__5620;
    wire N__5619;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5601;
    wire N__5592;
    wire N__5591;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5583;
    wire N__5580;
    wire N__5575;
    wire N__5572;
    wire N__5571;
    wire N__5568;
    wire N__5563;
    wire N__5560;
    wire N__5555;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5532;
    wire N__5529;
    wire N__5528;
    wire N__5525;
    wire N__5524;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5496;
    wire N__5495;
    wire N__5494;
    wire N__5491;
    wire N__5490;
    wire N__5487;
    wire N__5482;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5457;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5436;
    wire N__5435;
    wire N__5434;
    wire N__5433;
    wire N__5432;
    wire N__5431;
    wire N__5430;
    wire N__5427;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5403;
    wire N__5402;
    wire N__5397;
    wire N__5394;
    wire N__5393;
    wire N__5392;
    wire N__5389;
    wire N__5384;
    wire N__5379;
    wire N__5376;
    wire N__5373;
    wire N__5370;
    wire N__5367;
    wire N__5364;
    wire N__5363;
    wire N__5362;
    wire N__5359;
    wire N__5358;
    wire N__5355;
    wire N__5352;
    wire N__5351;
    wire N__5348;
    wire N__5345;
    wire N__5340;
    wire N__5337;
    wire N__5332;
    wire N__5327;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5309;
    wire N__5308;
    wire N__5305;
    wire N__5300;
    wire N__5295;
    wire N__5292;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5280;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5265;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5205;
    wire N__5202;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5184;
    wire N__5181;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5168;
    wire N__5163;
    wire N__5160;
    wire N__5157;
    wire N__5156;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5146;
    wire N__5139;
    wire N__5138;
    wire N__5137;
    wire N__5136;
    wire N__5133;
    wire N__5126;
    wire N__5121;
    wire N__5120;
    wire N__5119;
    wire N__5118;
    wire N__5115;
    wire N__5112;
    wire N__5107;
    wire N__5100;
    wire N__5099;
    wire N__5098;
    wire N__5095;
    wire N__5090;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5076;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire N__5068;
    wire N__5067;
    wire N__5062;
    wire N__5057;
    wire N__5052;
    wire N__5051;
    wire N__5050;
    wire N__5049;
    wire N__5048;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5034;
    wire N__5029;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5013;
    wire N__5012;
    wire N__5007;
    wire N__5004;
    wire N__5001;
    wire N__4998;
    wire N__4995;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4987;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4931;
    wire N__4930;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4908;
    wire N__4905;
    wire N__4904;
    wire N__4903;
    wire N__4900;
    wire N__4897;
    wire N__4894;
    wire N__4887;
    wire N__4884;
    wire N__4881;
    wire N__4878;
    wire N__4877;
    wire N__4876;
    wire N__4873;
    wire N__4868;
    wire N__4863;
    wire N__4862;
    wire N__4861;
    wire N__4858;
    wire N__4857;
    wire N__4852;
    wire N__4847;
    wire N__4842;
    wire N__4839;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4823;
    wire N__4822;
    wire N__4817;
    wire N__4816;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4800;
    wire N__4799;
    wire N__4798;
    wire N__4793;
    wire N__4790;
    wire N__4785;
    wire N__4784;
    wire N__4783;
    wire N__4782;
    wire N__4781;
    wire N__4780;
    wire N__4775;
    wire N__4772;
    wire N__4765;
    wire N__4758;
    wire N__4757;
    wire N__4756;
    wire N__4753;
    wire N__4750;
    wire N__4749;
    wire N__4746;
    wire N__4739;
    wire N__4734;
    wire N__4733;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4716;
    wire N__4715;
    wire N__4714;
    wire N__4713;
    wire N__4712;
    wire N__4711;
    wire N__4704;
    wire N__4697;
    wire N__4694;
    wire N__4689;
    wire N__4688;
    wire N__4687;
    wire N__4686;
    wire N__4683;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4675;
    wire N__4668;
    wire N__4661;
    wire N__4656;
    wire N__4655;
    wire N__4654;
    wire N__4653;
    wire N__4652;
    wire N__4647;
    wire N__4640;
    wire N__4635;
    wire N__4634;
    wire N__4633;
    wire N__4632;
    wire N__4631;
    wire N__4628;
    wire N__4621;
    wire N__4618;
    wire N__4611;
    wire N__4610;
    wire N__4609;
    wire N__4606;
    wire N__4605;
    wire N__4604;
    wire N__4601;
    wire N__4594;
    wire N__4591;
    wire N__4584;
    wire N__4583;
    wire N__4582;
    wire N__4581;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4565;
    wire N__4564;
    wire N__4563;
    wire N__4560;
    wire N__4557;
    wire N__4554;
    wire N__4551;
    wire N__4542;
    wire N__4541;
    wire N__4540;
    wire N__4539;
    wire N__4538;
    wire N__4537;
    wire N__4534;
    wire N__4531;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4506;
    wire N__4505;
    wire N__4504;
    wire N__4503;
    wire N__4500;
    wire N__4497;
    wire N__4494;
    wire N__4491;
    wire N__4488;
    wire N__4485;
    wire N__4476;
    wire N__4475;
    wire N__4474;
    wire N__4473;
    wire N__4468;
    wire N__4465;
    wire N__4464;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4437;
    wire N__4434;
    wire N__4431;
    wire N__4428;
    wire N__4425;
    wire N__4424;
    wire N__4421;
    wire N__4420;
    wire N__4417;
    wire N__4416;
    wire N__4415;
    wire N__4412;
    wire N__4407;
    wire N__4404;
    wire N__4401;
    wire N__4392;
    wire N__4389;
    wire N__4386;
    wire N__4383;
    wire N__4382;
    wire N__4381;
    wire N__4380;
    wire N__4379;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4349;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4323;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4311;
    wire N__4308;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4287;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4275;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4263;
    wire N__4260;
    wire N__4257;
    wire N__4254;
    wire N__4251;
    wire N__4248;
    wire N__4245;
    wire N__4242;
    wire N__4239;
    wire N__4238;
    wire N__4235;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4217;
    wire N__4212;
    wire N__4209;
    wire N__4208;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4167;
    wire N__4164;
    wire N__4161;
    wire N__4158;
    wire N__4155;
    wire N__4152;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4140;
    wire N__4137;
    wire N__4134;
    wire N__4131;
    wire N__4128;
    wire N__4125;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4107;
    wire N__4104;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4092;
    wire N__4089;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4050;
    wire N__4047;
    wire N__4044;
    wire N__4041;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4029;
    wire N__4026;
    wire N__4023;
    wire N__4020;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4007;
    wire N__4002;
    wire N__3999;
    wire N__3996;
    wire N__3993;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3981;
    wire N__3980;
    wire N__3979;
    wire N__3978;
    wire N__3977;
    wire N__3976;
    wire N__3975;
    wire N__3972;
    wire N__3965;
    wire N__3964;
    wire N__3963;
    wire N__3960;
    wire N__3955;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3939;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3921;
    wire N__3918;
    wire N__3915;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3902;
    wire N__3901;
    wire N__3900;
    wire N__3899;
    wire N__3898;
    wire N__3895;
    wire N__3894;
    wire N__3889;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3877;
    wire N__3876;
    wire N__3875;
    wire N__3872;
    wire N__3865;
    wire N__3862;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3845;
    wire N__3838;
    wire N__3835;
    wire N__3830;
    wire N__3825;
    wire N__3824;
    wire N__3823;
    wire N__3820;
    wire N__3819;
    wire N__3818;
    wire N__3817;
    wire N__3816;
    wire N__3813;
    wire N__3808;
    wire N__3807;
    wire N__3806;
    wire N__3805;
    wire N__3802;
    wire N__3799;
    wire N__3794;
    wire N__3791;
    wire N__3788;
    wire N__3783;
    wire N__3780;
    wire N__3773;
    wire N__3764;
    wire N__3761;
    wire N__3758;
    wire N__3753;
    wire N__3750;
    wire N__3747;
    wire N__3744;
    wire N__3741;
    wire N__3738;
    wire N__3735;
    wire N__3732;
    wire N__3729;
    wire N__3726;
    wire N__3723;
    wire N__3720;
    wire N__3717;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3695;
    wire N__3694;
    wire N__3689;
    wire N__3686;
    wire N__3685;
    wire N__3684;
    wire N__3681;
    wire N__3678;
    wire N__3675;
    wire N__3672;
    wire N__3669;
    wire N__3666;
    wire N__3663;
    wire N__3660;
    wire N__3659;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3630;
    wire N__3627;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3615;
    wire N__3612;
    wire N__3609;
    wire N__3608;
    wire N__3607;
    wire N__3606;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3596;
    wire N__3595;
    wire N__3588;
    wire N__3585;
    wire N__3582;
    wire N__3579;
    wire N__3576;
    wire N__3571;
    wire N__3568;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3552;
    wire N__3549;
    wire N__3548;
    wire N__3547;
    wire N__3546;
    wire N__3545;
    wire N__3540;
    wire N__3537;
    wire N__3534;
    wire N__3533;
    wire N__3530;
    wire N__3525;
    wire N__3522;
    wire N__3519;
    wire N__3516;
    wire N__3509;
    wire N__3506;
    wire N__3503;
    wire N__3500;
    wire N__3497;
    wire N__3494;
    wire N__3489;
    wire N__3486;
    wire N__3483;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3471;
    wire N__3468;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3456;
    wire N__3455;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3438;
    wire N__3435;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3427;
    wire N__3426;
    wire N__3423;
    wire N__3420;
    wire N__3417;
    wire N__3414;
    wire N__3413;
    wire N__3412;
    wire N__3407;
    wire N__3402;
    wire N__3397;
    wire N__3396;
    wire N__3393;
    wire N__3388;
    wire N__3385;
    wire N__3378;
    wire N__3375;
    wire N__3372;
    wire N__3369;
    wire N__3366;
    wire N__3365;
    wire N__3362;
    wire N__3361;
    wire N__3358;
    wire N__3357;
    wire N__3356;
    wire N__3353;
    wire N__3350;
    wire N__3347;
    wire N__3344;
    wire N__3341;
    wire N__3336;
    wire N__3329;
    wire N__3326;
    wire N__3323;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3309;
    wire N__3306;
    wire N__3305;
    wire N__3304;
    wire N__3299;
    wire N__3296;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3281;
    wire N__3280;
    wire N__3279;
    wire N__3274;
    wire N__3269;
    wire N__3264;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3248;
    wire N__3247;
    wire N__3240;
    wire N__3237;
    wire N__3234;
    wire N__3231;
    wire N__3228;
    wire N__3225;
    wire N__3222;
    wire N__3219;
    wire N__3216;
    wire N__3215;
    wire N__3212;
    wire N__3209;
    wire N__3204;
    wire N__3203;
    wire N__3200;
    wire N__3197;
    wire N__3192;
    wire N__3189;
    wire N__3186;
    wire N__3183;
    wire N__3182;
    wire N__3179;
    wire N__3176;
    wire N__3173;
    wire N__3170;
    wire N__3167;
    wire N__3164;
    wire N__3161;
    wire N__3156;
    wire N__3153;
    wire N__3150;
    wire N__3147;
    wire N__3144;
    wire N__3141;
    wire N__3138;
    wire N__3135;
    wire N__3132;
    wire N__3129;
    wire N__3126;
    wire N__3123;
    wire N__3120;
    wire N__3117;
    wire N__3114;
    wire N__3111;
    wire N__3110;
    wire N__3105;
    wire N__3102;
    wire N__3099;
    wire N__3096;
    wire N__3093;
    wire N__3092;
    wire N__3087;
    wire N__3084;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3072;
    wire N__3069;
    wire N__3066;
    wire N__3063;
    wire N__3062;
    wire N__3057;
    wire N__3054;
    wire N__3051;
    wire N__3048;
    wire N__3045;
    wire N__3042;
    wire N__3041;
    wire N__3036;
    wire N__3033;
    wire N__3030;
    wire N__3027;
    wire N__3024;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3009;
    wire N__3006;
    wire N__3003;
    wire N__3000;
    wire N__2999;
    wire N__2994;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire N__2979;
    wire N__2976;
    wire N__2975;
    wire N__2970;
    wire N__2967;
    wire N__2964;
    wire N__2961;
    wire N__2958;
    wire N__2955;
    wire N__2954;
    wire N__2949;
    wire N__2946;
    wire N__2943;
    wire N__2940;
    wire N__2937;
    wire N__2934;
    wire N__2931;
    wire N__2928;
    wire N__2925;
    wire N__2922;
    wire N__2919;
    wire N__2916;
    wire N__2913;
    wire N__2910;
    wire N__2909;
    wire N__2904;
    wire N__2901;
    wire N__2900;
    wire N__2899;
    wire N__2898;
    wire N__2897;
    wire N__2896;
    wire N__2895;
    wire N__2894;
    wire N__2893;
    wire N__2892;
    wire N__2891;
    wire N__2868;
    wire CLK80_OUT;
    wire GNDG0;
    wire VCCG0;
    wire A_c_31;
    wire A_c_30;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_ ;
    wire A_c_26;
    wire A_c_24;
    wire A_c_27;
    wire A_c_25;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_3 ;
    wire A_c_29;
    wire \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_4_cascade_ ;
    wire A_c_28;
    wire U409_ADDRESS_DECODE_un1_RTC_ENn_i;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_1 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_1_cascade_ ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3 ;
    wire A_c_16;
    wire A_c_17;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3_cascade_ ;
    wire U409_ADDRESS_DECODE_AUTOVECTOR_5_cascade_;
    wire A_c_18;
    wire \U409_ADDRESS_DECODE.AUTOVECTOR_16 ;
    wire TT_c_1;
    wire TT_c_0;
    wire U409_ADDRESS_DECODE_AUTOVECTOR_4;
    wire \U409_TRANSFER_ACK.N_38 ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3Z0Z_2_cascade_ ;
    wire \U409_ADDRESS_DECODE.CIA_SPACE_6 ;
    wire \U409_ADDRESS_DECODE.un1_RTC_ENn_2_cascade_ ;
    wire A_c_20;
    wire \U409_ADDRESS_DECODE.REGISTER_SPACEZ0 ;
    wire \U409_ADDRESS_DECODE.RANGER_SPACEZ0Z_2_cascade_ ;
    wire A_c_19;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ;
    wire \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1 ;
    wire OVL_c;
    wire \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0_cascade_ ;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn_i;
    wire U409_ADDRESS_DECODE_un1_RTC_ENn;
    wire PORTSIZE_0_i;
    wire A_c_23;
    wire \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0 ;
    wire A_c_22;
    wire A_c_21;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn_cascade_;
    wire U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_5;
    wire U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_7;
    wire AGNUS_SPACE_0_cascade_;
    wire U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_6;
    wire BUFENn_c;
    wire TM_c_0;
    wire \U409_ADDRESS_DECODE.un2_REGSPACEn_0 ;
    wire \U409_ADDRESS_DECODE.Z2_SPACEZ0 ;
    wire TM_c_1;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn_i;
    wire CIA_SPACE;
    wire \U409_CIA.VMA_RNOZ0Z_0_cascade_ ;
    wire \U409_CIA.un1_CIA_CLK_COUNT_3_1 ;
    wire bfn_9_8_0_;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_1 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_3 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_5 ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_6 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ;
    wire U409_ADDRESS_DECODE_un1_REGSPACEn;
    wire U409_ADDRESS_DECODE_un1_RAMSPACEn;
    wire TACKn_in;
    wire A_c_13;
    wire U409_ADDRESS_DECODE_un1_CIACS1n_i;
    wire A_c_12;
    wire U409_ADDRESS_DECODE_un1_CIACS0n_i;
    wire CIA_ENABLE;
    wire \U409_CIA.CLK_CIA6_0 ;
    wire \U409_CIA.CLK_CIA6_cascade_ ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_0 ;
    wire \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ;
    wire \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO ;
    wire \U409_CIA.CIA_CLK_COUNT11_3 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_2 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_5 ;
    wire CLK28_IN_c_g;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_6 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_0 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_7 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_1 ;
    wire \U409_CIA.CLK_CIA6_3 ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_4 ;
    wire \U409_CIA.un1_CIA_CLK_COUNT_2_1 ;
    wire \U409_CIA.CLK_CIA6_3_cascade_ ;
    wire \U409_CIA.CIA_CLK_COUNTZ0Z_3 ;
    wire \U409_CIA.CLK_CIA_RNOZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_6_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ;
    wire \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ;
    wire \U409_TRANSFER_ACK.m8_ns_1_cascade_ ;
    wire \U409_TRANSFER_ACK.i6_mux_0_cascade_ ;
    wire \U409_TRANSFER_ACK.N_9 ;
    wire \INVU409_TRANSFER_ACK.CIA_STATE_1C_net ;
    wire \U409_TRANSFER_ACK.N_4 ;
    wire \U409_TRANSFER_ACK.N_4_cascade_ ;
    wire \U409_TRANSFER_ACK.N_5 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ;
    wire CLK_CIA_c;
    wire \U409_CIA.VMAZ0 ;
    wire \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ;
    wire \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_0 ;
    wire \U409_TRANSFER_ACK.LASTCLKZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_EN_e_1 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ;
    wire \U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ;
    wire \U409_TRANSFER_ACK.N_138 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_0 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_cascade_ ;
    wire \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_ENZ0 ;
    wire \U409_TRANSFER_ACK.CIA_TACK_ENZ0 ;
    wire CONSTANT_ONE_NET;
    wire \U409_TRANSFER_ACK.N_18 ;
    wire \U409_TRANSFER_ACK.N_24 ;
    wire \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_0 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ;
    wire ROMENn_c;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ;
    wire \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ;
    wire TSn_c;
    wire U409_ADDRESS_DECODE_ROMEN_1;
    wire CLK40_IN_c;
    wire \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ;
    wire \U409_TRANSFER_ACK.N_28_4 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ;
    wire \INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC_net ;
    wire \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_0 ;
    wire RESETn_c_i;
    wire \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ;
    wire TACK_OUTn;
    wire \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ;
    wire \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ;
    wire RESETn_c;
    wire \U409_TRANSFER_ACK.TACK_COUNTER6 ;
    wire \INVU409_TRANSFER_ACK.TACK_EN_iC_net ;
    wire \U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en ;
    wire \U409_TICK.TICK603_8_cascade_ ;
    wire \U409_TICK.TICK603_14_cascade_ ;
    wire \U409_TICK.TICK603_9_cascade_ ;
    wire TICK60_c;
    wire \U409_TICK.TICK603_10_cascade_ ;
    wire \U409_TICK.TICK603_11 ;
    wire \U409_TICK.TICK603_14 ;
    wire \U409_TICK.TICK603_9 ;
    wire \U409_TICK.TICK603_10 ;
    wire bfn_14_1_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_1 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_2 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_3 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_4 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_5 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_6 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_7 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_8 ;
    wire bfn_14_2_0_;
    wire \U409_TICK.un2_COUNTER50_1_cry_9 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_10 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_11 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_12 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_13 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_14 ;
    wire \U409_TICK.un2_COUNTER50_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_1 ;
    wire \U409_TICK.COUNTER60Z0Z_0 ;
    wire bfn_14_4_0_;
    wire \U409_TICK.COUNTER60Z0Z_2 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_1 ;
    wire \U409_TICK.COUNTER60Z0Z_3 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_2 ;
    wire \U409_TICK.COUNTER60Z0Z_4 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_4 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_3 ;
    wire \U409_TICK.COUNTER60Z0Z_5 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_4 ;
    wire \U409_TICK.COUNTER60Z0Z_6 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_6 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_5 ;
    wire \U409_TICK.COUNTER60Z0Z_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_6 ;
    wire \U409_TICK.COUNTER60Z0Z_8 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_8 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_7 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_8 ;
    wire \U409_TICK.COUNTER60Z0Z_9 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_9 ;
    wire bfn_14_5_0_;
    wire \U409_TICK.COUNTER60Z0Z_10 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_9 ;
    wire \U409_TICK.COUNTER60Z0Z_11 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_10 ;
    wire \U409_TICK.COUNTER60Z0Z_12 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_11 ;
    wire \U409_TICK.COUNTER60Z0Z_13 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_12 ;
    wire \U409_TICK.COUNTER60Z0Z_14 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_13 ;
    wire \U409_TICK.COUNTER60Z0Z_15 ;
    wire \U409_TICK.COUNTER60_RNO_0Z0Z_15 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_14 ;
    wire \U409_TICK.un3_COUNTER60_1_cry_15 ;
    wire \U409_TICK.COUNTER60Z0Z_16 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_6 ;
    wire \U409_TICK.COUNTER50Z0Z_3 ;
    wire \U409_TICK.COUNTER50Z0Z_0 ;
    wire \U409_TICK.COUNTER50Z0Z_12 ;
    wire \U409_TICK.TICK503_8_cascade_ ;
    wire \U409_TICK.COUNTER50Z0Z_10 ;
    wire \U409_TICK.TICK503_14_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_5 ;
    wire \U409_TICK.COUNTER50Z0Z_8 ;
    wire \U409_TICK.COUNTER50Z0Z_2 ;
    wire \U409_TICK.COUNTER50Z0Z_1 ;
    wire \U409_TICK.COUNTER50Z0Z_16 ;
    wire \U409_TICK.TICK503_11 ;
    wire TICK50_c;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_9 ;
    wire \U409_TICK.COUNTER50Z0Z_9 ;
    wire \U409_TICK.COUNTER50Z0Z_6 ;
    wire \U409_TICK.TICK503_9_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_13 ;
    wire \U409_TICK.COUNTER50Z0Z_13 ;
    wire \U409_TICK.COUNTER50Z0Z_7 ;
    wire \U409_TICK.COUNTER50Z0Z_4 ;
    wire \U409_TICK.TICK503_10_cascade_ ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_11 ;
    wire \U409_TICK.COUNTER50Z0Z_11 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_15 ;
    wire \U409_TICK.COUNTER50Z0Z_15 ;
    wire \U409_TICK.TICK503_14 ;
    wire \U409_TICK.TICK503_10 ;
    wire \U409_TICK.COUNTER50_RNO_0Z0Z_14 ;
    wire \U409_TICK.TICK503_9 ;
    wire \U409_TICK.COUNTER50Z0Z_14 ;
    wire CLK6_c_g;
    wire TACK_EN_i;
    wire N_475_i;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0001111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__5529),
            .RESETB(N__5253),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(CLK80_OUT));
    PRE_IO_GBUF CLK28_IN_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__7373),
            .GLOBALBUFFEROUTPUT(CLK28_IN_c_g));
    IO_PAD CLK28_IN_ibuf_gb_io_iopad (
            .OE(N__7375),
            .DIN(N__7374),
            .DOUT(N__7373),
            .PACKAGEPIN(CLK28_IN));
    defparam CLK28_IN_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK28_IN_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK28_IN_ibuf_gb_io_preio (
            .PADOEN(N__7375),
            .PADOUT(N__7374),
            .PADIN(N__7373),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF CLK6_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__7363),
            .GLOBALBUFFEROUTPUT(CLK6_c_g));
    IO_PAD CLK6_ibuf_gb_io_iopad (
            .OE(N__7365),
            .DIN(N__7364),
            .DOUT(N__7363),
            .PACKAGEPIN(CLK6));
    defparam CLK6_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK6_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK6_ibuf_gb_io_preio (
            .PADOEN(N__7365),
            .PADOUT(N__7364),
            .PADIN(N__7363),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_0_iopad (
            .OE(N__7354),
            .DIN(N__7353),
            .DOUT(N__7352),
            .PACKAGEPIN(TT[0]));
    defparam TT_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_0_preio (
            .PADOEN(N__7354),
            .PADOUT(N__7353),
            .PADIN(N__7352),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_6_iopad (
            .OE(N__7345),
            .DIN(N__7344),
            .DOUT(N__7343),
            .PACKAGEPIN(D[6]));
    defparam D_obuft_6_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_6_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_6_preio (
            .PADOEN(N__7345),
            .PADOUT(N__7344),
            .PADIN(N__7343),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RTC_ENn_obuf_iopad (
            .OE(N__7336),
            .DIN(N__7335),
            .DOUT(N__7334),
            .PACKAGEPIN(RTC_ENn));
    defparam RTC_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RTC_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RTC_ENn_obuf_preio (
            .PADOEN(N__7336),
            .PADOUT(N__7335),
            .PADIN(N__7334),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2934),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_24_iopad (
            .OE(N__7327),
            .DIN(N__7326),
            .DOUT(N__7325),
            .PACKAGEPIN(A[24]));
    defparam A_ibuf_24_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_24_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_24_preio (
            .PADOEN(N__7327),
            .PADOUT(N__7326),
            .PADIN(N__7325),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_24),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_5_iopad (
            .OE(N__7318),
            .DIN(N__7317),
            .DOUT(N__7316),
            .PACKAGEPIN(D[5]));
    defparam D_obuft_5_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_5_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_5_preio (
            .PADOEN(N__7318),
            .PADOUT(N__7317),
            .PADIN(N__7316),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_1_iopad (
            .OE(N__7309),
            .DIN(N__7308),
            .DOUT(N__7307),
            .PACKAGEPIN(TM[1]));
    defparam TM_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_1_preio (
            .PADOEN(N__7309),
            .PADOUT(N__7308),
            .PADIN(N__7307),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__7300),
            .DIN(N__7299),
            .DOUT(N__7298),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__7300),
            .PADOUT(N__7299),
            .PADIN(N__7298),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_CIA_obuf_iopad (
            .OE(N__7291),
            .DIN(N__7290),
            .DOUT(N__7289),
            .PACKAGEPIN(CLK_CIA));
    defparam CLK_CIA_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_CIA_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_CIA_obuf_preio (
            .PADOEN(N__7291),
            .PADOUT(N__7290),
            .PADIN(N__7289),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4920),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_21_iopad (
            .OE(N__7282),
            .DIN(N__7281),
            .DOUT(N__7280),
            .PACKAGEPIN(A[21]));
    defparam A_ibuf_21_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_21_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_21_preio (
            .PADOEN(N__7282),
            .PADOUT(N__7281),
            .PADIN(N__7280),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_21),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_obuf_iopad (
            .OE(N__7273),
            .DIN(N__7272),
            .DOUT(N__7271),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMSPACEn_obuf_preio (
            .PADOEN(N__7273),
            .PADOUT(N__7272),
            .PADIN(N__7271),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4044),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_iobuf_iopad (
            .OE(N__7264),
            .DIN(N__7263),
            .DOUT(N__7262),
            .PACKAGEPIN(TACKn));
    defparam TACKn_iobuf_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_iobuf_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_iobuf_preio (
            .PADOEN(N__7264),
            .PADOUT(N__7263),
            .PADIN(N__7262),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__6726),
            .DIN0(TACKn_in),
            .DOUT0(N__5319),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__7255),
            .DIN(N__7254),
            .DOUT(N__7253),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__7255),
            .PADOUT(N__7254),
            .PADIN(N__7253),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ROMENn_obuf_iopad (
            .OE(N__7246),
            .DIN(N__7245),
            .DOUT(N__7244),
            .PACKAGEPIN(ROMENn));
    defparam ROMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ROMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ROMENn_obuf_preio (
            .PADOEN(N__7246),
            .PADOUT(N__7245),
            .PADIN(N__7244),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5193),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_0_iopad (
            .OE(N__7237),
            .DIN(N__7236),
            .DOUT(N__7235),
            .PACKAGEPIN(D[0]));
    defparam D_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_0_preio (
            .PADOEN(N__7237),
            .PADOUT(N__7236),
            .PADIN(N__7235),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TT_ibuf_1_iopad (
            .OE(N__7228),
            .DIN(N__7227),
            .DOUT(N__7226),
            .PACKAGEPIN(TT[1]));
    defparam TT_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam TT_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO TT_ibuf_1_preio (
            .PADOEN(N__7228),
            .PADOUT(N__7227),
            .PADIN(N__7226),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TT_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__7219),
            .DIN(N__7218),
            .DOUT(N__7217),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__7219),
            .PADOUT(N__7218),
            .PADIN(N__7217),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUFENn_obuf_iopad (
            .OE(N__7210),
            .DIN(N__7209),
            .DOUT(N__7208),
            .PACKAGEPIN(BUFENn));
    defparam BUFENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BUFENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BUFENn_obuf_preio (
            .PADOEN(N__7210),
            .PADOUT(N__7209),
            .PADIN(N__7208),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3717),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORTSIZE_obuf_iopad (
            .OE(N__7201),
            .DIN(N__7200),
            .DOUT(N__7199),
            .PACKAGEPIN(PORTSIZE));
    defparam PORTSIZE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORTSIZE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORTSIZE_obuf_preio (
            .PADOEN(N__7201),
            .PADOUT(N__7200),
            .PADIN(N__7199),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4002),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_7_iopad (
            .OE(N__7192),
            .DIN(N__7191),
            .DOUT(N__7190),
            .PACKAGEPIN(D[7]));
    defparam D_obuft_7_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_7_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_7_preio (
            .PADOEN(N__7192),
            .PADOUT(N__7191),
            .PADIN(N__7190),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__7183),
            .DIN(N__7182),
            .DOUT(N__7181),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__7183),
            .PADOUT(N__7182),
            .PADIN(N__7181),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_29_iopad (
            .OE(N__7174),
            .DIN(N__7173),
            .DOUT(N__7172),
            .PACKAGEPIN(A[29]));
    defparam A_ibuf_29_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_29_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_29_preio (
            .PADOEN(N__7174),
            .PADOUT(N__7173),
            .PADIN(N__7172),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_29),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_22_iopad (
            .OE(N__7165),
            .DIN(N__7164),
            .DOUT(N__7163),
            .PACKAGEPIN(A[22]));
    defparam A_ibuf_22_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_22_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_22_preio (
            .PADOEN(N__7165),
            .PADOUT(N__7164),
            .PADIN(N__7163),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_22),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_27_iopad (
            .OE(N__7156),
            .DIN(N__7155),
            .DOUT(N__7154),
            .PACKAGEPIN(A[27]));
    defparam A_ibuf_27_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_27_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_27_preio (
            .PADOEN(N__7156),
            .PADOUT(N__7155),
            .PADIN(N__7154),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_27),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__7147),
            .DIN(N__7146),
            .DOUT(N__7145),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__7147),
            .PADOUT(N__7146),
            .PADIN(N__7145),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_2_iopad (
            .OE(N__7138),
            .DIN(N__7137),
            .DOUT(N__7136),
            .PACKAGEPIN(D[2]));
    defparam D_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_2_preio (
            .PADOEN(N__7138),
            .PADOUT(N__7137),
            .PADIN(N__7136),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__7129),
            .DIN(N__7128),
            .DOUT(N__7127),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__7129),
            .PADOUT(N__7128),
            .PADIN(N__7127),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TM_ibuf_0_iopad (
            .OE(N__7120),
            .DIN(N__7119),
            .DOUT(N__7118),
            .PACKAGEPIN(TM[0]));
    defparam TM_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam TM_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO TM_ibuf_0_preio (
            .PADOEN(N__7120),
            .PADOUT(N__7119),
            .PADIN(N__7118),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TM_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__7111),
            .DIN(N__7110),
            .DOUT(N__7109),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__7111),
            .PADOUT(N__7110),
            .PADIN(N__7109),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__7102),
            .DIN(N__7101),
            .DOUT(N__7100),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__7102),
            .PADOUT(N__7101),
            .PADIN(N__7100),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_25_iopad (
            .OE(N__7093),
            .DIN(N__7092),
            .DOUT(N__7091),
            .PACKAGEPIN(A[25]));
    defparam A_ibuf_25_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_25_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_25_preio (
            .PADOEN(N__7093),
            .PADOUT(N__7092),
            .PADIN(N__7091),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_25),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_1_iopad (
            .OE(N__7084),
            .DIN(N__7083),
            .DOUT(N__7082),
            .PACKAGEPIN(D[1]));
    defparam D_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_1_preio (
            .PADOEN(N__7084),
            .PADOUT(N__7083),
            .PADIN(N__7082),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS0n_obuf_iopad (
            .OE(N__7075),
            .DIN(N__7074),
            .DOUT(N__7073),
            .PACKAGEPIN(CIACS0n));
    defparam CIACS0n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS0n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS0n_obuf_preio (
            .PADOEN(N__7075),
            .PADOUT(N__7074),
            .PADIN(N__7073),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4311),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_4_iopad (
            .OE(N__7066),
            .DIN(N__7065),
            .DOUT(N__7064),
            .PACKAGEPIN(D[4]));
    defparam D_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_4_preio (
            .PADOEN(N__7066),
            .PADOUT(N__7065),
            .PADIN(N__7064),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK50_obuf_iopad (
            .OE(N__7057),
            .DIN(N__7056),
            .DOUT(N__7055),
            .PACKAGEPIN(TICK50));
    defparam TICK50_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK50_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK50_obuf_preio (
            .PADOEN(N__7057),
            .PADOUT(N__7056),
            .PADIN(N__7055),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6624),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__7048),
            .DIN(N__7047),
            .DOUT(N__7046),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__7048),
            .PADOUT(N__7047),
            .PADIN(N__7046),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_28_iopad (
            .OE(N__7039),
            .DIN(N__7038),
            .DOUT(N__7037),
            .PACKAGEPIN(A[28]));
    defparam A_ibuf_28_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_28_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_28_preio (
            .PADOEN(N__7039),
            .PADOUT(N__7038),
            .PADIN(N__7037),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_28),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_30_iopad (
            .OE(N__7030),
            .DIN(N__7029),
            .DOUT(N__7028),
            .PACKAGEPIN(A[30]));
    defparam A_ibuf_30_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_30_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_30_preio (
            .PADOEN(N__7030),
            .PADOUT(N__7029),
            .PADIN(N__7028),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_30),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD OVL_ibuf_iopad (
            .OE(N__7021),
            .DIN(N__7020),
            .DOUT(N__7019),
            .PACKAGEPIN(OVL));
    defparam OVL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam OVL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO OVL_ibuf_preio (
            .PADOEN(N__7021),
            .PADOUT(N__7020),
            .PADIN(N__7019),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(OVL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__7012),
            .DIN(N__7011),
            .DOUT(N__7010),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__7012),
            .PADOUT(N__7011),
            .PADIN(N__7010),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TICK60_obuf_iopad (
            .OE(N__7003),
            .DIN(N__7002),
            .DOUT(N__7001),
            .PACKAGEPIN(TICK60));
    defparam TICK60_obuf_preio.NEG_TRIGGER=1'b0;
    defparam TICK60_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO TICK60_obuf_preio (
            .PADOEN(N__7003),
            .PADOUT(N__7002),
            .PADIN(N__7001),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6072),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_26_iopad (
            .OE(N__6994),
            .DIN(N__6993),
            .DOUT(N__6992),
            .PACKAGEPIN(A[26]));
    defparam A_ibuf_26_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_26_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_26_preio (
            .PADOEN(N__6994),
            .PADOUT(N__6993),
            .PADIN(N__6992),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_26),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD D_obuft_3_iopad (
            .OE(N__6985),
            .DIN(N__6984),
            .DOUT(N__6983),
            .PACKAGEPIN(D[3]));
    defparam D_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam D_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO D_obuft_3_preio (
            .PADOEN(N__6985),
            .PADOUT(N__6984),
            .PADIN(N__6983),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_23_iopad (
            .OE(N__6976),
            .DIN(N__6975),
            .DOUT(N__6974),
            .PACKAGEPIN(A[23]));
    defparam A_ibuf_23_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_23_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_23_preio (
            .PADOEN(N__6976),
            .PADOUT(N__6975),
            .PADIN(N__6974),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_23),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_31_iopad (
            .OE(N__6967),
            .DIN(N__6966),
            .DOUT(N__6965),
            .PACKAGEPIN(A[31]));
    defparam A_ibuf_31_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_31_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_31_preio (
            .PADOEN(N__6967),
            .PADOUT(N__6966),
            .PADIN(N__6965),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_31),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CIACS1n_obuf_iopad (
            .OE(N__6958),
            .DIN(N__6957),
            .DOUT(N__6956),
            .PACKAGEPIN(CIACS1n));
    defparam CIACS1n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CIACS1n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CIACS1n_obuf_preio (
            .PADOEN(N__6958),
            .PADOUT(N__6957),
            .PADIN(N__6956),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4149),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_obuf_iopad (
            .OE(N__6949),
            .DIN(N__6948),
            .DOUT(N__6947),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGSPACEn_obuf_preio (
            .PADOEN(N__6949),
            .PADOUT(N__6948),
            .PADIN(N__6947),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3489),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1603 (
            .O(N__6930),
            .I(N__6927));
    LocalMux I__1602 (
            .O(N__6927),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ));
    InMux I__1601 (
            .O(N__6924),
            .I(N__6920));
    InMux I__1600 (
            .O(N__6923),
            .I(N__6917));
    LocalMux I__1599 (
            .O(N__6920),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    LocalMux I__1598 (
            .O(N__6917),
            .I(\U409_TICK.COUNTER50Z0Z_15 ));
    InMux I__1597 (
            .O(N__6912),
            .I(N__6894));
    InMux I__1596 (
            .O(N__6911),
            .I(N__6894));
    InMux I__1595 (
            .O(N__6910),
            .I(N__6894));
    InMux I__1594 (
            .O(N__6909),
            .I(N__6894));
    InMux I__1593 (
            .O(N__6908),
            .I(N__6894));
    InMux I__1592 (
            .O(N__6907),
            .I(N__6887));
    InMux I__1591 (
            .O(N__6906),
            .I(N__6887));
    InMux I__1590 (
            .O(N__6905),
            .I(N__6887));
    LocalMux I__1589 (
            .O(N__6894),
            .I(\U409_TICK.TICK503_14 ));
    LocalMux I__1588 (
            .O(N__6887),
            .I(\U409_TICK.TICK503_14 ));
    InMux I__1587 (
            .O(N__6882),
            .I(N__6866));
    InMux I__1586 (
            .O(N__6881),
            .I(N__6866));
    InMux I__1585 (
            .O(N__6880),
            .I(N__6866));
    InMux I__1584 (
            .O(N__6879),
            .I(N__6866));
    InMux I__1583 (
            .O(N__6878),
            .I(N__6857));
    InMux I__1582 (
            .O(N__6877),
            .I(N__6857));
    InMux I__1581 (
            .O(N__6876),
            .I(N__6857));
    InMux I__1580 (
            .O(N__6875),
            .I(N__6857));
    LocalMux I__1579 (
            .O(N__6866),
            .I(\U409_TICK.TICK503_10 ));
    LocalMux I__1578 (
            .O(N__6857),
            .I(\U409_TICK.TICK503_10 ));
    CascadeMux I__1577 (
            .O(N__6852),
            .I(N__6849));
    InMux I__1576 (
            .O(N__6849),
            .I(N__6846));
    LocalMux I__1575 (
            .O(N__6846),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ));
    CascadeMux I__1574 (
            .O(N__6843),
            .I(N__6840));
    InMux I__1573 (
            .O(N__6840),
            .I(N__6830));
    InMux I__1572 (
            .O(N__6839),
            .I(N__6830));
    CascadeMux I__1571 (
            .O(N__6838),
            .I(N__6827));
    CascadeMux I__1570 (
            .O(N__6837),
            .I(N__6824));
    CascadeMux I__1569 (
            .O(N__6836),
            .I(N__6821));
    CascadeMux I__1568 (
            .O(N__6835),
            .I(N__6816));
    LocalMux I__1567 (
            .O(N__6830),
            .I(N__6813));
    InMux I__1566 (
            .O(N__6827),
            .I(N__6808));
    InMux I__1565 (
            .O(N__6824),
            .I(N__6808));
    InMux I__1564 (
            .O(N__6821),
            .I(N__6799));
    InMux I__1563 (
            .O(N__6820),
            .I(N__6799));
    InMux I__1562 (
            .O(N__6819),
            .I(N__6799));
    InMux I__1561 (
            .O(N__6816),
            .I(N__6799));
    Odrv4 I__1560 (
            .O(N__6813),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1559 (
            .O(N__6808),
            .I(\U409_TICK.TICK503_9 ));
    LocalMux I__1558 (
            .O(N__6799),
            .I(\U409_TICK.TICK503_9 ));
    CascadeMux I__1557 (
            .O(N__6792),
            .I(N__6789));
    InMux I__1556 (
            .O(N__6789),
            .I(N__6785));
    InMux I__1555 (
            .O(N__6788),
            .I(N__6782));
    LocalMux I__1554 (
            .O(N__6785),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    LocalMux I__1553 (
            .O(N__6782),
            .I(\U409_TICK.COUNTER50Z0Z_14 ));
    ClkMux I__1552 (
            .O(N__6777),
            .I(N__6750));
    ClkMux I__1551 (
            .O(N__6776),
            .I(N__6750));
    ClkMux I__1550 (
            .O(N__6775),
            .I(N__6750));
    ClkMux I__1549 (
            .O(N__6774),
            .I(N__6750));
    ClkMux I__1548 (
            .O(N__6773),
            .I(N__6750));
    ClkMux I__1547 (
            .O(N__6772),
            .I(N__6750));
    ClkMux I__1546 (
            .O(N__6771),
            .I(N__6750));
    ClkMux I__1545 (
            .O(N__6770),
            .I(N__6750));
    ClkMux I__1544 (
            .O(N__6769),
            .I(N__6750));
    GlobalMux I__1543 (
            .O(N__6750),
            .I(N__6747));
    gio2CtrlBuf I__1542 (
            .O(N__6747),
            .I(CLK6_c_g));
    InMux I__1541 (
            .O(N__6744),
            .I(N__6741));
    LocalMux I__1540 (
            .O(N__6741),
            .I(N__6738));
    Span4Mux_v I__1539 (
            .O(N__6738),
            .I(N__6735));
    Span4Mux_h I__1538 (
            .O(N__6735),
            .I(N__6732));
    Span4Mux_h I__1537 (
            .O(N__6732),
            .I(N__6729));
    Odrv4 I__1536 (
            .O(N__6729),
            .I(TACK_EN_i));
    IoInMux I__1535 (
            .O(N__6726),
            .I(N__6723));
    LocalMux I__1534 (
            .O(N__6723),
            .I(N__6720));
    Span4Mux_s1_v I__1533 (
            .O(N__6720),
            .I(N__6717));
    Span4Mux_h I__1532 (
            .O(N__6717),
            .I(N__6714));
    Span4Mux_v I__1531 (
            .O(N__6714),
            .I(N__6711));
    Odrv4 I__1530 (
            .O(N__6711),
            .I(N_475_i));
    CascadeMux I__1529 (
            .O(N__6708),
            .I(\U409_TICK.TICK503_14_cascade_ ));
    InMux I__1528 (
            .O(N__6705),
            .I(N__6702));
    LocalMux I__1527 (
            .O(N__6702),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ));
    InMux I__1526 (
            .O(N__6699),
            .I(N__6695));
    InMux I__1525 (
            .O(N__6698),
            .I(N__6692));
    LocalMux I__1524 (
            .O(N__6695),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    LocalMux I__1523 (
            .O(N__6692),
            .I(\U409_TICK.COUNTER50Z0Z_5 ));
    InMux I__1522 (
            .O(N__6687),
            .I(N__6683));
    InMux I__1521 (
            .O(N__6686),
            .I(N__6680));
    LocalMux I__1520 (
            .O(N__6683),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    LocalMux I__1519 (
            .O(N__6680),
            .I(\U409_TICK.COUNTER50Z0Z_8 ));
    InMux I__1518 (
            .O(N__6675),
            .I(N__6671));
    InMux I__1517 (
            .O(N__6674),
            .I(N__6668));
    LocalMux I__1516 (
            .O(N__6671),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    LocalMux I__1515 (
            .O(N__6668),
            .I(\U409_TICK.COUNTER50Z0Z_2 ));
    CascadeMux I__1514 (
            .O(N__6663),
            .I(N__6659));
    CascadeMux I__1513 (
            .O(N__6662),
            .I(N__6656));
    InMux I__1512 (
            .O(N__6659),
            .I(N__6650));
    InMux I__1511 (
            .O(N__6656),
            .I(N__6650));
    InMux I__1510 (
            .O(N__6655),
            .I(N__6647));
    LocalMux I__1509 (
            .O(N__6650),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    LocalMux I__1508 (
            .O(N__6647),
            .I(\U409_TICK.COUNTER50Z0Z_1 ));
    InMux I__1507 (
            .O(N__6642),
            .I(N__6638));
    InMux I__1506 (
            .O(N__6641),
            .I(N__6635));
    LocalMux I__1505 (
            .O(N__6638),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    LocalMux I__1504 (
            .O(N__6635),
            .I(\U409_TICK.COUNTER50Z0Z_16 ));
    InMux I__1503 (
            .O(N__6630),
            .I(N__6627));
    LocalMux I__1502 (
            .O(N__6627),
            .I(\U409_TICK.TICK503_11 ));
    IoInMux I__1501 (
            .O(N__6624),
            .I(N__6621));
    LocalMux I__1500 (
            .O(N__6621),
            .I(N__6618));
    Span4Mux_s3_v I__1499 (
            .O(N__6618),
            .I(N__6615));
    Span4Mux_h I__1498 (
            .O(N__6615),
            .I(N__6611));
    InMux I__1497 (
            .O(N__6614),
            .I(N__6608));
    Odrv4 I__1496 (
            .O(N__6611),
            .I(TICK50_c));
    LocalMux I__1495 (
            .O(N__6608),
            .I(TICK50_c));
    InMux I__1494 (
            .O(N__6603),
            .I(N__6600));
    LocalMux I__1493 (
            .O(N__6600),
            .I(N__6597));
    Odrv4 I__1492 (
            .O(N__6597),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ));
    InMux I__1491 (
            .O(N__6594),
            .I(N__6590));
    InMux I__1490 (
            .O(N__6593),
            .I(N__6587));
    LocalMux I__1489 (
            .O(N__6590),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    LocalMux I__1488 (
            .O(N__6587),
            .I(\U409_TICK.COUNTER50Z0Z_9 ));
    CascadeMux I__1487 (
            .O(N__6582),
            .I(N__6579));
    InMux I__1486 (
            .O(N__6579),
            .I(N__6575));
    InMux I__1485 (
            .O(N__6578),
            .I(N__6572));
    LocalMux I__1484 (
            .O(N__6575),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    LocalMux I__1483 (
            .O(N__6572),
            .I(\U409_TICK.COUNTER50Z0Z_6 ));
    CascadeMux I__1482 (
            .O(N__6567),
            .I(\U409_TICK.TICK503_9_cascade_ ));
    InMux I__1481 (
            .O(N__6564),
            .I(N__6561));
    LocalMux I__1480 (
            .O(N__6561),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ));
    InMux I__1479 (
            .O(N__6558),
            .I(N__6554));
    InMux I__1478 (
            .O(N__6557),
            .I(N__6551));
    LocalMux I__1477 (
            .O(N__6554),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    LocalMux I__1476 (
            .O(N__6551),
            .I(\U409_TICK.COUNTER50Z0Z_13 ));
    InMux I__1475 (
            .O(N__6546),
            .I(N__6542));
    InMux I__1474 (
            .O(N__6545),
            .I(N__6539));
    LocalMux I__1473 (
            .O(N__6542),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    LocalMux I__1472 (
            .O(N__6539),
            .I(\U409_TICK.COUNTER50Z0Z_7 ));
    InMux I__1471 (
            .O(N__6534),
            .I(N__6530));
    InMux I__1470 (
            .O(N__6533),
            .I(N__6527));
    LocalMux I__1469 (
            .O(N__6530),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    LocalMux I__1468 (
            .O(N__6527),
            .I(\U409_TICK.COUNTER50Z0Z_4 ));
    CascadeMux I__1467 (
            .O(N__6522),
            .I(\U409_TICK.TICK503_10_cascade_ ));
    InMux I__1466 (
            .O(N__6519),
            .I(N__6516));
    LocalMux I__1465 (
            .O(N__6516),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ));
    InMux I__1464 (
            .O(N__6513),
            .I(N__6509));
    InMux I__1463 (
            .O(N__6512),
            .I(N__6506));
    LocalMux I__1462 (
            .O(N__6509),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    LocalMux I__1461 (
            .O(N__6506),
            .I(\U409_TICK.COUNTER50Z0Z_11 ));
    InMux I__1460 (
            .O(N__6501),
            .I(N__6497));
    InMux I__1459 (
            .O(N__6500),
            .I(N__6494));
    LocalMux I__1458 (
            .O(N__6497),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    LocalMux I__1457 (
            .O(N__6494),
            .I(\U409_TICK.COUNTER60Z0Z_13 ));
    InMux I__1456 (
            .O(N__6489),
            .I(\U409_TICK.un3_COUNTER60_1_cry_12 ));
    InMux I__1455 (
            .O(N__6486),
            .I(N__6482));
    InMux I__1454 (
            .O(N__6485),
            .I(N__6479));
    LocalMux I__1453 (
            .O(N__6482),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    LocalMux I__1452 (
            .O(N__6479),
            .I(\U409_TICK.COUNTER60Z0Z_14 ));
    InMux I__1451 (
            .O(N__6474),
            .I(N__6471));
    LocalMux I__1450 (
            .O(N__6471),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ));
    InMux I__1449 (
            .O(N__6468),
            .I(\U409_TICK.un3_COUNTER60_1_cry_13 ));
    InMux I__1448 (
            .O(N__6465),
            .I(N__6461));
    InMux I__1447 (
            .O(N__6464),
            .I(N__6458));
    LocalMux I__1446 (
            .O(N__6461),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    LocalMux I__1445 (
            .O(N__6458),
            .I(\U409_TICK.COUNTER60Z0Z_15 ));
    InMux I__1444 (
            .O(N__6453),
            .I(N__6450));
    LocalMux I__1443 (
            .O(N__6450),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ));
    InMux I__1442 (
            .O(N__6447),
            .I(\U409_TICK.un3_COUNTER60_1_cry_14 ));
    InMux I__1441 (
            .O(N__6444),
            .I(\U409_TICK.un3_COUNTER60_1_cry_15 ));
    InMux I__1440 (
            .O(N__6441),
            .I(N__6437));
    InMux I__1439 (
            .O(N__6440),
            .I(N__6434));
    LocalMux I__1438 (
            .O(N__6437),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    LocalMux I__1437 (
            .O(N__6434),
            .I(\U409_TICK.COUNTER60Z0Z_16 ));
    InMux I__1436 (
            .O(N__6429),
            .I(N__6426));
    LocalMux I__1435 (
            .O(N__6426),
            .I(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ));
    InMux I__1434 (
            .O(N__6423),
            .I(N__6419));
    InMux I__1433 (
            .O(N__6422),
            .I(N__6416));
    LocalMux I__1432 (
            .O(N__6419),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    LocalMux I__1431 (
            .O(N__6416),
            .I(\U409_TICK.COUNTER50Z0Z_3 ));
    CascadeMux I__1430 (
            .O(N__6411),
            .I(N__6405));
    InMux I__1429 (
            .O(N__6410),
            .I(N__6398));
    InMux I__1428 (
            .O(N__6409),
            .I(N__6398));
    InMux I__1427 (
            .O(N__6408),
            .I(N__6398));
    InMux I__1426 (
            .O(N__6405),
            .I(N__6395));
    LocalMux I__1425 (
            .O(N__6398),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    LocalMux I__1424 (
            .O(N__6395),
            .I(\U409_TICK.COUNTER50Z0Z_0 ));
    InMux I__1423 (
            .O(N__6390),
            .I(N__6386));
    InMux I__1422 (
            .O(N__6389),
            .I(N__6383));
    LocalMux I__1421 (
            .O(N__6386),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    LocalMux I__1420 (
            .O(N__6383),
            .I(\U409_TICK.COUNTER50Z0Z_12 ));
    CascadeMux I__1419 (
            .O(N__6378),
            .I(\U409_TICK.TICK503_8_cascade_ ));
    InMux I__1418 (
            .O(N__6375),
            .I(N__6371));
    InMux I__1417 (
            .O(N__6374),
            .I(N__6368));
    LocalMux I__1416 (
            .O(N__6371),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    LocalMux I__1415 (
            .O(N__6368),
            .I(\U409_TICK.COUNTER50Z0Z_10 ));
    InMux I__1414 (
            .O(N__6363),
            .I(N__6359));
    InMux I__1413 (
            .O(N__6362),
            .I(N__6356));
    LocalMux I__1412 (
            .O(N__6359),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    LocalMux I__1411 (
            .O(N__6356),
            .I(\U409_TICK.COUNTER60Z0Z_5 ));
    InMux I__1410 (
            .O(N__6351),
            .I(\U409_TICK.un3_COUNTER60_1_cry_4 ));
    InMux I__1409 (
            .O(N__6348),
            .I(N__6344));
    InMux I__1408 (
            .O(N__6347),
            .I(N__6341));
    LocalMux I__1407 (
            .O(N__6344),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    LocalMux I__1406 (
            .O(N__6341),
            .I(\U409_TICK.COUNTER60Z0Z_6 ));
    InMux I__1405 (
            .O(N__6336),
            .I(N__6333));
    LocalMux I__1404 (
            .O(N__6333),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ));
    InMux I__1403 (
            .O(N__6330),
            .I(\U409_TICK.un3_COUNTER60_1_cry_5 ));
    CascadeMux I__1402 (
            .O(N__6327),
            .I(N__6324));
    InMux I__1401 (
            .O(N__6324),
            .I(N__6320));
    InMux I__1400 (
            .O(N__6323),
            .I(N__6317));
    LocalMux I__1399 (
            .O(N__6320),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    LocalMux I__1398 (
            .O(N__6317),
            .I(\U409_TICK.COUNTER60Z0Z_7 ));
    InMux I__1397 (
            .O(N__6312),
            .I(\U409_TICK.un3_COUNTER60_1_cry_6 ));
    CascadeMux I__1396 (
            .O(N__6309),
            .I(N__6306));
    InMux I__1395 (
            .O(N__6306),
            .I(N__6302));
    InMux I__1394 (
            .O(N__6305),
            .I(N__6299));
    LocalMux I__1393 (
            .O(N__6302),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    LocalMux I__1392 (
            .O(N__6299),
            .I(\U409_TICK.COUNTER60Z0Z_8 ));
    InMux I__1391 (
            .O(N__6294),
            .I(N__6291));
    LocalMux I__1390 (
            .O(N__6291),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ));
    InMux I__1389 (
            .O(N__6288),
            .I(\U409_TICK.un3_COUNTER60_1_cry_7 ));
    InMux I__1388 (
            .O(N__6285),
            .I(N__6281));
    InMux I__1387 (
            .O(N__6284),
            .I(N__6278));
    LocalMux I__1386 (
            .O(N__6281),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    LocalMux I__1385 (
            .O(N__6278),
            .I(\U409_TICK.COUNTER60Z0Z_9 ));
    CascadeMux I__1384 (
            .O(N__6273),
            .I(N__6270));
    InMux I__1383 (
            .O(N__6270),
            .I(N__6267));
    LocalMux I__1382 (
            .O(N__6267),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ));
    InMux I__1381 (
            .O(N__6264),
            .I(bfn_14_5_0_));
    InMux I__1380 (
            .O(N__6261),
            .I(N__6257));
    InMux I__1379 (
            .O(N__6260),
            .I(N__6254));
    LocalMux I__1378 (
            .O(N__6257),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    LocalMux I__1377 (
            .O(N__6254),
            .I(\U409_TICK.COUNTER60Z0Z_10 ));
    InMux I__1376 (
            .O(N__6249),
            .I(\U409_TICK.un3_COUNTER60_1_cry_9 ));
    InMux I__1375 (
            .O(N__6246),
            .I(N__6242));
    InMux I__1374 (
            .O(N__6245),
            .I(N__6239));
    LocalMux I__1373 (
            .O(N__6242),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    LocalMux I__1372 (
            .O(N__6239),
            .I(\U409_TICK.COUNTER60Z0Z_11 ));
    InMux I__1371 (
            .O(N__6234),
            .I(\U409_TICK.un3_COUNTER60_1_cry_10 ));
    InMux I__1370 (
            .O(N__6231),
            .I(N__6227));
    InMux I__1369 (
            .O(N__6230),
            .I(N__6224));
    LocalMux I__1368 (
            .O(N__6227),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    LocalMux I__1367 (
            .O(N__6224),
            .I(\U409_TICK.COUNTER60Z0Z_12 ));
    InMux I__1366 (
            .O(N__6219),
            .I(\U409_TICK.un3_COUNTER60_1_cry_11 ));
    InMux I__1365 (
            .O(N__6216),
            .I(\U409_TICK.un2_COUNTER50_1_cry_11 ));
    InMux I__1364 (
            .O(N__6213),
            .I(\U409_TICK.un2_COUNTER50_1_cry_12 ));
    InMux I__1363 (
            .O(N__6210),
            .I(\U409_TICK.un2_COUNTER50_1_cry_13 ));
    InMux I__1362 (
            .O(N__6207),
            .I(\U409_TICK.un2_COUNTER50_1_cry_14 ));
    InMux I__1361 (
            .O(N__6204),
            .I(\U409_TICK.un2_COUNTER50_1_cry_15 ));
    CascadeMux I__1360 (
            .O(N__6201),
            .I(N__6197));
    CascadeMux I__1359 (
            .O(N__6200),
            .I(N__6194));
    InMux I__1358 (
            .O(N__6197),
            .I(N__6190));
    InMux I__1357 (
            .O(N__6194),
            .I(N__6187));
    InMux I__1356 (
            .O(N__6193),
            .I(N__6184));
    LocalMux I__1355 (
            .O(N__6190),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__1354 (
            .O(N__6187),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    LocalMux I__1353 (
            .O(N__6184),
            .I(\U409_TICK.COUNTER60Z0Z_1 ));
    CascadeMux I__1352 (
            .O(N__6177),
            .I(N__6171));
    InMux I__1351 (
            .O(N__6176),
            .I(N__6164));
    InMux I__1350 (
            .O(N__6175),
            .I(N__6164));
    InMux I__1349 (
            .O(N__6174),
            .I(N__6164));
    InMux I__1348 (
            .O(N__6171),
            .I(N__6161));
    LocalMux I__1347 (
            .O(N__6164),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    LocalMux I__1346 (
            .O(N__6161),
            .I(\U409_TICK.COUNTER60Z0Z_0 ));
    InMux I__1345 (
            .O(N__6156),
            .I(N__6152));
    InMux I__1344 (
            .O(N__6155),
            .I(N__6149));
    LocalMux I__1343 (
            .O(N__6152),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    LocalMux I__1342 (
            .O(N__6149),
            .I(\U409_TICK.COUNTER60Z0Z_2 ));
    InMux I__1341 (
            .O(N__6144),
            .I(\U409_TICK.un3_COUNTER60_1_cry_1 ));
    InMux I__1340 (
            .O(N__6141),
            .I(N__6137));
    InMux I__1339 (
            .O(N__6140),
            .I(N__6134));
    LocalMux I__1338 (
            .O(N__6137),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    LocalMux I__1337 (
            .O(N__6134),
            .I(\U409_TICK.COUNTER60Z0Z_3 ));
    InMux I__1336 (
            .O(N__6129),
            .I(\U409_TICK.un3_COUNTER60_1_cry_2 ));
    InMux I__1335 (
            .O(N__6126),
            .I(N__6122));
    InMux I__1334 (
            .O(N__6125),
            .I(N__6119));
    LocalMux I__1333 (
            .O(N__6122),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    LocalMux I__1332 (
            .O(N__6119),
            .I(\U409_TICK.COUNTER60Z0Z_4 ));
    CascadeMux I__1331 (
            .O(N__6114),
            .I(N__6111));
    InMux I__1330 (
            .O(N__6111),
            .I(N__6108));
    LocalMux I__1329 (
            .O(N__6108),
            .I(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ));
    InMux I__1328 (
            .O(N__6105),
            .I(\U409_TICK.un3_COUNTER60_1_cry_3 ));
    InMux I__1327 (
            .O(N__6102),
            .I(\U409_TICK.un2_COUNTER50_1_cry_2 ));
    InMux I__1326 (
            .O(N__6099),
            .I(\U409_TICK.un2_COUNTER50_1_cry_3 ));
    InMux I__1325 (
            .O(N__6096),
            .I(\U409_TICK.un2_COUNTER50_1_cry_4 ));
    InMux I__1324 (
            .O(N__6093),
            .I(\U409_TICK.un2_COUNTER50_1_cry_5 ));
    InMux I__1323 (
            .O(N__6090),
            .I(\U409_TICK.un2_COUNTER50_1_cry_6 ));
    InMux I__1322 (
            .O(N__6087),
            .I(\U409_TICK.un2_COUNTER50_1_cry_7 ));
    InMux I__1321 (
            .O(N__6084),
            .I(bfn_14_2_0_));
    InMux I__1320 (
            .O(N__6081),
            .I(\U409_TICK.un2_COUNTER50_1_cry_9 ));
    InMux I__1319 (
            .O(N__6078),
            .I(\U409_TICK.un2_COUNTER50_1_cry_10 ));
    CascadeMux I__1318 (
            .O(N__6075),
            .I(\U409_TICK.TICK603_9_cascade_ ));
    IoInMux I__1317 (
            .O(N__6072),
            .I(N__6069));
    LocalMux I__1316 (
            .O(N__6069),
            .I(N__6066));
    Span4Mux_s3_v I__1315 (
            .O(N__6066),
            .I(N__6063));
    Span4Mux_v I__1314 (
            .O(N__6063),
            .I(N__6060));
    Span4Mux_h I__1313 (
            .O(N__6060),
            .I(N__6056));
    InMux I__1312 (
            .O(N__6059),
            .I(N__6053));
    Odrv4 I__1311 (
            .O(N__6056),
            .I(TICK60_c));
    LocalMux I__1310 (
            .O(N__6053),
            .I(TICK60_c));
    CascadeMux I__1309 (
            .O(N__6048),
            .I(\U409_TICK.TICK603_10_cascade_ ));
    InMux I__1308 (
            .O(N__6045),
            .I(N__6042));
    LocalMux I__1307 (
            .O(N__6042),
            .I(\U409_TICK.TICK603_11 ));
    InMux I__1306 (
            .O(N__6039),
            .I(N__6030));
    InMux I__1305 (
            .O(N__6038),
            .I(N__6023));
    InMux I__1304 (
            .O(N__6037),
            .I(N__6023));
    InMux I__1303 (
            .O(N__6036),
            .I(N__6023));
    InMux I__1302 (
            .O(N__6035),
            .I(N__6016));
    InMux I__1301 (
            .O(N__6034),
            .I(N__6016));
    InMux I__1300 (
            .O(N__6033),
            .I(N__6016));
    LocalMux I__1299 (
            .O(N__6030),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1298 (
            .O(N__6023),
            .I(\U409_TICK.TICK603_14 ));
    LocalMux I__1297 (
            .O(N__6016),
            .I(\U409_TICK.TICK603_14 ));
    CascadeMux I__1296 (
            .O(N__6009),
            .I(N__6002));
    InMux I__1295 (
            .O(N__6008),
            .I(N__5997));
    InMux I__1294 (
            .O(N__6007),
            .I(N__5990));
    InMux I__1293 (
            .O(N__6006),
            .I(N__5990));
    InMux I__1292 (
            .O(N__6005),
            .I(N__5990));
    InMux I__1291 (
            .O(N__6002),
            .I(N__5983));
    InMux I__1290 (
            .O(N__6001),
            .I(N__5983));
    InMux I__1289 (
            .O(N__6000),
            .I(N__5983));
    LocalMux I__1288 (
            .O(N__5997),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__1287 (
            .O(N__5990),
            .I(\U409_TICK.TICK603_9 ));
    LocalMux I__1286 (
            .O(N__5983),
            .I(\U409_TICK.TICK603_9 ));
    CascadeMux I__1285 (
            .O(N__5976),
            .I(N__5972));
    CascadeMux I__1284 (
            .O(N__5975),
            .I(N__5969));
    InMux I__1283 (
            .O(N__5972),
            .I(N__5961));
    InMux I__1282 (
            .O(N__5969),
            .I(N__5956));
    InMux I__1281 (
            .O(N__5968),
            .I(N__5956));
    InMux I__1280 (
            .O(N__5967),
            .I(N__5947));
    InMux I__1279 (
            .O(N__5966),
            .I(N__5947));
    InMux I__1278 (
            .O(N__5965),
            .I(N__5947));
    InMux I__1277 (
            .O(N__5964),
            .I(N__5947));
    LocalMux I__1276 (
            .O(N__5961),
            .I(N__5944));
    LocalMux I__1275 (
            .O(N__5956),
            .I(\U409_TICK.TICK603_10 ));
    LocalMux I__1274 (
            .O(N__5947),
            .I(\U409_TICK.TICK603_10 ));
    Odrv4 I__1273 (
            .O(N__5944),
            .I(\U409_TICK.TICK603_10 ));
    InMux I__1272 (
            .O(N__5937),
            .I(\U409_TICK.un2_COUNTER50_1_cry_1 ));
    CascadeMux I__1271 (
            .O(N__5934),
            .I(N__5927));
    CascadeMux I__1270 (
            .O(N__5933),
            .I(N__5924));
    InMux I__1269 (
            .O(N__5932),
            .I(N__5921));
    InMux I__1268 (
            .O(N__5931),
            .I(N__5912));
    InMux I__1267 (
            .O(N__5930),
            .I(N__5912));
    InMux I__1266 (
            .O(N__5927),
            .I(N__5912));
    InMux I__1265 (
            .O(N__5924),
            .I(N__5912));
    LocalMux I__1264 (
            .O(N__5921),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    LocalMux I__1263 (
            .O(N__5912),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ));
    InMux I__1262 (
            .O(N__5907),
            .I(N__5900));
    InMux I__1261 (
            .O(N__5906),
            .I(N__5891));
    InMux I__1260 (
            .O(N__5905),
            .I(N__5891));
    InMux I__1259 (
            .O(N__5904),
            .I(N__5891));
    InMux I__1258 (
            .O(N__5903),
            .I(N__5891));
    LocalMux I__1257 (
            .O(N__5900),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    LocalMux I__1256 (
            .O(N__5891),
            .I(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ));
    InMux I__1255 (
            .O(N__5886),
            .I(N__5882));
    CascadeMux I__1254 (
            .O(N__5885),
            .I(N__5879));
    LocalMux I__1253 (
            .O(N__5882),
            .I(N__5874));
    InMux I__1252 (
            .O(N__5879),
            .I(N__5871));
    InMux I__1251 (
            .O(N__5878),
            .I(N__5867));
    CascadeMux I__1250 (
            .O(N__5877),
            .I(N__5864));
    Span4Mux_v I__1249 (
            .O(N__5874),
            .I(N__5861));
    LocalMux I__1248 (
            .O(N__5871),
            .I(N__5858));
    InMux I__1247 (
            .O(N__5870),
            .I(N__5855));
    LocalMux I__1246 (
            .O(N__5867),
            .I(N__5852));
    InMux I__1245 (
            .O(N__5864),
            .I(N__5849));
    Span4Mux_h I__1244 (
            .O(N__5861),
            .I(N__5839));
    Span4Mux_v I__1243 (
            .O(N__5858),
            .I(N__5839));
    LocalMux I__1242 (
            .O(N__5855),
            .I(N__5839));
    Span4Mux_h I__1241 (
            .O(N__5852),
            .I(N__5832));
    LocalMux I__1240 (
            .O(N__5849),
            .I(N__5832));
    CascadeMux I__1239 (
            .O(N__5848),
            .I(N__5829));
    CascadeMux I__1238 (
            .O(N__5847),
            .I(N__5823));
    CascadeMux I__1237 (
            .O(N__5846),
            .I(N__5819));
    Span4Mux_v I__1236 (
            .O(N__5839),
            .I(N__5816));
    InMux I__1235 (
            .O(N__5838),
            .I(N__5813));
    InMux I__1234 (
            .O(N__5837),
            .I(N__5810));
    Span4Mux_h I__1233 (
            .O(N__5832),
            .I(N__5807));
    InMux I__1232 (
            .O(N__5829),
            .I(N__5804));
    InMux I__1231 (
            .O(N__5828),
            .I(N__5801));
    InMux I__1230 (
            .O(N__5827),
            .I(N__5794));
    InMux I__1229 (
            .O(N__5826),
            .I(N__5794));
    InMux I__1228 (
            .O(N__5823),
            .I(N__5794));
    InMux I__1227 (
            .O(N__5822),
            .I(N__5789));
    InMux I__1226 (
            .O(N__5819),
            .I(N__5789));
    Sp12to4 I__1225 (
            .O(N__5816),
            .I(N__5785));
    LocalMux I__1224 (
            .O(N__5813),
            .I(N__5780));
    LocalMux I__1223 (
            .O(N__5810),
            .I(N__5780));
    Sp12to4 I__1222 (
            .O(N__5807),
            .I(N__5771));
    LocalMux I__1221 (
            .O(N__5804),
            .I(N__5771));
    LocalMux I__1220 (
            .O(N__5801),
            .I(N__5771));
    LocalMux I__1219 (
            .O(N__5794),
            .I(N__5771));
    LocalMux I__1218 (
            .O(N__5789),
            .I(N__5768));
    InMux I__1217 (
            .O(N__5788),
            .I(N__5765));
    Span12Mux_h I__1216 (
            .O(N__5785),
            .I(N__5762));
    Span4Mux_v I__1215 (
            .O(N__5780),
            .I(N__5759));
    Span12Mux_v I__1214 (
            .O(N__5771),
            .I(N__5752));
    Sp12to4 I__1213 (
            .O(N__5768),
            .I(N__5752));
    LocalMux I__1212 (
            .O(N__5765),
            .I(N__5752));
    Span12Mux_v I__1211 (
            .O(N__5762),
            .I(N__5749));
    Sp12to4 I__1210 (
            .O(N__5759),
            .I(N__5746));
    Span12Mux_v I__1209 (
            .O(N__5752),
            .I(N__5743));
    Span12Mux_h I__1208 (
            .O(N__5749),
            .I(N__5740));
    Span12Mux_h I__1207 (
            .O(N__5746),
            .I(N__5737));
    Span12Mux_h I__1206 (
            .O(N__5743),
            .I(N__5734));
    Odrv12 I__1205 (
            .O(N__5740),
            .I(RESETn_c));
    Odrv12 I__1204 (
            .O(N__5737),
            .I(RESETn_c));
    Odrv12 I__1203 (
            .O(N__5734),
            .I(RESETn_c));
    InMux I__1202 (
            .O(N__5727),
            .I(N__5724));
    LocalMux I__1201 (
            .O(N__5724),
            .I(N__5718));
    InMux I__1200 (
            .O(N__5723),
            .I(N__5711));
    InMux I__1199 (
            .O(N__5722),
            .I(N__5711));
    InMux I__1198 (
            .O(N__5721),
            .I(N__5711));
    Odrv4 I__1197 (
            .O(N__5718),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    LocalMux I__1196 (
            .O(N__5711),
            .I(\U409_TRANSFER_ACK.TACK_COUNTER6 ));
    CEMux I__1195 (
            .O(N__5706),
            .I(N__5703));
    LocalMux I__1194 (
            .O(N__5703),
            .I(N__5700));
    Odrv4 I__1193 (
            .O(N__5700),
            .I(\U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en ));
    CascadeMux I__1192 (
            .O(N__5697),
            .I(\U409_TICK.TICK603_8_cascade_ ));
    CascadeMux I__1191 (
            .O(N__5694),
            .I(\U409_TICK.TICK603_14_cascade_ ));
    CascadeMux I__1190 (
            .O(N__5691),
            .I(N__5686));
    CascadeMux I__1189 (
            .O(N__5690),
            .I(N__5683));
    CascadeMux I__1188 (
            .O(N__5689),
            .I(N__5678));
    InMux I__1187 (
            .O(N__5686),
            .I(N__5672));
    InMux I__1186 (
            .O(N__5683),
            .I(N__5672));
    InMux I__1185 (
            .O(N__5682),
            .I(N__5669));
    InMux I__1184 (
            .O(N__5681),
            .I(N__5662));
    InMux I__1183 (
            .O(N__5678),
            .I(N__5662));
    InMux I__1182 (
            .O(N__5677),
            .I(N__5662));
    LocalMux I__1181 (
            .O(N__5672),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1180 (
            .O(N__5669),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    LocalMux I__1179 (
            .O(N__5662),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ));
    InMux I__1178 (
            .O(N__5655),
            .I(N__5646));
    InMux I__1177 (
            .O(N__5654),
            .I(N__5639));
    InMux I__1176 (
            .O(N__5653),
            .I(N__5639));
    InMux I__1175 (
            .O(N__5652),
            .I(N__5639));
    InMux I__1174 (
            .O(N__5651),
            .I(N__5632));
    InMux I__1173 (
            .O(N__5650),
            .I(N__5632));
    InMux I__1172 (
            .O(N__5649),
            .I(N__5632));
    LocalMux I__1171 (
            .O(N__5646),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1170 (
            .O(N__5639),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    LocalMux I__1169 (
            .O(N__5632),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ));
    InMux I__1168 (
            .O(N__5625),
            .I(N__5612));
    InMux I__1167 (
            .O(N__5624),
            .I(N__5612));
    InMux I__1166 (
            .O(N__5623),
            .I(N__5612));
    InMux I__1165 (
            .O(N__5622),
            .I(N__5609));
    InMux I__1164 (
            .O(N__5621),
            .I(N__5606));
    InMux I__1163 (
            .O(N__5620),
            .I(N__5601));
    InMux I__1162 (
            .O(N__5619),
            .I(N__5601));
    LocalMux I__1161 (
            .O(N__5612),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1160 (
            .O(N__5609),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1159 (
            .O(N__5606),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    LocalMux I__1158 (
            .O(N__5601),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ));
    CascadeMux I__1157 (
            .O(N__5592),
            .I(N__5587));
    CascadeMux I__1156 (
            .O(N__5591),
            .I(N__5584));
    InMux I__1155 (
            .O(N__5590),
            .I(N__5580));
    InMux I__1154 (
            .O(N__5587),
            .I(N__5575));
    InMux I__1153 (
            .O(N__5584),
            .I(N__5575));
    InMux I__1152 (
            .O(N__5583),
            .I(N__5572));
    LocalMux I__1151 (
            .O(N__5580),
            .I(N__5568));
    LocalMux I__1150 (
            .O(N__5575),
            .I(N__5563));
    LocalMux I__1149 (
            .O(N__5572),
            .I(N__5563));
    InMux I__1148 (
            .O(N__5571),
            .I(N__5560));
    Span4Mux_v I__1147 (
            .O(N__5568),
            .I(N__5555));
    Span4Mux_v I__1146 (
            .O(N__5563),
            .I(N__5555));
    LocalMux I__1145 (
            .O(N__5560),
            .I(N__5550));
    Sp12to4 I__1144 (
            .O(N__5555),
            .I(N__5550));
    Span12Mux_h I__1143 (
            .O(N__5550),
            .I(N__5547));
    Span12Mux_v I__1142 (
            .O(N__5547),
            .I(N__5544));
    Odrv12 I__1141 (
            .O(N__5544),
            .I(TSn_c));
    InMux I__1140 (
            .O(N__5541),
            .I(N__5538));
    LocalMux I__1139 (
            .O(N__5538),
            .I(N__5535));
    Span12Mux_h I__1138 (
            .O(N__5535),
            .I(N__5532));
    Odrv12 I__1137 (
            .O(N__5532),
            .I(U409_ADDRESS_DECODE_ROMEN_1));
    IoInMux I__1136 (
            .O(N__5529),
            .I(N__5525));
    CascadeMux I__1135 (
            .O(N__5528),
            .I(N__5520));
    LocalMux I__1134 (
            .O(N__5525),
            .I(N__5517));
    CascadeMux I__1133 (
            .O(N__5524),
            .I(N__5514));
    InMux I__1132 (
            .O(N__5523),
            .I(N__5511));
    InMux I__1131 (
            .O(N__5520),
            .I(N__5508));
    IoSpan4Mux I__1130 (
            .O(N__5517),
            .I(N__5504));
    InMux I__1129 (
            .O(N__5514),
            .I(N__5501));
    LocalMux I__1128 (
            .O(N__5511),
            .I(N__5496));
    LocalMux I__1127 (
            .O(N__5508),
            .I(N__5496));
    CascadeMux I__1126 (
            .O(N__5507),
            .I(N__5491));
    Span4Mux_s0_v I__1125 (
            .O(N__5504),
            .I(N__5487));
    LocalMux I__1124 (
            .O(N__5501),
            .I(N__5482));
    Span4Mux_v I__1123 (
            .O(N__5496),
            .I(N__5482));
    InMux I__1122 (
            .O(N__5495),
            .I(N__5477));
    InMux I__1121 (
            .O(N__5494),
            .I(N__5477));
    InMux I__1120 (
            .O(N__5491),
            .I(N__5474));
    InMux I__1119 (
            .O(N__5490),
            .I(N__5471));
    Sp12to4 I__1118 (
            .O(N__5487),
            .I(N__5468));
    Sp12to4 I__1117 (
            .O(N__5482),
            .I(N__5465));
    LocalMux I__1116 (
            .O(N__5477),
            .I(N__5462));
    LocalMux I__1115 (
            .O(N__5474),
            .I(N__5457));
    LocalMux I__1114 (
            .O(N__5471),
            .I(N__5457));
    Span12Mux_v I__1113 (
            .O(N__5468),
            .I(N__5450));
    Span12Mux_h I__1112 (
            .O(N__5465),
            .I(N__5450));
    Sp12to4 I__1111 (
            .O(N__5462),
            .I(N__5450));
    Sp12to4 I__1110 (
            .O(N__5457),
            .I(N__5447));
    Span12Mux_v I__1109 (
            .O(N__5450),
            .I(N__5444));
    Span12Mux_v I__1108 (
            .O(N__5447),
            .I(N__5441));
    Odrv12 I__1107 (
            .O(N__5444),
            .I(CLK40_IN_c));
    Odrv12 I__1106 (
            .O(N__5441),
            .I(CLK40_IN_c));
    InMux I__1105 (
            .O(N__5436),
            .I(N__5427));
    InMux I__1104 (
            .O(N__5435),
            .I(N__5418));
    InMux I__1103 (
            .O(N__5434),
            .I(N__5418));
    InMux I__1102 (
            .O(N__5433),
            .I(N__5418));
    InMux I__1101 (
            .O(N__5432),
            .I(N__5418));
    InMux I__1100 (
            .O(N__5431),
            .I(N__5415));
    InMux I__1099 (
            .O(N__5430),
            .I(N__5412));
    LocalMux I__1098 (
            .O(N__5427),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1097 (
            .O(N__5418),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1096 (
            .O(N__5415),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    LocalMux I__1095 (
            .O(N__5412),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ));
    InMux I__1094 (
            .O(N__5403),
            .I(N__5397));
    InMux I__1093 (
            .O(N__5402),
            .I(N__5397));
    LocalMux I__1092 (
            .O(N__5397),
            .I(\U409_TRANSFER_ACK.N_28_4 ));
    InMux I__1091 (
            .O(N__5394),
            .I(N__5389));
    InMux I__1090 (
            .O(N__5393),
            .I(N__5384));
    InMux I__1089 (
            .O(N__5392),
            .I(N__5384));
    LocalMux I__1088 (
            .O(N__5389),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    LocalMux I__1087 (
            .O(N__5384),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ));
    InMux I__1086 (
            .O(N__5379),
            .I(N__5376));
    LocalMux I__1085 (
            .O(N__5376),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ));
    CEMux I__1084 (
            .O(N__5373),
            .I(N__5370));
    LocalMux I__1083 (
            .O(N__5370),
            .I(N__5367));
    Odrv12 I__1082 (
            .O(N__5367),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_0 ));
    SRMux I__1081 (
            .O(N__5364),
            .I(N__5359));
    InMux I__1080 (
            .O(N__5363),
            .I(N__5355));
    SRMux I__1079 (
            .O(N__5362),
            .I(N__5352));
    LocalMux I__1078 (
            .O(N__5359),
            .I(N__5348));
    SRMux I__1077 (
            .O(N__5358),
            .I(N__5345));
    LocalMux I__1076 (
            .O(N__5355),
            .I(N__5340));
    LocalMux I__1075 (
            .O(N__5352),
            .I(N__5340));
    SRMux I__1074 (
            .O(N__5351),
            .I(N__5337));
    Span4Mux_v I__1073 (
            .O(N__5348),
            .I(N__5332));
    LocalMux I__1072 (
            .O(N__5345),
            .I(N__5332));
    Span4Mux_v I__1071 (
            .O(N__5340),
            .I(N__5327));
    LocalMux I__1070 (
            .O(N__5337),
            .I(N__5327));
    Odrv4 I__1069 (
            .O(N__5332),
            .I(RESETn_c_i));
    Odrv4 I__1068 (
            .O(N__5327),
            .I(RESETn_c_i));
    CascadeMux I__1067 (
            .O(N__5322),
            .I(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ));
    IoInMux I__1066 (
            .O(N__5319),
            .I(N__5316));
    LocalMux I__1065 (
            .O(N__5316),
            .I(N__5313));
    Span12Mux_s3_v I__1064 (
            .O(N__5313),
            .I(N__5310));
    Span12Mux_v I__1063 (
            .O(N__5310),
            .I(N__5305));
    InMux I__1062 (
            .O(N__5309),
            .I(N__5300));
    InMux I__1061 (
            .O(N__5308),
            .I(N__5300));
    Odrv12 I__1060 (
            .O(N__5305),
            .I(TACK_OUTn));
    LocalMux I__1059 (
            .O(N__5300),
            .I(TACK_OUTn));
    CascadeMux I__1058 (
            .O(N__5295),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_cascade_ ));
    InMux I__1057 (
            .O(N__5292),
            .I(N__5288));
    InMux I__1056 (
            .O(N__5291),
            .I(N__5285));
    LocalMux I__1055 (
            .O(N__5288),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    LocalMux I__1054 (
            .O(N__5285),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ));
    CascadeMux I__1053 (
            .O(N__5280),
            .I(N__5276));
    InMux I__1052 (
            .O(N__5279),
            .I(N__5273));
    InMux I__1051 (
            .O(N__5276),
            .I(N__5270));
    LocalMux I__1050 (
            .O(N__5273),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    LocalMux I__1049 (
            .O(N__5270),
            .I(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ));
    InMux I__1048 (
            .O(N__5265),
            .I(N__5261));
    InMux I__1047 (
            .O(N__5264),
            .I(N__5258));
    LocalMux I__1046 (
            .O(N__5261),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    LocalMux I__1045 (
            .O(N__5258),
            .I(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ));
    IoInMux I__1044 (
            .O(N__5253),
            .I(N__5250));
    LocalMux I__1043 (
            .O(N__5250),
            .I(N__5247));
    Span4Mux_s2_v I__1042 (
            .O(N__5247),
            .I(N__5244));
    Span4Mux_v I__1041 (
            .O(N__5244),
            .I(N__5241));
    Odrv4 I__1040 (
            .O(N__5241),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1039 (
            .O(N__5238),
            .I(N__5234));
    CascadeMux I__1038 (
            .O(N__5237),
            .I(N__5231));
    InMux I__1037 (
            .O(N__5234),
            .I(N__5228));
    InMux I__1036 (
            .O(N__5231),
            .I(N__5225));
    LocalMux I__1035 (
            .O(N__5228),
            .I(N__5220));
    LocalMux I__1034 (
            .O(N__5225),
            .I(N__5220));
    Span4Mux_v I__1033 (
            .O(N__5220),
            .I(N__5217));
    Span4Mux_h I__1032 (
            .O(N__5217),
            .I(N__5214));
    Odrv4 I__1031 (
            .O(N__5214),
            .I(\U409_TRANSFER_ACK.N_18 ));
    InMux I__1030 (
            .O(N__5211),
            .I(N__5208));
    LocalMux I__1029 (
            .O(N__5208),
            .I(\U409_TRANSFER_ACK.N_24 ));
    InMux I__1028 (
            .O(N__5205),
            .I(N__5202));
    LocalMux I__1027 (
            .O(N__5202),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_0 ));
    InMux I__1026 (
            .O(N__5199),
            .I(N__5196));
    LocalMux I__1025 (
            .O(N__5196),
            .I(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ));
    IoInMux I__1024 (
            .O(N__5193),
            .I(N__5190));
    LocalMux I__1023 (
            .O(N__5190),
            .I(N__5187));
    Span4Mux_s2_v I__1022 (
            .O(N__5187),
            .I(N__5184));
    Span4Mux_h I__1021 (
            .O(N__5184),
            .I(N__5181));
    Span4Mux_v I__1020 (
            .O(N__5181),
            .I(N__5177));
    CascadeMux I__1019 (
            .O(N__5180),
            .I(N__5174));
    Sp12to4 I__1018 (
            .O(N__5177),
            .I(N__5171));
    InMux I__1017 (
            .O(N__5174),
            .I(N__5168));
    Odrv12 I__1016 (
            .O(N__5171),
            .I(ROMENn_c));
    LocalMux I__1015 (
            .O(N__5168),
            .I(ROMENn_c));
    InMux I__1014 (
            .O(N__5163),
            .I(N__5160));
    LocalMux I__1013 (
            .O(N__5160),
            .I(N__5157));
    Span4Mux_v I__1012 (
            .O(N__5157),
            .I(N__5152));
    InMux I__1011 (
            .O(N__5156),
            .I(N__5149));
    InMux I__1010 (
            .O(N__5155),
            .I(N__5146));
    Odrv4 I__1009 (
            .O(N__5152),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__1008 (
            .O(N__5149),
            .I(\U409_CIA.VMAZ0 ));
    LocalMux I__1007 (
            .O(N__5146),
            .I(\U409_CIA.VMAZ0 ));
    InMux I__1006 (
            .O(N__5139),
            .I(N__5133));
    InMux I__1005 (
            .O(N__5138),
            .I(N__5126));
    InMux I__1004 (
            .O(N__5137),
            .I(N__5126));
    InMux I__1003 (
            .O(N__5136),
            .I(N__5126));
    LocalMux I__1002 (
            .O(N__5133),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    LocalMux I__1001 (
            .O(N__5126),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ));
    InMux I__1000 (
            .O(N__5121),
            .I(N__5115));
    InMux I__999 (
            .O(N__5120),
            .I(N__5112));
    InMux I__998 (
            .O(N__5119),
            .I(N__5107));
    InMux I__997 (
            .O(N__5118),
            .I(N__5107));
    LocalMux I__996 (
            .O(N__5115),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__995 (
            .O(N__5112),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    LocalMux I__994 (
            .O(N__5107),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ));
    InMux I__993 (
            .O(N__5100),
            .I(N__5095));
    InMux I__992 (
            .O(N__5099),
            .I(N__5090));
    InMux I__991 (
            .O(N__5098),
            .I(N__5090));
    LocalMux I__990 (
            .O(N__5095),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    LocalMux I__989 (
            .O(N__5090),
            .I(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ));
    CascadeMux I__988 (
            .O(N__5085),
            .I(N__5082));
    InMux I__987 (
            .O(N__5082),
            .I(N__5079));
    LocalMux I__986 (
            .O(N__5079),
            .I(\U409_TRANSFER_ACK.ROM_TACK_EN_e_1 ));
    InMux I__985 (
            .O(N__5076),
            .I(N__5072));
    InMux I__984 (
            .O(N__5075),
            .I(N__5069));
    LocalMux I__983 (
            .O(N__5072),
            .I(N__5062));
    LocalMux I__982 (
            .O(N__5069),
            .I(N__5062));
    InMux I__981 (
            .O(N__5068),
            .I(N__5057));
    InMux I__980 (
            .O(N__5067),
            .I(N__5057));
    Odrv4 I__979 (
            .O(N__5062),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    LocalMux I__978 (
            .O(N__5057),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ));
    InMux I__977 (
            .O(N__5052),
            .I(N__5045));
    InMux I__976 (
            .O(N__5051),
            .I(N__5042));
    InMux I__975 (
            .O(N__5050),
            .I(N__5039));
    InMux I__974 (
            .O(N__5049),
            .I(N__5034));
    InMux I__973 (
            .O(N__5048),
            .I(N__5034));
    LocalMux I__972 (
            .O(N__5045),
            .I(N__5029));
    LocalMux I__971 (
            .O(N__5042),
            .I(N__5029));
    LocalMux I__970 (
            .O(N__5039),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    LocalMux I__969 (
            .O(N__5034),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    Odrv4 I__968 (
            .O(N__5029),
            .I(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ));
    CascadeMux I__967 (
            .O(N__5022),
            .I(N__5019));
    InMux I__966 (
            .O(N__5019),
            .I(N__5016));
    LocalMux I__965 (
            .O(N__5016),
            .I(\U409_TRANSFER_ACK.N_138 ));
    InMux I__964 (
            .O(N__5013),
            .I(N__5007));
    InMux I__963 (
            .O(N__5012),
            .I(N__5007));
    LocalMux I__962 (
            .O(N__5007),
            .I(N__5004));
    Span4Mux_v I__961 (
            .O(N__5004),
            .I(N__5001));
    Sp12to4 I__960 (
            .O(N__5001),
            .I(N__4998));
    Odrv12 I__959 (
            .O(N__4998),
            .I(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_0 ));
    SRMux I__958 (
            .O(N__4995),
            .I(N__4991));
    SRMux I__957 (
            .O(N__4994),
            .I(N__4988));
    LocalMux I__956 (
            .O(N__4991),
            .I(N__4982));
    LocalMux I__955 (
            .O(N__4988),
            .I(N__4982));
    SRMux I__954 (
            .O(N__4987),
            .I(N__4979));
    Span4Mux_v I__953 (
            .O(N__4982),
            .I(N__4976));
    LocalMux I__952 (
            .O(N__4979),
            .I(N__4973));
    Sp12to4 I__951 (
            .O(N__4976),
            .I(N__4970));
    Sp12to4 I__950 (
            .O(N__4973),
            .I(N__4967));
    Odrv12 I__949 (
            .O(N__4970),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    Odrv12 I__948 (
            .O(N__4967),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ));
    CascadeMux I__947 (
            .O(N__4962),
            .I(\U409_TRANSFER_ACK.m8_ns_1_cascade_ ));
    CascadeMux I__946 (
            .O(N__4959),
            .I(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ));
    InMux I__945 (
            .O(N__4956),
            .I(N__4953));
    LocalMux I__944 (
            .O(N__4953),
            .I(\U409_TRANSFER_ACK.N_9 ));
    InMux I__943 (
            .O(N__4950),
            .I(N__4947));
    LocalMux I__942 (
            .O(N__4947),
            .I(\U409_TRANSFER_ACK.N_4 ));
    CascadeMux I__941 (
            .O(N__4944),
            .I(\U409_TRANSFER_ACK.N_4_cascade_ ));
    InMux I__940 (
            .O(N__4941),
            .I(N__4938));
    LocalMux I__939 (
            .O(N__4938),
            .I(\U409_TRANSFER_ACK.N_5 ));
    CascadeMux I__938 (
            .O(N__4935),
            .I(N__4932));
    InMux I__937 (
            .O(N__4932),
            .I(N__4923));
    InMux I__936 (
            .O(N__4931),
            .I(N__4923));
    InMux I__935 (
            .O(N__4930),
            .I(N__4923));
    LocalMux I__934 (
            .O(N__4923),
            .I(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ));
    IoInMux I__933 (
            .O(N__4920),
            .I(N__4917));
    LocalMux I__932 (
            .O(N__4917),
            .I(N__4914));
    IoSpan4Mux I__931 (
            .O(N__4914),
            .I(N__4911));
    Sp12to4 I__930 (
            .O(N__4911),
            .I(N__4908));
    Span12Mux_s6_v I__929 (
            .O(N__4908),
            .I(N__4905));
    Span12Mux_v I__928 (
            .O(N__4905),
            .I(N__4900));
    InMux I__927 (
            .O(N__4904),
            .I(N__4897));
    InMux I__926 (
            .O(N__4903),
            .I(N__4894));
    Odrv12 I__925 (
            .O(N__4900),
            .I(CLK_CIA_c));
    LocalMux I__924 (
            .O(N__4897),
            .I(CLK_CIA_c));
    LocalMux I__923 (
            .O(N__4894),
            .I(CLK_CIA_c));
    CascadeMux I__922 (
            .O(N__4887),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ));
    InMux I__921 (
            .O(N__4884),
            .I(N__4881));
    LocalMux I__920 (
            .O(N__4881),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ));
    InMux I__919 (
            .O(N__4878),
            .I(N__4873));
    InMux I__918 (
            .O(N__4877),
            .I(N__4868));
    InMux I__917 (
            .O(N__4876),
            .I(N__4868));
    LocalMux I__916 (
            .O(N__4873),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    LocalMux I__915 (
            .O(N__4868),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ));
    CascadeMux I__914 (
            .O(N__4863),
            .I(N__4858));
    InMux I__913 (
            .O(N__4862),
            .I(N__4852));
    InMux I__912 (
            .O(N__4861),
            .I(N__4852));
    InMux I__911 (
            .O(N__4858),
            .I(N__4847));
    InMux I__910 (
            .O(N__4857),
            .I(N__4847));
    LocalMux I__909 (
            .O(N__4852),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    LocalMux I__908 (
            .O(N__4847),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ));
    CascadeMux I__907 (
            .O(N__4842),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_6_cascade_ ));
    InMux I__906 (
            .O(N__4839),
            .I(N__4836));
    LocalMux I__905 (
            .O(N__4836),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1 ));
    InMux I__904 (
            .O(N__4833),
            .I(N__4830));
    LocalMux I__903 (
            .O(N__4830),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ));
    CascadeMux I__902 (
            .O(N__4827),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ));
    InMux I__901 (
            .O(N__4824),
            .I(N__4817));
    InMux I__900 (
            .O(N__4823),
            .I(N__4817));
    InMux I__899 (
            .O(N__4822),
            .I(N__4813));
    LocalMux I__898 (
            .O(N__4817),
            .I(N__4810));
    InMux I__897 (
            .O(N__4816),
            .I(N__4807));
    LocalMux I__896 (
            .O(N__4813),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    Odrv4 I__895 (
            .O(N__4810),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    LocalMux I__894 (
            .O(N__4807),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ));
    InMux I__893 (
            .O(N__4800),
            .I(N__4793));
    InMux I__892 (
            .O(N__4799),
            .I(N__4793));
    InMux I__891 (
            .O(N__4798),
            .I(N__4790));
    LocalMux I__890 (
            .O(N__4793),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    LocalMux I__889 (
            .O(N__4790),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ));
    InMux I__888 (
            .O(N__4785),
            .I(N__4775));
    InMux I__887 (
            .O(N__4784),
            .I(N__4775));
    InMux I__886 (
            .O(N__4783),
            .I(N__4772));
    InMux I__885 (
            .O(N__4782),
            .I(N__4765));
    InMux I__884 (
            .O(N__4781),
            .I(N__4765));
    InMux I__883 (
            .O(N__4780),
            .I(N__4765));
    LocalMux I__882 (
            .O(N__4775),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__881 (
            .O(N__4772),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    LocalMux I__880 (
            .O(N__4765),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ));
    CascadeMux I__879 (
            .O(N__4758),
            .I(N__4753));
    CascadeMux I__878 (
            .O(N__4757),
            .I(N__4750));
    InMux I__877 (
            .O(N__4756),
            .I(N__4746));
    InMux I__876 (
            .O(N__4753),
            .I(N__4739));
    InMux I__875 (
            .O(N__4750),
            .I(N__4739));
    InMux I__874 (
            .O(N__4749),
            .I(N__4739));
    LocalMux I__873 (
            .O(N__4746),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    LocalMux I__872 (
            .O(N__4739),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ));
    InMux I__871 (
            .O(N__4734),
            .I(N__4729));
    InMux I__870 (
            .O(N__4733),
            .I(N__4726));
    InMux I__869 (
            .O(N__4732),
            .I(N__4723));
    LocalMux I__868 (
            .O(N__4729),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__867 (
            .O(N__4726),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    LocalMux I__866 (
            .O(N__4723),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ));
    InMux I__865 (
            .O(N__4716),
            .I(N__4704));
    InMux I__864 (
            .O(N__4715),
            .I(N__4704));
    InMux I__863 (
            .O(N__4714),
            .I(N__4704));
    InMux I__862 (
            .O(N__4713),
            .I(N__4697));
    InMux I__861 (
            .O(N__4712),
            .I(N__4697));
    InMux I__860 (
            .O(N__4711),
            .I(N__4697));
    LocalMux I__859 (
            .O(N__4704),
            .I(N__4694));
    LocalMux I__858 (
            .O(N__4697),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    Odrv4 I__857 (
            .O(N__4694),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ));
    CascadeMux I__856 (
            .O(N__4689),
            .I(N__4683));
    CascadeMux I__855 (
            .O(N__4688),
            .I(N__4679));
    CascadeMux I__854 (
            .O(N__4687),
            .I(N__4676));
    InMux I__853 (
            .O(N__4686),
            .I(N__4668));
    InMux I__852 (
            .O(N__4683),
            .I(N__4668));
    InMux I__851 (
            .O(N__4682),
            .I(N__4668));
    InMux I__850 (
            .O(N__4679),
            .I(N__4661));
    InMux I__849 (
            .O(N__4676),
            .I(N__4661));
    InMux I__848 (
            .O(N__4675),
            .I(N__4661));
    LocalMux I__847 (
            .O(N__4668),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    LocalMux I__846 (
            .O(N__4661),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ));
    InMux I__845 (
            .O(N__4656),
            .I(N__4647));
    InMux I__844 (
            .O(N__4655),
            .I(N__4647));
    InMux I__843 (
            .O(N__4654),
            .I(N__4640));
    InMux I__842 (
            .O(N__4653),
            .I(N__4640));
    InMux I__841 (
            .O(N__4652),
            .I(N__4640));
    LocalMux I__840 (
            .O(N__4647),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    LocalMux I__839 (
            .O(N__4640),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ));
    InMux I__838 (
            .O(N__4635),
            .I(N__4628));
    InMux I__837 (
            .O(N__4634),
            .I(N__4621));
    InMux I__836 (
            .O(N__4633),
            .I(N__4621));
    InMux I__835 (
            .O(N__4632),
            .I(N__4621));
    InMux I__834 (
            .O(N__4631),
            .I(N__4618));
    LocalMux I__833 (
            .O(N__4628),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__832 (
            .O(N__4621),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    LocalMux I__831 (
            .O(N__4618),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ));
    CascadeMux I__830 (
            .O(N__4611),
            .I(N__4606));
    InMux I__829 (
            .O(N__4610),
            .I(N__4601));
    InMux I__828 (
            .O(N__4609),
            .I(N__4594));
    InMux I__827 (
            .O(N__4606),
            .I(N__4594));
    InMux I__826 (
            .O(N__4605),
            .I(N__4594));
    InMux I__825 (
            .O(N__4604),
            .I(N__4591));
    LocalMux I__824 (
            .O(N__4601),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__823 (
            .O(N__4594),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    LocalMux I__822 (
            .O(N__4591),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ));
    ClkMux I__821 (
            .O(N__4584),
            .I(N__4572));
    ClkMux I__820 (
            .O(N__4583),
            .I(N__4572));
    ClkMux I__819 (
            .O(N__4582),
            .I(N__4572));
    ClkMux I__818 (
            .O(N__4581),
            .I(N__4572));
    GlobalMux I__817 (
            .O(N__4572),
            .I(N__4569));
    gio2CtrlBuf I__816 (
            .O(N__4569),
            .I(CLK28_IN_c_g));
    InMux I__815 (
            .O(N__4566),
            .I(N__4560));
    InMux I__814 (
            .O(N__4565),
            .I(N__4557));
    InMux I__813 (
            .O(N__4564),
            .I(N__4554));
    InMux I__812 (
            .O(N__4563),
            .I(N__4551));
    LocalMux I__811 (
            .O(N__4560),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__810 (
            .O(N__4557),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__809 (
            .O(N__4554),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    LocalMux I__808 (
            .O(N__4551),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ));
    CascadeMux I__807 (
            .O(N__4542),
            .I(N__4534));
    InMux I__806 (
            .O(N__4541),
            .I(N__4531));
    InMux I__805 (
            .O(N__4540),
            .I(N__4526));
    InMux I__804 (
            .O(N__4539),
            .I(N__4526));
    InMux I__803 (
            .O(N__4538),
            .I(N__4523));
    InMux I__802 (
            .O(N__4537),
            .I(N__4520));
    InMux I__801 (
            .O(N__4534),
            .I(N__4517));
    LocalMux I__800 (
            .O(N__4531),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__799 (
            .O(N__4526),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__798 (
            .O(N__4523),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__797 (
            .O(N__4520),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    LocalMux I__796 (
            .O(N__4517),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ));
    CascadeMux I__795 (
            .O(N__4506),
            .I(N__4500));
    CascadeMux I__794 (
            .O(N__4505),
            .I(N__4497));
    InMux I__793 (
            .O(N__4504),
            .I(N__4494));
    InMux I__792 (
            .O(N__4503),
            .I(N__4491));
    InMux I__791 (
            .O(N__4500),
            .I(N__4488));
    InMux I__790 (
            .O(N__4497),
            .I(N__4485));
    LocalMux I__789 (
            .O(N__4494),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__788 (
            .O(N__4491),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__787 (
            .O(N__4488),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    LocalMux I__786 (
            .O(N__4485),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ));
    InMux I__785 (
            .O(N__4476),
            .I(N__4468));
    InMux I__784 (
            .O(N__4475),
            .I(N__4468));
    CascadeMux I__783 (
            .O(N__4474),
            .I(N__4465));
    InMux I__782 (
            .O(N__4473),
            .I(N__4460));
    LocalMux I__781 (
            .O(N__4468),
            .I(N__4457));
    InMux I__780 (
            .O(N__4465),
            .I(N__4454));
    InMux I__779 (
            .O(N__4464),
            .I(N__4451));
    InMux I__778 (
            .O(N__4463),
            .I(N__4448));
    LocalMux I__777 (
            .O(N__4460),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    Odrv12 I__776 (
            .O(N__4457),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__775 (
            .O(N__4454),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__774 (
            .O(N__4451),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    LocalMux I__773 (
            .O(N__4448),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ));
    InMux I__772 (
            .O(N__4437),
            .I(N__4434));
    LocalMux I__771 (
            .O(N__4434),
            .I(N__4431));
    Odrv4 I__770 (
            .O(N__4431),
            .I(\U409_CIA.CLK_CIA6_3 ));
    CascadeMux I__769 (
            .O(N__4428),
            .I(N__4425));
    InMux I__768 (
            .O(N__4425),
            .I(N__4421));
    CascadeMux I__767 (
            .O(N__4424),
            .I(N__4417));
    LocalMux I__766 (
            .O(N__4421),
            .I(N__4412));
    InMux I__765 (
            .O(N__4420),
            .I(N__4407));
    InMux I__764 (
            .O(N__4417),
            .I(N__4407));
    InMux I__763 (
            .O(N__4416),
            .I(N__4404));
    InMux I__762 (
            .O(N__4415),
            .I(N__4401));
    Odrv4 I__761 (
            .O(N__4412),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__760 (
            .O(N__4407),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__759 (
            .O(N__4404),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    LocalMux I__758 (
            .O(N__4401),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ));
    InMux I__757 (
            .O(N__4392),
            .I(N__4389));
    LocalMux I__756 (
            .O(N__4389),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_2_1 ));
    CascadeMux I__755 (
            .O(N__4386),
            .I(\U409_CIA.CLK_CIA6_3_cascade_ ));
    InMux I__754 (
            .O(N__4383),
            .I(N__4374));
    InMux I__753 (
            .O(N__4382),
            .I(N__4374));
    InMux I__752 (
            .O(N__4381),
            .I(N__4371));
    InMux I__751 (
            .O(N__4380),
            .I(N__4368));
    InMux I__750 (
            .O(N__4379),
            .I(N__4365));
    LocalMux I__749 (
            .O(N__4374),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__748 (
            .O(N__4371),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__747 (
            .O(N__4368),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    LocalMux I__746 (
            .O(N__4365),
            .I(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ));
    InMux I__745 (
            .O(N__4356),
            .I(N__4353));
    LocalMux I__744 (
            .O(N__4353),
            .I(\U409_CIA.CLK_CIA_RNOZ0Z_1 ));
    InMux I__743 (
            .O(N__4350),
            .I(N__4345));
    InMux I__742 (
            .O(N__4349),
            .I(N__4342));
    InMux I__741 (
            .O(N__4348),
            .I(N__4339));
    LocalMux I__740 (
            .O(N__4345),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__739 (
            .O(N__4342),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    LocalMux I__738 (
            .O(N__4339),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ));
    CascadeMux I__737 (
            .O(N__4332),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ));
    InMux I__736 (
            .O(N__4329),
            .I(N__4326));
    LocalMux I__735 (
            .O(N__4326),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ));
    InMux I__734 (
            .O(N__4323),
            .I(N__4320));
    LocalMux I__733 (
            .O(N__4320),
            .I(N__4317));
    Span12Mux_h I__732 (
            .O(N__4317),
            .I(N__4314));
    Odrv12 I__731 (
            .O(N__4314),
            .I(A_c_12));
    IoInMux I__730 (
            .O(N__4311),
            .I(N__4308));
    LocalMux I__729 (
            .O(N__4308),
            .I(N__4305));
    Span4Mux_s0_h I__728 (
            .O(N__4305),
            .I(N__4302));
    Sp12to4 I__727 (
            .O(N__4302),
            .I(N__4299));
    Span12Mux_s10_v I__726 (
            .O(N__4299),
            .I(N__4296));
    Span12Mux_h I__725 (
            .O(N__4296),
            .I(N__4293));
    Odrv12 I__724 (
            .O(N__4293),
            .I(U409_ADDRESS_DECODE_un1_CIACS0n_i));
    InMux I__723 (
            .O(N__4290),
            .I(N__4287));
    LocalMux I__722 (
            .O(N__4287),
            .I(N__4283));
    InMux I__721 (
            .O(N__4286),
            .I(N__4280));
    Odrv4 I__720 (
            .O(N__4283),
            .I(CIA_ENABLE));
    LocalMux I__719 (
            .O(N__4280),
            .I(CIA_ENABLE));
    InMux I__718 (
            .O(N__4275),
            .I(N__4271));
    InMux I__717 (
            .O(N__4274),
            .I(N__4268));
    LocalMux I__716 (
            .O(N__4271),
            .I(\U409_CIA.CLK_CIA6_0 ));
    LocalMux I__715 (
            .O(N__4268),
            .I(\U409_CIA.CLK_CIA6_0 ));
    CascadeMux I__714 (
            .O(N__4263),
            .I(\U409_CIA.CLK_CIA6_cascade_ ));
    InMux I__713 (
            .O(N__4260),
            .I(N__4257));
    LocalMux I__712 (
            .O(N__4257),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ));
    InMux I__711 (
            .O(N__4254),
            .I(N__4251));
    LocalMux I__710 (
            .O(N__4251),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0 ));
    CascadeMux I__709 (
            .O(N__4248),
            .I(\U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ));
    InMux I__708 (
            .O(N__4245),
            .I(N__4242));
    LocalMux I__707 (
            .O(N__4242),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO ));
    CascadeMux I__706 (
            .O(N__4239),
            .I(N__4235));
    InMux I__705 (
            .O(N__4238),
            .I(N__4230));
    InMux I__704 (
            .O(N__4235),
            .I(N__4230));
    LocalMux I__703 (
            .O(N__4230),
            .I(\U409_CIA.CIA_CLK_COUNT11_3 ));
    InMux I__702 (
            .O(N__4227),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ));
    CascadeMux I__701 (
            .O(N__4224),
            .I(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_ ));
    CascadeMux I__700 (
            .O(N__4221),
            .I(N__4218));
    InMux I__699 (
            .O(N__4218),
            .I(N__4212));
    InMux I__698 (
            .O(N__4217),
            .I(N__4212));
    LocalMux I__697 (
            .O(N__4212),
            .I(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ));
    InMux I__696 (
            .O(N__4209),
            .I(N__4204));
    InMux I__695 (
            .O(N__4208),
            .I(N__4201));
    InMux I__694 (
            .O(N__4207),
            .I(N__4198));
    LocalMux I__693 (
            .O(N__4204),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    LocalMux I__692 (
            .O(N__4201),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    LocalMux I__691 (
            .O(N__4198),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn));
    InMux I__690 (
            .O(N__4191),
            .I(N__4188));
    LocalMux I__689 (
            .O(N__4188),
            .I(N__4185));
    Odrv4 I__688 (
            .O(N__4185),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn));
    InMux I__687 (
            .O(N__4182),
            .I(N__4179));
    LocalMux I__686 (
            .O(N__4179),
            .I(N__4176));
    Span12Mux_h I__685 (
            .O(N__4176),
            .I(N__4173));
    Span12Mux_h I__684 (
            .O(N__4173),
            .I(N__4170));
    Span12Mux_v I__683 (
            .O(N__4170),
            .I(N__4167));
    Odrv12 I__682 (
            .O(N__4167),
            .I(TACKn_in));
    InMux I__681 (
            .O(N__4164),
            .I(N__4161));
    LocalMux I__680 (
            .O(N__4161),
            .I(N__4158));
    Span12Mux_v I__679 (
            .O(N__4158),
            .I(N__4155));
    Span12Mux_h I__678 (
            .O(N__4155),
            .I(N__4152));
    Odrv12 I__677 (
            .O(N__4152),
            .I(A_c_13));
    IoInMux I__676 (
            .O(N__4149),
            .I(N__4146));
    LocalMux I__675 (
            .O(N__4146),
            .I(N__4143));
    Span4Mux_s0_h I__674 (
            .O(N__4143),
            .I(N__4140));
    Sp12to4 I__673 (
            .O(N__4140),
            .I(N__4137));
    Span12Mux_s9_v I__672 (
            .O(N__4137),
            .I(N__4134));
    Span12Mux_h I__671 (
            .O(N__4134),
            .I(N__4131));
    Odrv12 I__670 (
            .O(N__4131),
            .I(U409_ADDRESS_DECODE_un1_CIACS1n_i));
    InMux I__669 (
            .O(N__4128),
            .I(N__4125));
    LocalMux I__668 (
            .O(N__4125),
            .I(N__4121));
    InMux I__667 (
            .O(N__4124),
            .I(N__4118));
    Span12Mux_h I__666 (
            .O(N__4121),
            .I(N__4115));
    LocalMux I__665 (
            .O(N__4118),
            .I(N__4112));
    Odrv12 I__664 (
            .O(N__4115),
            .I(CIA_SPACE));
    Odrv4 I__663 (
            .O(N__4112),
            .I(CIA_SPACE));
    CascadeMux I__662 (
            .O(N__4107),
            .I(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ));
    InMux I__661 (
            .O(N__4104),
            .I(N__4101));
    LocalMux I__660 (
            .O(N__4101),
            .I(\U409_CIA.un1_CIA_CLK_COUNT_3_1 ));
    InMux I__659 (
            .O(N__4098),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ));
    InMux I__658 (
            .O(N__4095),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ));
    InMux I__657 (
            .O(N__4092),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ));
    InMux I__656 (
            .O(N__4089),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ));
    InMux I__655 (
            .O(N__4086),
            .I(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ));
    InMux I__654 (
            .O(N__4083),
            .I(N__4080));
    LocalMux I__653 (
            .O(N__4080),
            .I(N__4076));
    InMux I__652 (
            .O(N__4079),
            .I(N__4073));
    Span4Mux_v I__651 (
            .O(N__4076),
            .I(N__4070));
    LocalMux I__650 (
            .O(N__4073),
            .I(N__4067));
    Sp12to4 I__649 (
            .O(N__4070),
            .I(N__4064));
    Sp12to4 I__648 (
            .O(N__4067),
            .I(N__4061));
    Span12Mux_h I__647 (
            .O(N__4064),
            .I(N__4058));
    Span12Mux_v I__646 (
            .O(N__4061),
            .I(N__4055));
    Span12Mux_v I__645 (
            .O(N__4058),
            .I(N__4050));
    Span12Mux_h I__644 (
            .O(N__4055),
            .I(N__4050));
    Odrv12 I__643 (
            .O(N__4050),
            .I(OVL_c));
    CascadeMux I__642 (
            .O(N__4047),
            .I(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0_cascade_ ));
    IoInMux I__641 (
            .O(N__4044),
            .I(N__4041));
    LocalMux I__640 (
            .O(N__4041),
            .I(N__4038));
    Span4Mux_s3_v I__639 (
            .O(N__4038),
            .I(N__4035));
    Sp12to4 I__638 (
            .O(N__4035),
            .I(N__4032));
    Span12Mux_h I__637 (
            .O(N__4032),
            .I(N__4029));
    Span12Mux_v I__636 (
            .O(N__4029),
            .I(N__4026));
    Odrv12 I__635 (
            .O(N__4026),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn_i));
    InMux I__634 (
            .O(N__4023),
            .I(N__4020));
    LocalMux I__633 (
            .O(N__4020),
            .I(N__4016));
    InMux I__632 (
            .O(N__4019),
            .I(N__4013));
    Span4Mux_v I__631 (
            .O(N__4016),
            .I(N__4010));
    LocalMux I__630 (
            .O(N__4013),
            .I(N__4007));
    Odrv4 I__629 (
            .O(N__4010),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn));
    Odrv4 I__628 (
            .O(N__4007),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn));
    IoInMux I__627 (
            .O(N__4002),
            .I(N__3999));
    LocalMux I__626 (
            .O(N__3999),
            .I(N__3996));
    Span4Mux_s2_v I__625 (
            .O(N__3996),
            .I(N__3993));
    Sp12to4 I__624 (
            .O(N__3993),
            .I(N__3990));
    Span12Mux_h I__623 (
            .O(N__3990),
            .I(N__3987));
    Span12Mux_v I__622 (
            .O(N__3987),
            .I(N__3984));
    Odrv12 I__621 (
            .O(N__3984),
            .I(PORTSIZE_0_i));
    InMux I__620 (
            .O(N__3981),
            .I(N__3972));
    InMux I__619 (
            .O(N__3980),
            .I(N__3965));
    InMux I__618 (
            .O(N__3979),
            .I(N__3965));
    InMux I__617 (
            .O(N__3978),
            .I(N__3965));
    InMux I__616 (
            .O(N__3977),
            .I(N__3960));
    InMux I__615 (
            .O(N__3976),
            .I(N__3955));
    InMux I__614 (
            .O(N__3975),
            .I(N__3955));
    LocalMux I__613 (
            .O(N__3972),
            .I(N__3950));
    LocalMux I__612 (
            .O(N__3965),
            .I(N__3950));
    InMux I__611 (
            .O(N__3964),
            .I(N__3947));
    InMux I__610 (
            .O(N__3963),
            .I(N__3944));
    LocalMux I__609 (
            .O(N__3960),
            .I(N__3939));
    LocalMux I__608 (
            .O(N__3955),
            .I(N__3939));
    Span4Mux_h I__607 (
            .O(N__3950),
            .I(N__3932));
    LocalMux I__606 (
            .O(N__3947),
            .I(N__3932));
    LocalMux I__605 (
            .O(N__3944),
            .I(N__3932));
    Span4Mux_v I__604 (
            .O(N__3939),
            .I(N__3929));
    Span4Mux_v I__603 (
            .O(N__3932),
            .I(N__3926));
    Sp12to4 I__602 (
            .O(N__3929),
            .I(N__3921));
    Sp12to4 I__601 (
            .O(N__3926),
            .I(N__3921));
    Odrv12 I__600 (
            .O(N__3921),
            .I(A_c_23));
    InMux I__599 (
            .O(N__3918),
            .I(N__3915));
    LocalMux I__598 (
            .O(N__3915),
            .I(N__3912));
    Odrv4 I__597 (
            .O(N__3912),
            .I(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0 ));
    CascadeMux I__596 (
            .O(N__3909),
            .I(N__3906));
    InMux I__595 (
            .O(N__3906),
            .I(N__3903));
    LocalMux I__594 (
            .O(N__3903),
            .I(N__3895));
    InMux I__593 (
            .O(N__3902),
            .I(N__3889));
    InMux I__592 (
            .O(N__3901),
            .I(N__3889));
    InMux I__591 (
            .O(N__3900),
            .I(N__3884));
    InMux I__590 (
            .O(N__3899),
            .I(N__3884));
    InMux I__589 (
            .O(N__3898),
            .I(N__3881));
    Span4Mux_v I__588 (
            .O(N__3895),
            .I(N__3878));
    InMux I__587 (
            .O(N__3894),
            .I(N__3872));
    LocalMux I__586 (
            .O(N__3889),
            .I(N__3865));
    LocalMux I__585 (
            .O(N__3884),
            .I(N__3865));
    LocalMux I__584 (
            .O(N__3881),
            .I(N__3865));
    Span4Mux_v I__583 (
            .O(N__3878),
            .I(N__3862));
    InMux I__582 (
            .O(N__3877),
            .I(N__3857));
    InMux I__581 (
            .O(N__3876),
            .I(N__3857));
    InMux I__580 (
            .O(N__3875),
            .I(N__3854));
    LocalMux I__579 (
            .O(N__3872),
            .I(N__3851));
    Span12Mux_h I__578 (
            .O(N__3865),
            .I(N__3848));
    Span4Mux_v I__577 (
            .O(N__3862),
            .I(N__3845));
    LocalMux I__576 (
            .O(N__3857),
            .I(N__3838));
    LocalMux I__575 (
            .O(N__3854),
            .I(N__3838));
    Sp12to4 I__574 (
            .O(N__3851),
            .I(N__3838));
    Span12Mux_v I__573 (
            .O(N__3848),
            .I(N__3835));
    Sp12to4 I__572 (
            .O(N__3845),
            .I(N__3830));
    Span12Mux_v I__571 (
            .O(N__3838),
            .I(N__3830));
    Odrv12 I__570 (
            .O(N__3835),
            .I(A_c_22));
    Odrv12 I__569 (
            .O(N__3830),
            .I(A_c_22));
    CascadeMux I__568 (
            .O(N__3825),
            .I(N__3820));
    InMux I__567 (
            .O(N__3824),
            .I(N__3813));
    InMux I__566 (
            .O(N__3823),
            .I(N__3808));
    InMux I__565 (
            .O(N__3820),
            .I(N__3808));
    InMux I__564 (
            .O(N__3819),
            .I(N__3802));
    InMux I__563 (
            .O(N__3818),
            .I(N__3799));
    InMux I__562 (
            .O(N__3817),
            .I(N__3794));
    InMux I__561 (
            .O(N__3816),
            .I(N__3794));
    LocalMux I__560 (
            .O(N__3813),
            .I(N__3791));
    LocalMux I__559 (
            .O(N__3808),
            .I(N__3788));
    InMux I__558 (
            .O(N__3807),
            .I(N__3783));
    InMux I__557 (
            .O(N__3806),
            .I(N__3783));
    InMux I__556 (
            .O(N__3805),
            .I(N__3780));
    LocalMux I__555 (
            .O(N__3802),
            .I(N__3773));
    LocalMux I__554 (
            .O(N__3799),
            .I(N__3773));
    LocalMux I__553 (
            .O(N__3794),
            .I(N__3773));
    Span4Mux_h I__552 (
            .O(N__3791),
            .I(N__3764));
    Span4Mux_h I__551 (
            .O(N__3788),
            .I(N__3764));
    LocalMux I__550 (
            .O(N__3783),
            .I(N__3764));
    LocalMux I__549 (
            .O(N__3780),
            .I(N__3764));
    Span4Mux_v I__548 (
            .O(N__3773),
            .I(N__3761));
    Span4Mux_v I__547 (
            .O(N__3764),
            .I(N__3758));
    Sp12to4 I__546 (
            .O(N__3761),
            .I(N__3753));
    Sp12to4 I__545 (
            .O(N__3758),
            .I(N__3753));
    Odrv12 I__544 (
            .O(N__3753),
            .I(A_c_21));
    CascadeMux I__543 (
            .O(N__3750),
            .I(U409_ADDRESS_DECODE_un1_RAMSPACEn_cascade_));
    InMux I__542 (
            .O(N__3747),
            .I(N__3744));
    LocalMux I__541 (
            .O(N__3744),
            .I(U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_5));
    InMux I__540 (
            .O(N__3741),
            .I(N__3738));
    LocalMux I__539 (
            .O(N__3738),
            .I(N__3735));
    Odrv4 I__538 (
            .O(N__3735),
            .I(U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_7));
    CascadeMux I__537 (
            .O(N__3732),
            .I(AGNUS_SPACE_0_cascade_));
    InMux I__536 (
            .O(N__3729),
            .I(N__3726));
    LocalMux I__535 (
            .O(N__3726),
            .I(N__3723));
    Span4Mux_v I__534 (
            .O(N__3723),
            .I(N__3720));
    Odrv4 I__533 (
            .O(N__3720),
            .I(U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_6));
    IoInMux I__532 (
            .O(N__3717),
            .I(N__3714));
    LocalMux I__531 (
            .O(N__3714),
            .I(N__3711));
    Span4Mux_s3_v I__530 (
            .O(N__3711),
            .I(N__3708));
    Span4Mux_h I__529 (
            .O(N__3708),
            .I(N__3705));
    Sp12to4 I__528 (
            .O(N__3705),
            .I(N__3702));
    Span12Mux_h I__527 (
            .O(N__3702),
            .I(N__3699));
    Odrv12 I__526 (
            .O(N__3699),
            .I(BUFENn_c));
    InMux I__525 (
            .O(N__3696),
            .I(N__3689));
    InMux I__524 (
            .O(N__3695),
            .I(N__3689));
    InMux I__523 (
            .O(N__3694),
            .I(N__3686));
    LocalMux I__522 (
            .O(N__3689),
            .I(N__3681));
    LocalMux I__521 (
            .O(N__3686),
            .I(N__3678));
    CascadeMux I__520 (
            .O(N__3685),
            .I(N__3675));
    CascadeMux I__519 (
            .O(N__3684),
            .I(N__3672));
    Span4Mux_v I__518 (
            .O(N__3681),
            .I(N__3669));
    Span4Mux_v I__517 (
            .O(N__3678),
            .I(N__3666));
    InMux I__516 (
            .O(N__3675),
            .I(N__3663));
    InMux I__515 (
            .O(N__3672),
            .I(N__3660));
    Sp12to4 I__514 (
            .O(N__3669),
            .I(N__3650));
    Sp12to4 I__513 (
            .O(N__3666),
            .I(N__3650));
    LocalMux I__512 (
            .O(N__3663),
            .I(N__3650));
    LocalMux I__511 (
            .O(N__3660),
            .I(N__3650));
    InMux I__510 (
            .O(N__3659),
            .I(N__3647));
    Span12Mux_h I__509 (
            .O(N__3650),
            .I(N__3644));
    LocalMux I__508 (
            .O(N__3647),
            .I(N__3641));
    Span12Mux_v I__507 (
            .O(N__3644),
            .I(N__3638));
    Span12Mux_h I__506 (
            .O(N__3641),
            .I(N__3635));
    Odrv12 I__505 (
            .O(N__3638),
            .I(TM_c_0));
    Odrv12 I__504 (
            .O(N__3635),
            .I(TM_c_0));
    InMux I__503 (
            .O(N__3630),
            .I(N__3627));
    LocalMux I__502 (
            .O(N__3627),
            .I(N__3623));
    InMux I__501 (
            .O(N__3626),
            .I(N__3620));
    Span4Mux_v I__500 (
            .O(N__3623),
            .I(N__3615));
    LocalMux I__499 (
            .O(N__3620),
            .I(N__3615));
    Span4Mux_v I__498 (
            .O(N__3615),
            .I(N__3612));
    Odrv4 I__497 (
            .O(N__3612),
            .I(\U409_ADDRESS_DECODE.un2_REGSPACEn_0 ));
    CascadeMux I__496 (
            .O(N__3609),
            .I(N__3602));
    InMux I__495 (
            .O(N__3608),
            .I(N__3599));
    InMux I__494 (
            .O(N__3607),
            .I(N__3596));
    InMux I__493 (
            .O(N__3606),
            .I(N__3588));
    InMux I__492 (
            .O(N__3605),
            .I(N__3588));
    InMux I__491 (
            .O(N__3602),
            .I(N__3588));
    LocalMux I__490 (
            .O(N__3599),
            .I(N__3585));
    LocalMux I__489 (
            .O(N__3596),
            .I(N__3582));
    CascadeMux I__488 (
            .O(N__3595),
            .I(N__3579));
    LocalMux I__487 (
            .O(N__3588),
            .I(N__3576));
    Span4Mux_h I__486 (
            .O(N__3585),
            .I(N__3571));
    Span4Mux_v I__485 (
            .O(N__3582),
            .I(N__3571));
    InMux I__484 (
            .O(N__3579),
            .I(N__3568));
    Span12Mux_h I__483 (
            .O(N__3576),
            .I(N__3565));
    Span4Mux_v I__482 (
            .O(N__3571),
            .I(N__3562));
    LocalMux I__481 (
            .O(N__3568),
            .I(N__3559));
    Odrv12 I__480 (
            .O(N__3565),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    Odrv4 I__479 (
            .O(N__3562),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    Odrv12 I__478 (
            .O(N__3559),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ));
    CascadeMux I__477 (
            .O(N__3552),
            .I(N__3549));
    InMux I__476 (
            .O(N__3549),
            .I(N__3540));
    InMux I__475 (
            .O(N__3548),
            .I(N__3540));
    InMux I__474 (
            .O(N__3547),
            .I(N__3537));
    InMux I__473 (
            .O(N__3546),
            .I(N__3534));
    InMux I__472 (
            .O(N__3545),
            .I(N__3530));
    LocalMux I__471 (
            .O(N__3540),
            .I(N__3525));
    LocalMux I__470 (
            .O(N__3537),
            .I(N__3525));
    LocalMux I__469 (
            .O(N__3534),
            .I(N__3522));
    InMux I__468 (
            .O(N__3533),
            .I(N__3519));
    LocalMux I__467 (
            .O(N__3530),
            .I(N__3516));
    Span4Mux_v I__466 (
            .O(N__3525),
            .I(N__3509));
    Span4Mux_h I__465 (
            .O(N__3522),
            .I(N__3509));
    LocalMux I__464 (
            .O(N__3519),
            .I(N__3509));
    Span4Mux_v I__463 (
            .O(N__3516),
            .I(N__3506));
    Span4Mux_h I__462 (
            .O(N__3509),
            .I(N__3503));
    Sp12to4 I__461 (
            .O(N__3506),
            .I(N__3500));
    Sp12to4 I__460 (
            .O(N__3503),
            .I(N__3497));
    Span12Mux_h I__459 (
            .O(N__3500),
            .I(N__3494));
    Odrv12 I__458 (
            .O(N__3497),
            .I(TM_c_1));
    Odrv12 I__457 (
            .O(N__3494),
            .I(TM_c_1));
    IoInMux I__456 (
            .O(N__3489),
            .I(N__3486));
    LocalMux I__455 (
            .O(N__3486),
            .I(N__3483));
    Span4Mux_s1_v I__454 (
            .O(N__3483),
            .I(N__3480));
    Span4Mux_h I__453 (
            .O(N__3480),
            .I(N__3477));
    Sp12to4 I__452 (
            .O(N__3477),
            .I(N__3474));
    Span12Mux_h I__451 (
            .O(N__3474),
            .I(N__3471));
    Odrv12 I__450 (
            .O(N__3471),
            .I(U409_ADDRESS_DECODE_un1_REGSPACEn_i));
    InMux I__449 (
            .O(N__3468),
            .I(N__3465));
    LocalMux I__448 (
            .O(N__3465),
            .I(\U409_TRANSFER_ACK.N_38 ));
    CascadeMux I__447 (
            .O(N__3462),
            .I(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3Z0Z_2_cascade_ ));
    InMux I__446 (
            .O(N__3459),
            .I(N__3456));
    LocalMux I__445 (
            .O(N__3456),
            .I(N__3451));
    InMux I__444 (
            .O(N__3455),
            .I(N__3448));
    InMux I__443 (
            .O(N__3454),
            .I(N__3445));
    Odrv4 I__442 (
            .O(N__3451),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_6 ));
    LocalMux I__441 (
            .O(N__3448),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_6 ));
    LocalMux I__440 (
            .O(N__3445),
            .I(\U409_ADDRESS_DECODE.CIA_SPACE_6 ));
    CascadeMux I__439 (
            .O(N__3438),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENn_2_cascade_ ));
    CascadeMux I__438 (
            .O(N__3435),
            .I(N__3431));
    CascadeMux I__437 (
            .O(N__3434),
            .I(N__3428));
    InMux I__436 (
            .O(N__3431),
            .I(N__3423));
    InMux I__435 (
            .O(N__3428),
            .I(N__3420));
    InMux I__434 (
            .O(N__3427),
            .I(N__3417));
    InMux I__433 (
            .O(N__3426),
            .I(N__3414));
    LocalMux I__432 (
            .O(N__3423),
            .I(N__3407));
    LocalMux I__431 (
            .O(N__3420),
            .I(N__3407));
    LocalMux I__430 (
            .O(N__3417),
            .I(N__3402));
    LocalMux I__429 (
            .O(N__3414),
            .I(N__3402));
    InMux I__428 (
            .O(N__3413),
            .I(N__3397));
    InMux I__427 (
            .O(N__3412),
            .I(N__3397));
    Span4Mux_v I__426 (
            .O(N__3407),
            .I(N__3393));
    Span4Mux_v I__425 (
            .O(N__3402),
            .I(N__3388));
    LocalMux I__424 (
            .O(N__3397),
            .I(N__3388));
    InMux I__423 (
            .O(N__3396),
            .I(N__3385));
    Sp12to4 I__422 (
            .O(N__3393),
            .I(N__3378));
    Sp12to4 I__421 (
            .O(N__3388),
            .I(N__3378));
    LocalMux I__420 (
            .O(N__3385),
            .I(N__3378));
    Odrv12 I__419 (
            .O(N__3378),
            .I(A_c_20));
    InMux I__418 (
            .O(N__3375),
            .I(N__3372));
    LocalMux I__417 (
            .O(N__3372),
            .I(\U409_ADDRESS_DECODE.REGISTER_SPACEZ0 ));
    CascadeMux I__416 (
            .O(N__3369),
            .I(\U409_ADDRESS_DECODE.RANGER_SPACEZ0Z_2_cascade_ ));
    InMux I__415 (
            .O(N__3366),
            .I(N__3362));
    InMux I__414 (
            .O(N__3365),
            .I(N__3358));
    LocalMux I__413 (
            .O(N__3362),
            .I(N__3353));
    InMux I__412 (
            .O(N__3361),
            .I(N__3350));
    LocalMux I__411 (
            .O(N__3358),
            .I(N__3347));
    InMux I__410 (
            .O(N__3357),
            .I(N__3344));
    InMux I__409 (
            .O(N__3356),
            .I(N__3341));
    Span4Mux_v I__408 (
            .O(N__3353),
            .I(N__3336));
    LocalMux I__407 (
            .O(N__3350),
            .I(N__3336));
    Span4Mux_v I__406 (
            .O(N__3347),
            .I(N__3329));
    LocalMux I__405 (
            .O(N__3344),
            .I(N__3329));
    LocalMux I__404 (
            .O(N__3341),
            .I(N__3329));
    Span4Mux_v I__403 (
            .O(N__3336),
            .I(N__3326));
    Span4Mux_v I__402 (
            .O(N__3329),
            .I(N__3323));
    Sp12to4 I__401 (
            .O(N__3326),
            .I(N__3318));
    Sp12to4 I__400 (
            .O(N__3323),
            .I(N__3318));
    Span12Mux_h I__399 (
            .O(N__3318),
            .I(N__3315));
    Span12Mux_v I__398 (
            .O(N__3315),
            .I(N__3312));
    Odrv12 I__397 (
            .O(N__3312),
            .I(A_c_19));
    CascadeMux I__396 (
            .O(N__3309),
            .I(N__3306));
    InMux I__395 (
            .O(N__3306),
            .I(N__3299));
    InMux I__394 (
            .O(N__3305),
            .I(N__3299));
    InMux I__393 (
            .O(N__3304),
            .I(N__3296));
    LocalMux I__392 (
            .O(N__3299),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ));
    LocalMux I__391 (
            .O(N__3296),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ));
    InMux I__390 (
            .O(N__3291),
            .I(N__3288));
    LocalMux I__389 (
            .O(N__3288),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1 ));
    CascadeMux I__388 (
            .O(N__3285),
            .I(N__3282));
    InMux I__387 (
            .O(N__3282),
            .I(N__3274));
    InMux I__386 (
            .O(N__3281),
            .I(N__3274));
    InMux I__385 (
            .O(N__3280),
            .I(N__3269));
    InMux I__384 (
            .O(N__3279),
            .I(N__3269));
    LocalMux I__383 (
            .O(N__3274),
            .I(N__3264));
    LocalMux I__382 (
            .O(N__3269),
            .I(N__3264));
    Span4Mux_v I__381 (
            .O(N__3264),
            .I(N__3261));
    Span4Mux_v I__380 (
            .O(N__3261),
            .I(N__3258));
    Span4Mux_v I__379 (
            .O(N__3258),
            .I(N__3255));
    Sp12to4 I__378 (
            .O(N__3255),
            .I(N__3252));
    Odrv12 I__377 (
            .O(N__3252),
            .I(A_c_16));
    InMux I__376 (
            .O(N__3249),
            .I(N__3240));
    InMux I__375 (
            .O(N__3248),
            .I(N__3240));
    InMux I__374 (
            .O(N__3247),
            .I(N__3240));
    LocalMux I__373 (
            .O(N__3240),
            .I(N__3237));
    Span4Mux_v I__372 (
            .O(N__3237),
            .I(N__3234));
    Sp12to4 I__371 (
            .O(N__3234),
            .I(N__3231));
    Span12Mux_v I__370 (
            .O(N__3231),
            .I(N__3228));
    Odrv12 I__369 (
            .O(N__3228),
            .I(A_c_17));
    CascadeMux I__368 (
            .O(N__3225),
            .I(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3_cascade_ ));
    CascadeMux I__367 (
            .O(N__3222),
            .I(U409_ADDRESS_DECODE_AUTOVECTOR_5_cascade_));
    CascadeMux I__366 (
            .O(N__3219),
            .I(N__3216));
    InMux I__365 (
            .O(N__3216),
            .I(N__3212));
    InMux I__364 (
            .O(N__3215),
            .I(N__3209));
    LocalMux I__363 (
            .O(N__3212),
            .I(N__3204));
    LocalMux I__362 (
            .O(N__3209),
            .I(N__3204));
    Span4Mux_v I__361 (
            .O(N__3204),
            .I(N__3200));
    InMux I__360 (
            .O(N__3203),
            .I(N__3197));
    Sp12to4 I__359 (
            .O(N__3200),
            .I(N__3192));
    LocalMux I__358 (
            .O(N__3197),
            .I(N__3192));
    Span12Mux_h I__357 (
            .O(N__3192),
            .I(N__3189));
    Span12Mux_v I__356 (
            .O(N__3189),
            .I(N__3186));
    Odrv12 I__355 (
            .O(N__3186),
            .I(A_c_18));
    InMux I__354 (
            .O(N__3183),
            .I(N__3179));
    InMux I__353 (
            .O(N__3182),
            .I(N__3176));
    LocalMux I__352 (
            .O(N__3179),
            .I(N__3173));
    LocalMux I__351 (
            .O(N__3176),
            .I(N__3170));
    Span4Mux_h I__350 (
            .O(N__3173),
            .I(N__3167));
    Span12Mux_h I__349 (
            .O(N__3170),
            .I(N__3164));
    Span4Mux_v I__348 (
            .O(N__3167),
            .I(N__3161));
    Odrv12 I__347 (
            .O(N__3164),
            .I(\U409_ADDRESS_DECODE.AUTOVECTOR_16 ));
    Odrv4 I__346 (
            .O(N__3161),
            .I(\U409_ADDRESS_DECODE.AUTOVECTOR_16 ));
    InMux I__345 (
            .O(N__3156),
            .I(N__3153));
    LocalMux I__344 (
            .O(N__3153),
            .I(N__3150));
    Span4Mux_v I__343 (
            .O(N__3150),
            .I(N__3147));
    Span4Mux_v I__342 (
            .O(N__3147),
            .I(N__3144));
    IoSpan4Mux I__341 (
            .O(N__3144),
            .I(N__3141));
    Odrv4 I__340 (
            .O(N__3141),
            .I(TT_c_1));
    InMux I__339 (
            .O(N__3138),
            .I(N__3135));
    LocalMux I__338 (
            .O(N__3135),
            .I(N__3132));
    Span4Mux_v I__337 (
            .O(N__3132),
            .I(N__3129));
    Span4Mux_v I__336 (
            .O(N__3129),
            .I(N__3126));
    IoSpan4Mux I__335 (
            .O(N__3126),
            .I(N__3123));
    Odrv4 I__334 (
            .O(N__3123),
            .I(TT_c_0));
    InMux I__333 (
            .O(N__3120),
            .I(N__3117));
    LocalMux I__332 (
            .O(N__3117),
            .I(N__3114));
    Odrv12 I__331 (
            .O(N__3114),
            .I(U409_ADDRESS_DECODE_AUTOVECTOR_4));
    InMux I__330 (
            .O(N__3111),
            .I(N__3105));
    InMux I__329 (
            .O(N__3110),
            .I(N__3105));
    LocalMux I__328 (
            .O(N__3105),
            .I(N__3102));
    Span4Mux_v I__327 (
            .O(N__3102),
            .I(N__3099));
    Span4Mux_h I__326 (
            .O(N__3099),
            .I(N__3096));
    Odrv4 I__325 (
            .O(N__3096),
            .I(A_c_31));
    InMux I__324 (
            .O(N__3093),
            .I(N__3087));
    InMux I__323 (
            .O(N__3092),
            .I(N__3087));
    LocalMux I__322 (
            .O(N__3087),
            .I(N__3084));
    Span4Mux_v I__321 (
            .O(N__3084),
            .I(N__3081));
    Sp12to4 I__320 (
            .O(N__3081),
            .I(N__3078));
    Odrv12 I__319 (
            .O(N__3078),
            .I(A_c_30));
    InMux I__318 (
            .O(N__3075),
            .I(N__3072));
    LocalMux I__317 (
            .O(N__3072),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ));
    CascadeMux I__316 (
            .O(N__3069),
            .I(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_ ));
    CascadeMux I__315 (
            .O(N__3066),
            .I(N__3063));
    InMux I__314 (
            .O(N__3063),
            .I(N__3057));
    InMux I__313 (
            .O(N__3062),
            .I(N__3057));
    LocalMux I__312 (
            .O(N__3057),
            .I(N__3054));
    Span4Mux_v I__311 (
            .O(N__3054),
            .I(N__3051));
    Span4Mux_v I__310 (
            .O(N__3051),
            .I(N__3048));
    Sp12to4 I__309 (
            .O(N__3048),
            .I(N__3045));
    Odrv12 I__308 (
            .O(N__3045),
            .I(A_c_26));
    InMux I__307 (
            .O(N__3042),
            .I(N__3036));
    InMux I__306 (
            .O(N__3041),
            .I(N__3036));
    LocalMux I__305 (
            .O(N__3036),
            .I(N__3033));
    Span4Mux_h I__304 (
            .O(N__3033),
            .I(N__3030));
    Span4Mux_v I__303 (
            .O(N__3030),
            .I(N__3027));
    Odrv4 I__302 (
            .O(N__3027),
            .I(A_c_24));
    CascadeMux I__301 (
            .O(N__3024),
            .I(N__3020));
    InMux I__300 (
            .O(N__3023),
            .I(N__3017));
    InMux I__299 (
            .O(N__3020),
            .I(N__3014));
    LocalMux I__298 (
            .O(N__3017),
            .I(N__3009));
    LocalMux I__297 (
            .O(N__3014),
            .I(N__3009));
    Span4Mux_v I__296 (
            .O(N__3009),
            .I(N__3006));
    Sp12to4 I__295 (
            .O(N__3006),
            .I(N__3003));
    Odrv12 I__294 (
            .O(N__3003),
            .I(A_c_27));
    InMux I__293 (
            .O(N__3000),
            .I(N__2994));
    InMux I__292 (
            .O(N__2999),
            .I(N__2994));
    LocalMux I__291 (
            .O(N__2994),
            .I(N__2991));
    Span4Mux_v I__290 (
            .O(N__2991),
            .I(N__2988));
    Span4Mux_h I__289 (
            .O(N__2988),
            .I(N__2985));
    Odrv4 I__288 (
            .O(N__2985),
            .I(A_c_25));
    InMux I__287 (
            .O(N__2982),
            .I(N__2979));
    LocalMux I__286 (
            .O(N__2979),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_3 ));
    InMux I__285 (
            .O(N__2976),
            .I(N__2970));
    InMux I__284 (
            .O(N__2975),
            .I(N__2970));
    LocalMux I__283 (
            .O(N__2970),
            .I(N__2967));
    Span4Mux_h I__282 (
            .O(N__2967),
            .I(N__2964));
    Span4Mux_v I__281 (
            .O(N__2964),
            .I(N__2961));
    Odrv4 I__280 (
            .O(N__2961),
            .I(A_c_29));
    CascadeMux I__279 (
            .O(N__2958),
            .I(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_4_cascade_ ));
    InMux I__278 (
            .O(N__2955),
            .I(N__2949));
    InMux I__277 (
            .O(N__2954),
            .I(N__2949));
    LocalMux I__276 (
            .O(N__2949),
            .I(N__2946));
    Span4Mux_v I__275 (
            .O(N__2946),
            .I(N__2943));
    Span4Mux_v I__274 (
            .O(N__2943),
            .I(N__2940));
    Sp12to4 I__273 (
            .O(N__2940),
            .I(N__2937));
    Odrv12 I__272 (
            .O(N__2937),
            .I(A_c_28));
    IoInMux I__271 (
            .O(N__2934),
            .I(N__2931));
    LocalMux I__270 (
            .O(N__2931),
            .I(N__2928));
    Span12Mux_s11_h I__269 (
            .O(N__2928),
            .I(N__2925));
    Span12Mux_h I__268 (
            .O(N__2925),
            .I(N__2922));
    Odrv12 I__267 (
            .O(N__2922),
            .I(U409_ADDRESS_DECODE_un1_RTC_ENn_i));
    InMux I__266 (
            .O(N__2919),
            .I(N__2916));
    LocalMux I__265 (
            .O(N__2916),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_1 ));
    CascadeMux I__264 (
            .O(N__2913),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_1_cascade_ ));
    InMux I__263 (
            .O(N__2910),
            .I(N__2904));
    InMux I__262 (
            .O(N__2909),
            .I(N__2904));
    LocalMux I__261 (
            .O(N__2904),
            .I(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3 ));
    ClkMux I__260 (
            .O(N__2901),
            .I(N__2868));
    ClkMux I__259 (
            .O(N__2900),
            .I(N__2868));
    ClkMux I__258 (
            .O(N__2899),
            .I(N__2868));
    ClkMux I__257 (
            .O(N__2898),
            .I(N__2868));
    ClkMux I__256 (
            .O(N__2897),
            .I(N__2868));
    ClkMux I__255 (
            .O(N__2896),
            .I(N__2868));
    ClkMux I__254 (
            .O(N__2895),
            .I(N__2868));
    ClkMux I__253 (
            .O(N__2894),
            .I(N__2868));
    ClkMux I__252 (
            .O(N__2893),
            .I(N__2868));
    ClkMux I__251 (
            .O(N__2892),
            .I(N__2868));
    ClkMux I__250 (
            .O(N__2891),
            .I(N__2868));
    GlobalMux I__249 (
            .O(N__2868),
            .I(CLK80_OUT));
    INV \INVU409_TRANSFER_ACK.TACK_EN_iC  (
            .O(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .I(N__2898));
    INV \INVU409_TRANSFER_ACK.TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .I(N__2896));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC_net ),
            .I(N__2894));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .I(N__2892));
    INV \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC  (
            .O(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .I(N__2897));
    INV \INVU409_TRANSFER_ACK.ROM_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .I(N__2895));
    INV \INVU409_TRANSFER_ACK.CIA_ENABLED_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .I(N__2893));
    INV \INVU409_TRANSFER_ACK.CIA_STATE_1C  (
            .O(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .I(N__2891));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .I(N__2901));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .I(N__2899));
    INV \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C  (
            .O(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .I(N__2900));
    defparam IN_MUX_bfv_14_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_4_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_1_0_));
    defparam IN_MUX_bfv_14_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_2_0_ (
            .carryinitin(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .carryinitout(bfn_14_2_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_17_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_17_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_1_17_0  (
            .in0(N__5886),
            .in1(N__3023),
            .in2(N__3066),
            .in3(N__3000),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_3_LC_1_17_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_3_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_3_LC_1_17_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_3_LC_1_17_3  (
            .in0(N__3092),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3110),
            .lcout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_4  (
            .in0(N__3111),
            .in1(N__3042),
            .in2(_gnd_net_),
            .in3(N__3093),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_17_5  (
            .in0(N__3075),
            .in1(N__2976),
            .in2(N__3069),
            .in3(N__2955),
            .lcout(\U409_ADDRESS_DECODE.Z2_SPACEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_4_LC_1_17_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_4_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_4_LC_1_17_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_4_LC_1_17_6  (
            .in0(N__3062),
            .in1(N__3041),
            .in2(N__3024),
            .in3(N__2999),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_LC_1_17_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_LC_1_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_14_LC_1_17_7  (
            .in0(N__2982),
            .in1(N__2975),
            .in2(N__2958),
            .in3(N__2954),
            .lcout(\U409_ADDRESS_DECODE.AUTOVECTOR_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_10_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_10_0 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_5_10_0  (
            .in0(N__3280),
            .in1(N__2910),
            .in2(N__3309),
            .in3(N__2919),
            .lcout(U409_ADDRESS_DECODE_un1_RTC_ENn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_1_LC_5_10_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_1_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_1_LC_5_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_1_LC_5_10_6  (
            .in0(N__3203),
            .in1(N__3898),
            .in2(N__3435),
            .in3(N__3356),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_1 ),
            .ltout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_10_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_10_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_5_10_7  (
            .in0(N__2909),
            .in1(N__3279),
            .in2(N__2913),
            .in3(N__3305),
            .lcout(U409_ADDRESS_DECODE_un1_RTC_ENn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_5_11_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_5_11_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_5_11_0  (
            .in0(N__3607),
            .in1(N__3249),
            .in2(_gnd_net_),
            .in3(N__3807),
            .lcout(\U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_6_LC_5_11_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_6_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_6_LC_5_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_6_LC_5_11_2  (
            .in0(N__3281),
            .in1(N__3806),
            .in2(N__3434),
            .in3(N__3247),
            .lcout(U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_11_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_11_6  (
            .in0(N__3357),
            .in1(N__3215),
            .in2(N__3285),
            .in3(N__3248),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACE_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_5_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_5_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_3_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__3805),
            .in2(_gnd_net_),
            .in3(N__3396),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_5_LC_5_12_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_5_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_5_LC_5_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_5_LC_5_12_4  (
            .in0(N__3454),
            .in1(N__3182),
            .in2(N__3225),
            .in3(N__3964),
            .lcout(),
            .ltout(U409_ADDRESS_DECODE_AUTOVECTOR_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_LC_5_12_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_LC_5_12_5 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_LC_5_12_5  (
            .in0(N__3120),
            .in1(N__4019),
            .in2(N__3222),
            .in3(N__5870),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxaZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_7_LC_5_13_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_7_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_7_LC_5_13_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_7_LC_5_13_1  (
            .in0(N__3365),
            .in1(N__3963),
            .in2(N__3219),
            .in3(N__3183),
            .lcout(U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_5_18_4 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_5_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_5_18_4  (
            .in0(N__3894),
            .in1(N__3156),
            .in2(N__5885),
            .in3(N__3138),
            .lcout(U409_ADDRESS_DECODE_AUTOVECTOR_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_0_LC_6_10_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_0_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_0_LC_6_10_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_0_LC_6_10_0  (
            .in0(N__4083),
            .in1(N__3979),
            .in2(N__3825),
            .in3(N__3899),
            .lcout(\U409_TRANSFER_ACK.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_10_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_10_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_6_10_2  (
            .in0(N__3547),
            .in1(N__3978),
            .in2(_gnd_net_),
            .in3(N__3694),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_2_LC_6_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_2_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_2_LC_6_10_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3_2_LC_6_10_5  (
            .in0(N__3980),
            .in1(N__3427),
            .in2(_gnd_net_),
            .in3(N__3823),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_6_10_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_6_10_6 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_o2_LC_6_10_6  (
            .in0(N__3468),
            .in1(N__3361),
            .in2(N__3462),
            .in3(N__3900),
            .lcout(\U409_TRANSFER_ACK.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_6_11_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_6_11_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_1_LC_6_11_6  (
            .in0(N__3455),
            .in1(N__3819),
            .in2(_gnd_net_),
            .in3(N__3426),
            .lcout(\U409_ADDRESS_DECODE.CIA_SPACEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.REGISTER_SPACE_3_LC_6_12_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.REGISTER_SPACE_3_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.REGISTER_SPACE_3_LC_6_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_ADDRESS_DECODE.REGISTER_SPACE_3_LC_6_12_2  (
            .in0(N__3876),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3413),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.un1_RTC_ENn_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.REGISTER_SPACE_LC_6_12_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.REGISTER_SPACE_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.REGISTER_SPACE_LC_6_12_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.REGISTER_SPACE_LC_6_12_3  (
            .in0(N__3459),
            .in1(N__3817),
            .in2(N__3438),
            .in3(N__3976),
            .lcout(\U409_ADDRESS_DECODE.REGISTER_SPACEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.RANGER_SPACE_2_LC_6_12_5 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.RANGER_SPACE_2_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.RANGER_SPACE_2_LC_6_12_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U409_ADDRESS_DECODE.RANGER_SPACE_2_LC_6_12_5  (
            .in0(N__3412),
            .in1(N__3975),
            .in2(_gnd_net_),
            .in3(N__3816),
            .lcout(),
            .ltout(\U409_ADDRESS_DECODE.RANGER_SPACEZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_LC_6_12_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un2_REGSPACEn_LC_6_12_6 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \U409_ADDRESS_DECODE.un2_REGSPACEn_LC_6_12_6  (
            .in0(N__3877),
            .in1(N__3375),
            .in2(N__3369),
            .in3(N__3366),
            .lcout(\U409_ADDRESS_DECODE.un2_REGSPACEn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_6_13_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_6_13_1 .LUT_INIT=16'b0001001000000000;
    LogicCell40 \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_5_LC_6_13_1  (
            .in0(N__3533),
            .in1(N__3875),
            .in2(N__3684),
            .in3(N__5878),
            .lcout(U409_ADDRESS_DECODE_AUTOCONFIG_SPACE_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_10_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_10_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_10_0  (
            .in0(N__3304),
            .in1(N__3901),
            .in2(N__3609),
            .in3(N__3291),
            .lcout(CIA_SPACE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.ROMEN_1_LC_7_10_3 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.ROMEN_1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.ROMEN_1_LC_7_10_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \U409_ADDRESS_DECODE.ROMEN_1_LC_7_10_3  (
            .in0(N__3695),
            .in1(N__3605),
            .in2(_gnd_net_),
            .in3(N__3548),
            .lcout(U409_ADDRESS_DECODE_ROMEN_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_0_LC_7_10_6 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_0_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_0_LC_7_10_6 .LUT_INIT=16'b0000000000101000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_0_LC_7_10_6  (
            .in0(N__3606),
            .in1(N__3696),
            .in2(N__3552),
            .in3(N__4079),
            .lcout(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0 ),
            .ltout(\U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_7_10_7 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_7_10_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_7_10_7  (
            .in0(N__3902),
            .in1(N__3981),
            .in2(N__4047),
            .in3(N__3824),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_12_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_12_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_7_12_1  (
            .in0(N__4124),
            .in1(N__4023),
            .in2(_gnd_net_),
            .in3(N__4209),
            .lcout(PORTSIZE_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_7_13_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_7_13_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_7_13_0  (
            .in0(N__3977),
            .in1(N__3918),
            .in2(N__3909),
            .in3(N__3818),
            .lcout(U409_ADDRESS_DECODE_un1_RAMSPACEn),
            .ltout(U409_ADDRESS_DECODE_un1_RAMSPACEn_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_7_13_1 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_7_13_1 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_7_13_1  (
            .in0(N__4207),
            .in1(_gnd_net_),
            .in2(N__3750),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(AGNUS_SPACE_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_DATA_BUFFERS.un1_BUFENn_LC_7_13_2 .C_ON=1'b0;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \U409_DATA_BUFFERS.un1_BUFENn_LC_7_13_2 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_DATA_BUFFERS.un1_BUFENn_LC_7_13_2  (
            .in0(N__3747),
            .in1(N__3741),
            .in2(N__3732),
            .in3(N__3729),
            .lcout(BUFENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_8_13_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_8_13_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_8_13_0  (
            .in0(N__3626),
            .in1(N__3608),
            .in2(N__3685),
            .in3(N__3546),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_8_17_0 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_8_17_0 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_8_17_0  (
            .in0(N__3659),
            .in1(N__3630),
            .in2(N__3595),
            .in3(N__3545),
            .lcout(U409_ADDRESS_DECODE_un1_REGSPACEn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_0_LC_9_6_0 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_0_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_0_LC_9_6_0 .LUT_INIT=16'b0000100010000000;
    LogicCell40 \U409_CIA.VMA_RNO_0_LC_9_6_0  (
            .in0(N__4104),
            .in1(N__4275),
            .in2(N__4428),
            .in3(N__4475),
            .lcout(),
            .ltout(\U409_CIA.VMA_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_LC_9_6_1 .C_ON=1'b0;
    defparam \U409_CIA.VMA_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.VMA_LC_9_6_1 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \U409_CIA.VMA_LC_9_6_1  (
            .in0(N__4476),
            .in1(N__4128),
            .in2(N__4107),
            .in3(N__5155),
            .lcout(\U409_CIA.VMAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4584),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNO_1_LC_9_7_1 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNO_1_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNO_1_LC_9_7_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_CIA.VMA_RNO_1_LC_9_7_1  (
            .in0(N__4564),
            .in1(N__4635),
            .in2(N__4506),
            .in3(N__4538),
            .lcout(\U409_CIA.un1_CIA_CLK_COUNT_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_9_8_0 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_9_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__4463),
            .in2(N__4542),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_9_8_1 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_2_LC_9_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_2_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__4631),
            .in2(_gnd_net_),
            .in3(N__4098),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_1 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .clk(N__4583),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_9_8_2 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_9_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__4380),
            .in2(_gnd_net_),
            .in3(N__4095),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_2 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_9_8_3 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_4_LC_9_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_4_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__4415),
            .in2(_gnd_net_),
            .in3(N__4092),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_3 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .clk(N__4583),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_9_8_4 .C_ON=1'b1;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_9_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__4610),
            .in2(_gnd_net_),
            .in3(N__4089),
            .lcout(\U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_4 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_9_8_5 .C_ON=1'b1;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_6_LC_9_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_6_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__4566),
            .in2(_gnd_net_),
            .in3(N__4086),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(\U409_CIA.un2_CIA_CLK_COUNT_cry_5 ),
            .carryout(\U409_CIA.un2_CIA_CLK_COUNT_cry_6 ),
            .clk(N__4583),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_9_8_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_7_LC_9_8_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_7_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__4504),
            .in2(_gnd_net_),
            .in3(N__4227),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4583),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_9_9_6 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_1_LC_9_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_1_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__4541),
            .in2(_gnd_net_),
            .in3(N__4473),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4581),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_11_0 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_11_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_9_11_0  (
            .in0(N__4884),
            .in1(N__4350),
            .in2(_gnd_net_),
            .in3(N__4682),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__4987));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_9_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_9_11_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_9_11_1 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__4217),
            .in2(N__4689),
            .in3(N__4861),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__4987));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_9_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_9_11_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_9_11_6 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_9_11_6  (
            .in0(N__4862),
            .in1(N__4878),
            .in2(N__4221),
            .in3(N__4686),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net ),
            .ce(),
            .sr(N__4987));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIF4AR_5_LC_9_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIF4AR_5_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIF4AR_5_LC_9_12_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIF4AR_5_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__4816),
            .in2(_gnd_net_),
            .in3(N__4348),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_3_LC_9_12_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_3_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_3_LC_9_12_3 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_3_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__4783),
            .in2(N__4224),
            .in3(N__4798),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_1 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_13_1  (
            .in0(N__4208),
            .in1(N__4191),
            .in2(N__5877),
            .in3(N__4182),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_10_4_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_10_4_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_10_4_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_10_4_2  (
            .in0(_gnd_net_),
            .in1(N__4164),
            .in2(_gnd_net_),
            .in3(N__4290),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS1n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_10_5_2 .C_ON=1'b0;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_10_5_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_10_5_2  (
            .in0(N__4286),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4323),
            .lcout(U409_ADDRESS_DECODE_un1_CIACS0n_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.VMA_RNI692L_0_LC_10_6_6 .C_ON=1'b0;
    defparam \U409_CIA.VMA_RNI692L_0_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.VMA_RNI692L_0_LC_10_6_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U409_CIA.VMA_RNI692L_0_LC_10_6_6  (
            .in0(N__5837),
            .in1(N__5156),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CIA_ENABLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNICGRM_3_LC_10_7_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNICGRM_3_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNICGRM_3_LC_10_7_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNICGRM_3_LC_10_7_4  (
            .in0(_gnd_net_),
            .in1(N__4604),
            .in2(_gnd_net_),
            .in3(N__4379),
            .lcout(\U409_CIA.CLK_CIA6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_10_8_0 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_0_LC_10_8_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_0_LC_10_8_0  (
            .in0(N__4274),
            .in1(N__4634),
            .in2(N__4424),
            .in3(N__4437),
            .lcout(),
            .ltout(\U409_CIA.CLK_CIA6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_LC_10_8_1 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CLK_CIA_LC_10_8_1 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \U409_CIA.CLK_CIA_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(N__4903),
            .in2(N__4263),
            .in3(N__4356),
            .lcout(CLK_CIA_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4582),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_10_8_2 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_10_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_3_LC_10_8_2 .LUT_INIT=16'b0001010100101010;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_3_LC_10_8_2  (
            .in0(N__4383),
            .in1(N__4254),
            .in2(N__4239),
            .in3(N__4260),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4582),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_3_LC_10_8_3 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_3_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_3_LC_10_8_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_3_LC_10_8_3  (
            .in0(N__4633),
            .in1(N__4382),
            .in2(N__4611),
            .in3(N__4539),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_2_0 ),
            .ltout(\U409_CIA.CIA_CLK_COUNT11_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_10_8_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_5_LC_10_8_4 .LUT_INIT=16'b0001001101001100;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_5_LC_10_8_4  (
            .in0(N__4238),
            .in1(N__4609),
            .in2(N__4248),
            .in3(N__4245),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4582),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_10_8_5 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_10_8_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_10_8_5  (
            .in0(N__4565),
            .in1(N__4503),
            .in2(N__4474),
            .in3(N__4420),
            .lcout(\U409_CIA.CIA_CLK_COUNT11_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_10_8_6 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_2_LC_10_8_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_2_LC_10_8_6  (
            .in0(_gnd_net_),
            .in1(N__4632),
            .in2(_gnd_net_),
            .in3(N__4605),
            .lcout(\U409_CIA.un1_CIA_CLK_COUNT_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_10_8_7 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_10_8_7 .SEQ_MODE=4'b1000;
    defparam \U409_CIA.CIA_CLK_COUNT_0_LC_10_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_0_LC_10_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4540),
            .lcout(\U409_CIA.CIA_CLK_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4582),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMUMD1_7_LC_10_9_4 .C_ON=1'b0;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMUMD1_7_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CIA_CLK_COUNT_RNIMUMD1_7_LC_10_9_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_CIA.CIA_CLK_COUNT_RNIMUMD1_7_LC_10_9_4  (
            .in0(N__4563),
            .in1(N__4537),
            .in2(N__4505),
            .in3(N__4464),
            .lcout(\U409_CIA.CLK_CIA6_3 ),
            .ltout(\U409_CIA.CLK_CIA6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_10_9_5 .C_ON=1'b0;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U409_CIA.CLK_CIA_RNO_1_LC_10_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_CIA.CLK_CIA_RNO_1_LC_10_9_5  (
            .in0(N__4416),
            .in1(N__4392),
            .in2(N__4386),
            .in3(N__4381),
            .lcout(\U409_CIA.CLK_CIA_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_4 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_10_4  (
            .in0(N__5292),
            .in1(N__4733),
            .in2(_gnd_net_),
            .in3(N__4833),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net ),
            .ce(),
            .sr(N__4995));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_5_LC_10_11_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_5_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_5_LC_10_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_5_LC_10_11_0  (
            .in0(N__4876),
            .in1(N__4823),
            .in2(N__4863),
            .in3(N__4349),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_0_LC_10_11_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_0_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_0_LC_10_11_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_0_LC_10_11_1  (
            .in0(N__4781),
            .in1(N__4716),
            .in2(N__4332),
            .in3(N__4329),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_11_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__4652),
            .in2(_gnd_net_),
            .in3(N__4749),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_11_3 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_11_3  (
            .in0(N__4653),
            .in1(N__4714),
            .in2(N__4758),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3 ),
            .ltout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_10_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_10_11_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(N__4824),
            .in2(N__4887),
            .in3(N__4782),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_11_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_11_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_10_11_5  (
            .in0(N__4654),
            .in1(N__4877),
            .in2(N__4757),
            .in3(N__4857),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_LC_10_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_LC_10_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_LC_10_11_6  (
            .in0(N__4715),
            .in1(N__4780),
            .in2(N__4842),
            .in3(N__4839),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22 ),
            .ltout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_0_LC_10_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_0_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_0_LC_10_11_7 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_0_LC_10_11_7  (
            .in0(N__5523),
            .in1(N__5590),
            .in2(N__4827),
            .in3(N__4732),
            .lcout(\U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_12_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_12_1 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_12_1 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_12_1  (
            .in0(N__4800),
            .in1(N__4785),
            .in2(N__4688),
            .in3(N__4822),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .ce(),
            .sr(N__4994));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_12_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_12_2 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_12_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_12_2  (
            .in0(N__4784),
            .in1(N__4799),
            .in2(_gnd_net_),
            .in3(N__4675),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .ce(),
            .sr(N__4994));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_12_4 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_12_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_12_4  (
            .in0(N__4655),
            .in1(N__4713),
            .in2(_gnd_net_),
            .in3(N__4756),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .ce(),
            .sr(N__4994));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_12_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_12_6 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_12_6 .LUT_INIT=16'b0000000001110011;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_12_6  (
            .in0(N__5583),
            .in1(N__4734),
            .in2(N__5528),
            .in3(N__4711),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .ce(),
            .sr(N__4994));
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_12_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_12_7 .SEQ_MODE=4'b1010;
    defparam \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_12_7 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_12_7  (
            .in0(N__4712),
            .in1(_gnd_net_),
            .in2(N__4687),
            .in3(N__4656),
            .lcout(\U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net ),
            .ce(),
            .sr(N__4994));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_1_LC_11_6_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_1_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_1_LC_11_6_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_1_LC_11_6_0  (
            .in0(N__5490),
            .in1(N__5119),
            .in2(_gnd_net_),
            .in3(N__5099),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.m8_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_LC_11_6_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_LC_11_6_1 .LUT_INIT=16'b0000010100100111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m8_ns_LC_11_6_1  (
            .in0(N__5067),
            .in1(N__4931),
            .in2(N__4962),
            .in3(N__5137),
            .lcout(\U409_TRANSFER_ACK.N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_11_6_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_11_6_2 .LUT_INIT=16'b0000010000110111;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_11_6_2  (
            .in0(N__5138),
            .in1(N__5048),
            .in2(N__4935),
            .in3(N__4950),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.i6_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_6_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_6_3 .LUT_INIT=16'b0010101000001000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_6_3  (
            .in0(N__5822),
            .in1(N__5076),
            .in2(N__4959),
            .in3(N__5050),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_6_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_6_5 .LUT_INIT=16'b0111000000100000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_6_5  (
            .in0(N__5049),
            .in1(N__4956),
            .in2(N__5846),
            .in3(N__4941),
            .lcout(\U409_TRANSFER_ACK.CIA_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_STATE_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_6_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_6_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(N__5118),
            .in2(_gnd_net_),
            .in3(N__5098),
            .lcout(\U409_TRANSFER_ACK.N_4 ),
            .ltout(\U409_TRANSFER_ACK.N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m4_LC_11_6_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m4_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m4_LC_11_6_7 .LUT_INIT=16'b0100111000001010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m4_LC_11_6_7  (
            .in0(N__5068),
            .in1(N__4930),
            .in2(N__4944),
            .in3(N__5136),
            .lcout(\U409_TRANSFER_ACK.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_7_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5139),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(N__5351));
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_11_7_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_0_LC_11_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_0_LC_11_7_1  (
            .in0(N__4904),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(N__5351));
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_11_7_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.LASTCLK_1_LC_11_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.LASTCLK_1_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5121),
            .lcout(\U409_TRANSFER_ACK.LASTCLKZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(N__5351));
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_7_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_7_5  (
            .in0(N__5163),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5838),
            .lcout(\U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net ),
            .ce(),
            .sr(N__5351));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_11_8_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_11_8_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__5682),
            .in2(_gnd_net_),
            .in3(N__5622),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_EN_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_8_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_RNO_0_LC_11_8_6  (
            .in0(N__5051),
            .in1(N__5120),
            .in2(N__5507),
            .in3(N__5100),
            .lcout(\U409_TRANSFER_ACK.N_138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_9_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_9_6 .LUT_INIT=16'b1011111100100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_EN_LC_11_9_6  (
            .in0(N__5436),
            .in1(N__5655),
            .in2(N__5085),
            .in3(N__5279),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(N__5362));
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_9_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_9_7 .LUT_INIT=16'b0100011101000000;
    LogicCell40 \U409_TRANSFER_ACK.CIA_TACK_EN_LC_11_9_7  (
            .in0(N__5075),
            .in1(N__5052),
            .in2(N__5022),
            .in3(N__5265),
            .lcout(\U409_TRANSFER_ACK.CIA_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_ENC_net ),
            .ce(),
            .sr(N__5362));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_11_10_1 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_11_10_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_11_10_1  (
            .in0(N__5012),
            .in1(N__5495),
            .in2(N__5591),
            .in3(N__5393),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNIG3KDC_LC_11_10_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNIG3KDC_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNIG3KDC_LC_11_10_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNIG3KDC_LC_11_10_3  (
            .in0(N__5013),
            .in1(N__5494),
            .in2(N__5592),
            .in3(N__5392),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNO_LC_11_10_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNO_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNO_LC_11_10_4 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNO_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5295),
            .in3(N__5363),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNIECRR_LC_11_10_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNIECRR_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNIECRR_LC_11_10_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_RNIECRR_LC_11_10_7  (
            .in0(N__5379),
            .in1(N__5291),
            .in2(N__5280),
            .in3(N__5264),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTER6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_7_0.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_7_0.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_7_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_7_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5788),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_12_7_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_12_7_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_12_7_2  (
            .in0(N__5677),
            .in1(N__5619),
            .in2(_gnd_net_),
            .in3(N__5649),
            .lcout(\U409_TRANSFER_ACK.N_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_7_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_7_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_7_4  (
            .in0(N__5621),
            .in1(N__5430),
            .in2(N__5689),
            .in3(N__5650),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_7_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_7_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_12_7_6  (
            .in0(N__5681),
            .in1(N__5620),
            .in2(N__5238),
            .in3(N__5651),
            .lcout(\U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_8_0 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_8_0 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_8_0  (
            .in0(N__5403),
            .in1(N__5435),
            .in2(N__5237),
            .in3(N__5211),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5358));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_12_8_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_12_8_2 .LUT_INIT=16'b0111100010110000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_12_8_2  (
            .in0(N__5625),
            .in1(N__5434),
            .in2(N__5691),
            .in3(N__5654),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5358));
    defparam \U409_TRANSFER_ACK.ROMENn_LC_12_8_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_12_8_3 .SEQ_MODE=4'b1001;
    defparam \U409_TRANSFER_ACK.ROMENn_LC_12_8_3 .LUT_INIT=16'b1111111101110000;
    LogicCell40 \U409_TRANSFER_ACK.ROMENn_LC_12_8_3  (
            .in0(N__5205),
            .in1(N__5402),
            .in2(N__5180),
            .in3(N__5199),
            .lcout(ROMENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5358));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_8_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_8_4 .LUT_INIT=16'b0011001110001100;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_8_4  (
            .in0(N__5623),
            .in1(N__5432),
            .in2(N__5690),
            .in3(N__5652),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5358));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_8_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_8_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_8_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_8_6  (
            .in0(N__5624),
            .in1(N__5433),
            .in2(_gnd_net_),
            .in3(N__5653),
            .lcout(\U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net ),
            .ce(),
            .sr(N__5358));
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIPTM34_0_LC_12_9_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIPTM34_0_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIPTM34_0_LC_12_9_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIPTM34_0_LC_12_9_2  (
            .in0(N__5571),
            .in1(N__5541),
            .in2(N__5524),
            .in3(N__5431),
            .lcout(\U409_TRANSFER_ACK.N_28_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_LC_12_10_5 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_LC_12_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U409_TRANSFER_ACK.IRQ_TACK_EN_nesr_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5394),
            .lcout(\U409_TRANSFER_ACK.IRQ_TACK_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.IRQ_TACK_EN_nesrC_net ),
            .ce(N__5373),
            .sr(N__5364));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_11_2 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_11_2 .LUT_INIT=16'b0000000011010000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_11_2  (
            .in0(N__5723),
            .in1(N__5931),
            .in2(N__5847),
            .in3(N__5906),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_12_11_3 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_12_11_3 .LUT_INIT=16'b0010001100100111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_12_11_3  (
            .in0(N__5903),
            .in1(N__5308),
            .in2(N__5933),
            .in3(N__5721),
            .lcout(),
            .ltout(\U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_12_11_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_12_11_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_OUTn_LC_12_11_4 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \U409_TRANSFER_ACK.TACK_OUTn_LC_12_11_4  (
            .in0(N__5309),
            .in1(_gnd_net_),
            .in2(N__5322),
            .in3(N__5828),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_11_6 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_11_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_11_6  (
            .in0(N__5826),
            .in1(N__5930),
            .in2(_gnd_net_),
            .in3(N__5905),
            .lcout(\U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_12_11_7 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_12_11_7 .LUT_INIT=16'b1011001110110111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_12_11_7  (
            .in0(N__5904),
            .in1(N__5827),
            .in2(N__5934),
            .in3(N__5722),
            .lcout(\U409_TRANSFER_ACK.TACK_OUTn_0_sqmuxa_0_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_12_12_4 .C_ON=1'b0;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \U409_TRANSFER_ACK.TACK_EN_i_LC_12_12_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \U409_TRANSFER_ACK.TACK_EN_i_LC_12_12_4  (
            .in0(N__5932),
            .in1(N__5907),
            .in2(N__5848),
            .in3(N__5727),
            .lcout(TACK_EN_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU409_TRANSFER_ACK.TACK_EN_iC_net ),
            .ce(N__5706),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_8_LC_13_3_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_8_LC_13_3_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_8_LC_13_3_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_8_LC_13_3_4  (
            .in0(N__6008),
            .in1(N__6039),
            .in2(N__5976),
            .in3(N__6294),
            .lcout(\U409_TICK.COUNTER60Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6770),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_4_LC_13_4_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_4_LC_13_4_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_4_LC_13_4_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_4_LC_13_4_0  (
            .in0(N__5965),
            .in1(N__6035),
            .in2(N__6114),
            .in3(N__6001),
            .lcout(\U409_TICK.COUNTER60Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6773),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_6_LC_13_4_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_6_LC_13_4_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_6_LC_13_4_1 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_6_LC_13_4_1  (
            .in0(N__6033),
            .in1(N__5966),
            .in2(N__6009),
            .in3(N__6336),
            .lcout(\U409_TICK.COUNTER60Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6773),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_4_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_4_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_4_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U409_TICK.COUNTER60_RNIHJU51_4_LC_13_4_2  (
            .in0(N__6363),
            .in1(N__6126),
            .in2(_gnd_net_),
            .in3(N__6174),
            .lcout(),
            .ltout(\U409_TICK.TICK603_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_4_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_4_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI335G2_11_LC_13_4_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI335G2_11_LC_13_4_3  (
            .in0(N__6246),
            .in1(N__6045),
            .in2(N__5697),
            .in3(N__6141),
            .lcout(\U409_TICK.TICK603_14 ),
            .ltout(\U409_TICK.TICK603_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_0_LC_13_4_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_0_LC_13_4_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_0_LC_13_4_4 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER60_0_LC_13_4_4  (
            .in0(N__5964),
            .in1(N__6000),
            .in2(N__5694),
            .in3(N__6175),
            .lcout(\U409_TICK.COUNTER60Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6773),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_1_LC_13_4_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_1_LC_13_4_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_1_LC_13_4_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER60_1_LC_13_4_5  (
            .in0(N__6176),
            .in1(_gnd_net_),
            .in2(N__6201),
            .in3(_gnd_net_),
            .lcout(\U409_TICK.COUNTER60Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6773),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_13_4_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_13_4_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNICDC71_14_LC_13_4_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER60_RNICDC71_14_LC_13_4_6  (
            .in0(N__6285),
            .in1(N__6486),
            .in2(N__6309),
            .in3(N__6348),
            .lcout(\U409_TICK.TICK603_9 ),
            .ltout(\U409_TICK.TICK603_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK60_LC_13_4_7 .C_ON=1'b0;
    defparam \U409_TICK.TICK60_LC_13_4_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK60_LC_13_4_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK60_LC_13_4_7  (
            .in0(N__6034),
            .in1(N__6059),
            .in2(N__6075),
            .in3(N__5967),
            .lcout(TICK60_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6773),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_9_LC_13_5_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_9_LC_13_5_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_9_LC_13_5_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER60_9_LC_13_5_0  (
            .in0(N__6007),
            .in1(N__5968),
            .in2(N__6273),
            .in3(N__6038),
            .lcout(\U409_TICK.COUNTER60Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6775),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_5_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNI2USG_10_LC_13_5_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U409_TICK.COUNTER60_RNI2USG_10_LC_13_5_1  (
            .in0(N__6501),
            .in1(N__6261),
            .in2(N__6327),
            .in3(N__6465),
            .lcout(\U409_TICK.TICK603_10 ),
            .ltout(\U409_TICK.TICK603_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_14_LC_13_5_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_14_LC_13_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_14_LC_13_5_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_14_LC_13_5_2  (
            .in0(N__6005),
            .in1(N__6037),
            .in2(N__6048),
            .in3(N__6474),
            .lcout(\U409_TICK.COUNTER60Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6775),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_5_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_5_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER60_RNIDB4S_16_LC_13_5_5  (
            .in0(N__6231),
            .in1(N__6156),
            .in2(N__6200),
            .in3(N__6440),
            .lcout(\U409_TICK.TICK603_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_15_LC_13_5_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_15_LC_13_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_15_LC_13_5_7 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER60_15_LC_13_5_7  (
            .in0(N__6036),
            .in1(N__6006),
            .in2(N__5975),
            .in3(N__6453),
            .lcout(\U409_TICK.COUNTER60Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6775),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_1_0 .C_ON=1'b1;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_1_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_1_0  (
            .in0(_gnd_net_),
            .in1(N__6655),
            .in2(N__6411),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_1_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_2_LC_14_1_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_2_LC_14_1_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_2_LC_14_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_2_LC_14_1_1  (
            .in0(_gnd_net_),
            .in1(N__6674),
            .in2(_gnd_net_),
            .in3(N__5937),
            .lcout(\U409_TICK.COUNTER50Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_1 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .clk(N__6769),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_3_LC_14_1_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_3_LC_14_1_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_3_LC_14_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_3_LC_14_1_2  (
            .in0(_gnd_net_),
            .in1(N__6422),
            .in2(_gnd_net_),
            .in3(N__6102),
            .lcout(\U409_TICK.COUNTER50Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_2 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .clk(N__6769),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_4_LC_14_1_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_4_LC_14_1_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_4_LC_14_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_4_LC_14_1_3  (
            .in0(_gnd_net_),
            .in1(N__6533),
            .in2(_gnd_net_),
            .in3(N__6099),
            .lcout(\U409_TICK.COUNTER50Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_3 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .clk(N__6769),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_1_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_1_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_5_LC_14_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_5_LC_14_1_4  (
            .in0(_gnd_net_),
            .in1(N__6698),
            .in2(_gnd_net_),
            .in3(N__6096),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_4 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_1_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_1_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_6_LC_14_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_6_LC_14_1_5  (
            .in0(_gnd_net_),
            .in1(N__6578),
            .in2(_gnd_net_),
            .in3(N__6093),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_5 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_7_LC_14_1_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_7_LC_14_1_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_7_LC_14_1_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_7_LC_14_1_6  (
            .in0(_gnd_net_),
            .in1(N__6545),
            .in2(_gnd_net_),
            .in3(N__6090),
            .lcout(\U409_TICK.COUNTER50Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_6 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .clk(N__6769),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_8_LC_14_1_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_8_LC_14_1_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_8_LC_14_1_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_8_LC_14_1_7  (
            .in0(_gnd_net_),
            .in1(N__6686),
            .in2(_gnd_net_),
            .in3(N__6087),
            .lcout(\U409_TICK.COUNTER50Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_7 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_8 ),
            .clk(N__6769),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_2_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_2_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_9_LC_14_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_9_LC_14_2_0  (
            .in0(_gnd_net_),
            .in1(N__6593),
            .in2(_gnd_net_),
            .in3(N__6084),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_14_2_0_),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_10_LC_14_2_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_10_LC_14_2_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_10_LC_14_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_10_LC_14_2_1  (
            .in0(_gnd_net_),
            .in1(N__6374),
            .in2(_gnd_net_),
            .in3(N__6081),
            .lcout(\U409_TICK.COUNTER50Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_9 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .clk(N__6771),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_2_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_2_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_11_LC_14_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_11_LC_14_2_2  (
            .in0(_gnd_net_),
            .in1(N__6512),
            .in2(_gnd_net_),
            .in3(N__6078),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_10 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_12_LC_14_2_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_12_LC_14_2_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_12_LC_14_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_12_LC_14_2_3  (
            .in0(_gnd_net_),
            .in1(N__6389),
            .in2(_gnd_net_),
            .in3(N__6216),
            .lcout(\U409_TICK.COUNTER50Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_11 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .clk(N__6771),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_2_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_2_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_13_LC_14_2_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_13_LC_14_2_4  (
            .in0(_gnd_net_),
            .in1(N__6557),
            .in2(_gnd_net_),
            .in3(N__6213),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_12 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_2_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_2_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_14_LC_14_2_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_14_LC_14_2_5  (
            .in0(_gnd_net_),
            .in1(N__6788),
            .in2(_gnd_net_),
            .in3(N__6210),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_13 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_2_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_2_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNO_0_15_LC_14_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER50_RNO_0_15_LC_14_2_6  (
            .in0(_gnd_net_),
            .in1(N__6923),
            .in2(_gnd_net_),
            .in3(N__6207),
            .lcout(\U409_TICK.COUNTER50_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un2_COUNTER50_1_cry_14 ),
            .carryout(\U409_TICK.un2_COUNTER50_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_16_LC_14_2_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_16_LC_14_2_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_16_LC_14_2_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER50_16_LC_14_2_7  (
            .in0(_gnd_net_),
            .in1(N__6642),
            .in2(_gnd_net_),
            .in3(N__6204),
            .lcout(\U409_TICK.COUNTER50Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6771),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_4_0 .C_ON=1'b1;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_4_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_4_0  (
            .in0(_gnd_net_),
            .in1(N__6193),
            .in2(N__6177),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_4_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_2_LC_14_4_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_2_LC_14_4_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_2_LC_14_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_2_LC_14_4_1  (
            .in0(_gnd_net_),
            .in1(N__6155),
            .in2(_gnd_net_),
            .in3(N__6144),
            .lcout(\U409_TICK.COUNTER60Z0Z_2 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_1 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .clk(N__6776),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_3_LC_14_4_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_3_LC_14_4_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_3_LC_14_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_3_LC_14_4_2  (
            .in0(_gnd_net_),
            .in1(N__6140),
            .in2(_gnd_net_),
            .in3(N__6129),
            .lcout(\U409_TICK.COUNTER60Z0Z_3 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_2 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .clk(N__6776),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_14_4_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_14_4_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_4_LC_14_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_4_LC_14_4_3  (
            .in0(_gnd_net_),
            .in1(N__6125),
            .in2(_gnd_net_),
            .in3(N__6105),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_3 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_5_LC_14_4_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_5_LC_14_4_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_5_LC_14_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_5_LC_14_4_4  (
            .in0(_gnd_net_),
            .in1(N__6362),
            .in2(_gnd_net_),
            .in3(N__6351),
            .lcout(\U409_TICK.COUNTER60Z0Z_5 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_4 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .clk(N__6776),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_14_4_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_14_4_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_6_LC_14_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_6_LC_14_4_5  (
            .in0(_gnd_net_),
            .in1(N__6347),
            .in2(_gnd_net_),
            .in3(N__6330),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_5 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_7_LC_14_4_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_7_LC_14_4_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_7_LC_14_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_7_LC_14_4_6  (
            .in0(_gnd_net_),
            .in1(N__6323),
            .in2(_gnd_net_),
            .in3(N__6312),
            .lcout(\U409_TICK.COUNTER60Z0Z_7 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_6 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .clk(N__6776),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_14_4_7 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_14_4_7 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_8_LC_14_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_8_LC_14_4_7  (
            .in0(_gnd_net_),
            .in1(N__6305),
            .in2(_gnd_net_),
            .in3(N__6288),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_7 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_14_5_0 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_9_LC_14_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_9_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(N__6284),
            .in2(_gnd_net_),
            .in3(N__6264),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_10_LC_14_5_1 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_10_LC_14_5_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_10_LC_14_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_10_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(N__6260),
            .in2(_gnd_net_),
            .in3(N__6249),
            .lcout(\U409_TICK.COUNTER60Z0Z_10 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_9 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .clk(N__6777),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_11_LC_14_5_2 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_11_LC_14_5_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_11_LC_14_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_11_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(N__6245),
            .in2(_gnd_net_),
            .in3(N__6234),
            .lcout(\U409_TICK.COUNTER60Z0Z_11 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_10 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .clk(N__6777),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_12_LC_14_5_3 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_12_LC_14_5_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_12_LC_14_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_12_LC_14_5_3  (
            .in0(_gnd_net_),
            .in1(N__6230),
            .in2(_gnd_net_),
            .in3(N__6219),
            .lcout(\U409_TICK.COUNTER60Z0Z_12 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_11 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .clk(N__6777),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_13_LC_14_5_4 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_13_LC_14_5_4 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_13_LC_14_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_13_LC_14_5_4  (
            .in0(_gnd_net_),
            .in1(N__6500),
            .in2(_gnd_net_),
            .in3(N__6489),
            .lcout(\U409_TICK.COUNTER60Z0Z_13 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_12 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .clk(N__6777),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_14_5_5 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_14_LC_14_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_14_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(N__6485),
            .in2(_gnd_net_),
            .in3(N__6468),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_13 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_14_5_6 .C_ON=1'b1;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER60_RNO_0_15_LC_14_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U409_TICK.COUNTER60_RNO_0_15_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(N__6464),
            .in2(_gnd_net_),
            .in3(N__6447),
            .lcout(\U409_TICK.COUNTER60_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\U409_TICK.un3_COUNTER60_1_cry_14 ),
            .carryout(\U409_TICK.un3_COUNTER60_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER60_16_LC_14_5_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER60_16_LC_14_5_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER60_16_LC_14_5_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U409_TICK.COUNTER60_16_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(N__6441),
            .in2(_gnd_net_),
            .in3(N__6444),
            .lcout(\U409_TICK.COUNTER60Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6777),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_6_LC_15_1_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_6_LC_15_1_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_6_LC_15_1_0 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_6_LC_15_1_0  (
            .in0(N__6906),
            .in1(N__6881),
            .in2(N__6843),
            .in3(N__6429),
            .lcout(\U409_TICK.COUNTER50Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6772),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_0_LC_15_1_1 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_0_LC_15_1_1 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_0_LC_15_1_1 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \U409_TICK.COUNTER50_0_LC_15_1_1  (
            .in0(N__6879),
            .in1(N__6905),
            .in2(N__6837),
            .in3(N__6409),
            .lcout(\U409_TICK.COUNTER50Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6772),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_1_LC_15_1_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_1_LC_15_1_2 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_1_LC_15_1_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \U409_TICK.COUNTER50_1_LC_15_1_2  (
            .in0(N__6410),
            .in1(_gnd_net_),
            .in2(N__6663),
            .in3(_gnd_net_),
            .lcout(\U409_TICK.COUNTER50Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6772),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_15_1_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_15_1_3 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNID6CP_3_LC_15_1_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U409_TICK.COUNTER50_RNID6CP_3_LC_15_1_3  (
            .in0(N__6699),
            .in1(N__6423),
            .in2(_gnd_net_),
            .in3(N__6408),
            .lcout(),
            .ltout(\U409_TICK.TICK503_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_15_1_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_15_1_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNITU182_10_LC_15_1_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNITU182_10_LC_15_1_4  (
            .in0(N__6630),
            .in1(N__6390),
            .in2(N__6378),
            .in3(N__6375),
            .lcout(\U409_TICK.TICK503_14 ),
            .ltout(\U409_TICK.TICK503_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_5_LC_15_1_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_5_LC_15_1_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_5_LC_15_1_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_5_LC_15_1_5  (
            .in0(N__6880),
            .in1(N__6839),
            .in2(N__6708),
            .in3(N__6705),
            .lcout(\U409_TICK.COUNTER50Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6772),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_15_1_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_15_1_6 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIUHF01_16_LC_15_1_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U409_TICK.COUNTER50_RNIUHF01_16_LC_15_1_6  (
            .in0(N__6687),
            .in1(N__6675),
            .in2(N__6662),
            .in3(N__6641),
            .lcout(\U409_TICK.TICK503_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.TICK50_LC_15_1_7 .C_ON=1'b0;
    defparam \U409_TICK.TICK50_LC_15_1_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.TICK50_LC_15_1_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \U409_TICK.TICK50_LC_15_1_7  (
            .in0(N__6882),
            .in1(N__6614),
            .in2(N__6838),
            .in3(N__6907),
            .lcout(TICK50_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6772),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_9_LC_15_2_0 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_9_LC_15_2_0 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_9_LC_15_2_0 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \U409_TICK.COUNTER50_9_LC_15_2_0  (
            .in0(N__6878),
            .in1(N__6603),
            .in2(N__6836),
            .in3(N__6912),
            .lcout(\U409_TICK.COUNTER50Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6774),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_15_2_2 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_15_2_2 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNIH14V_11_LC_15_2_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U409_TICK.COUNTER50_RNIH14V_11_LC_15_2_2  (
            .in0(N__6513),
            .in1(N__6594),
            .in2(N__6582),
            .in3(N__6558),
            .lcout(\U409_TICK.TICK503_9 ),
            .ltout(\U409_TICK.TICK503_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_13_LC_15_2_3 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_13_LC_15_2_3 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_13_LC_15_2_3 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_13_LC_15_2_3  (
            .in0(N__6909),
            .in1(N__6875),
            .in2(N__6567),
            .in3(N__6564),
            .lcout(\U409_TICK.COUNTER50Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6774),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_15_2_4 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_15_2_4 .SEQ_MODE=4'b0000;
    defparam \U409_TICK.COUNTER50_RNII24V_14_LC_15_2_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U409_TICK.COUNTER50_RNII24V_14_LC_15_2_4  (
            .in0(N__6924),
            .in1(N__6546),
            .in2(N__6792),
            .in3(N__6534),
            .lcout(\U409_TICK.TICK503_10 ),
            .ltout(\U409_TICK.TICK503_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_11_LC_15_2_5 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_11_LC_15_2_5 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_11_LC_15_2_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_11_LC_15_2_5  (
            .in0(N__6908),
            .in1(N__6819),
            .in2(N__6522),
            .in3(N__6519),
            .lcout(\U409_TICK.COUNTER50Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6774),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_15_LC_15_2_6 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_15_LC_15_2_6 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_15_LC_15_2_6 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \U409_TICK.COUNTER50_15_LC_15_2_6  (
            .in0(N__6877),
            .in1(N__6911),
            .in2(N__6835),
            .in3(N__6930),
            .lcout(\U409_TICK.COUNTER50Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6774),
            .ce(),
            .sr(_gnd_net_));
    defparam \U409_TICK.COUNTER50_14_LC_15_2_7 .C_ON=1'b0;
    defparam \U409_TICK.COUNTER50_14_LC_15_2_7 .SEQ_MODE=4'b1000;
    defparam \U409_TICK.COUNTER50_14_LC_15_2_7 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \U409_TICK.COUNTER50_14_LC_15_2_7  (
            .in0(N__6910),
            .in1(N__6876),
            .in2(N__6852),
            .in3(N__6820),
            .lcout(\U409_TICK.COUNTER50Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__6774),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_iobuf_RNO_LC_19_18_5.C_ON=1'b0;
    defparam TACKn_iobuf_RNO_LC_19_18_5.SEQ_MODE=4'b0000;
    defparam TACKn_iobuf_RNO_LC_19_18_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_iobuf_RNO_LC_19_18_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6744),
            .lcout(N_475_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U409_TOP

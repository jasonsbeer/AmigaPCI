// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 25 2025 20:17:12

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    CMA,
    DRA,
    SIZ,
    A,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    DBRn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    output [10:0] CMA;
    input [9:0] DRA;
    input [1:0] SIZ;
    input [20:0] A;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input DBRn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__12003;
    wire N__12002;
    wire N__12001;
    wire N__11994;
    wire N__11993;
    wire N__11992;
    wire N__11985;
    wire N__11984;
    wire N__11983;
    wire N__11976;
    wire N__11975;
    wire N__11974;
    wire N__11967;
    wire N__11966;
    wire N__11965;
    wire N__11958;
    wire N__11957;
    wire N__11956;
    wire N__11949;
    wire N__11948;
    wire N__11947;
    wire N__11940;
    wire N__11939;
    wire N__11938;
    wire N__11931;
    wire N__11930;
    wire N__11929;
    wire N__11922;
    wire N__11921;
    wire N__11920;
    wire N__11913;
    wire N__11912;
    wire N__11911;
    wire N__11904;
    wire N__11903;
    wire N__11902;
    wire N__11895;
    wire N__11894;
    wire N__11893;
    wire N__11886;
    wire N__11885;
    wire N__11884;
    wire N__11877;
    wire N__11876;
    wire N__11875;
    wire N__11868;
    wire N__11867;
    wire N__11866;
    wire N__11859;
    wire N__11858;
    wire N__11857;
    wire N__11850;
    wire N__11849;
    wire N__11848;
    wire N__11841;
    wire N__11840;
    wire N__11839;
    wire N__11832;
    wire N__11831;
    wire N__11830;
    wire N__11823;
    wire N__11822;
    wire N__11821;
    wire N__11814;
    wire N__11813;
    wire N__11812;
    wire N__11805;
    wire N__11804;
    wire N__11803;
    wire N__11796;
    wire N__11795;
    wire N__11794;
    wire N__11787;
    wire N__11786;
    wire N__11785;
    wire N__11778;
    wire N__11777;
    wire N__11776;
    wire N__11769;
    wire N__11768;
    wire N__11767;
    wire N__11760;
    wire N__11759;
    wire N__11758;
    wire N__11751;
    wire N__11750;
    wire N__11749;
    wire N__11742;
    wire N__11741;
    wire N__11740;
    wire N__11733;
    wire N__11732;
    wire N__11731;
    wire N__11724;
    wire N__11723;
    wire N__11722;
    wire N__11715;
    wire N__11714;
    wire N__11713;
    wire N__11706;
    wire N__11705;
    wire N__11704;
    wire N__11697;
    wire N__11696;
    wire N__11695;
    wire N__11688;
    wire N__11687;
    wire N__11686;
    wire N__11679;
    wire N__11678;
    wire N__11677;
    wire N__11670;
    wire N__11669;
    wire N__11668;
    wire N__11661;
    wire N__11660;
    wire N__11659;
    wire N__11652;
    wire N__11651;
    wire N__11650;
    wire N__11643;
    wire N__11642;
    wire N__11641;
    wire N__11634;
    wire N__11633;
    wire N__11632;
    wire N__11625;
    wire N__11624;
    wire N__11623;
    wire N__11616;
    wire N__11615;
    wire N__11614;
    wire N__11607;
    wire N__11606;
    wire N__11605;
    wire N__11598;
    wire N__11597;
    wire N__11596;
    wire N__11589;
    wire N__11588;
    wire N__11587;
    wire N__11580;
    wire N__11579;
    wire N__11578;
    wire N__11571;
    wire N__11570;
    wire N__11569;
    wire N__11562;
    wire N__11561;
    wire N__11560;
    wire N__11553;
    wire N__11552;
    wire N__11551;
    wire N__11544;
    wire N__11543;
    wire N__11542;
    wire N__11535;
    wire N__11534;
    wire N__11533;
    wire N__11526;
    wire N__11525;
    wire N__11524;
    wire N__11517;
    wire N__11516;
    wire N__11515;
    wire N__11508;
    wire N__11507;
    wire N__11506;
    wire N__11499;
    wire N__11498;
    wire N__11497;
    wire N__11490;
    wire N__11489;
    wire N__11488;
    wire N__11481;
    wire N__11480;
    wire N__11479;
    wire N__11472;
    wire N__11471;
    wire N__11470;
    wire N__11463;
    wire N__11462;
    wire N__11461;
    wire N__11454;
    wire N__11453;
    wire N__11452;
    wire N__11445;
    wire N__11444;
    wire N__11443;
    wire N__11436;
    wire N__11435;
    wire N__11434;
    wire N__11427;
    wire N__11426;
    wire N__11425;
    wire N__11418;
    wire N__11417;
    wire N__11416;
    wire N__11409;
    wire N__11408;
    wire N__11407;
    wire N__11400;
    wire N__11399;
    wire N__11398;
    wire N__11391;
    wire N__11390;
    wire N__11389;
    wire N__11382;
    wire N__11381;
    wire N__11380;
    wire N__11373;
    wire N__11372;
    wire N__11371;
    wire N__11364;
    wire N__11363;
    wire N__11362;
    wire N__11355;
    wire N__11354;
    wire N__11353;
    wire N__11346;
    wire N__11345;
    wire N__11344;
    wire N__11337;
    wire N__11336;
    wire N__11335;
    wire N__11328;
    wire N__11327;
    wire N__11326;
    wire N__11319;
    wire N__11318;
    wire N__11317;
    wire N__11310;
    wire N__11309;
    wire N__11308;
    wire N__11301;
    wire N__11300;
    wire N__11299;
    wire N__11292;
    wire N__11291;
    wire N__11290;
    wire N__11283;
    wire N__11282;
    wire N__11281;
    wire N__11274;
    wire N__11273;
    wire N__11272;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11256;
    wire N__11255;
    wire N__11254;
    wire N__11247;
    wire N__11246;
    wire N__11245;
    wire N__11238;
    wire N__11237;
    wire N__11236;
    wire N__11229;
    wire N__11228;
    wire N__11227;
    wire N__11220;
    wire N__11219;
    wire N__11218;
    wire N__11211;
    wire N__11210;
    wire N__11209;
    wire N__11192;
    wire N__11189;
    wire N__11188;
    wire N__11185;
    wire N__11184;
    wire N__11183;
    wire N__11182;
    wire N__11181;
    wire N__11178;
    wire N__11177;
    wire N__11174;
    wire N__11169;
    wire N__11164;
    wire N__11163;
    wire N__11158;
    wire N__11157;
    wire N__11156;
    wire N__11155;
    wire N__11154;
    wire N__11153;
    wire N__11152;
    wire N__11151;
    wire N__11150;
    wire N__11147;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11113;
    wire N__11112;
    wire N__11105;
    wire N__11100;
    wire N__11099;
    wire N__11088;
    wire N__11087;
    wire N__11084;
    wire N__11083;
    wire N__11080;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11048;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11026;
    wire N__11021;
    wire N__11020;
    wire N__11017;
    wire N__11014;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__11000;
    wire N__10997;
    wire N__10996;
    wire N__10995;
    wire N__10992;
    wire N__10991;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10963;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10942;
    wire N__10941;
    wire N__10940;
    wire N__10939;
    wire N__10938;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10918;
    wire N__10917;
    wire N__10916;
    wire N__10915;
    wire N__10914;
    wire N__10913;
    wire N__10912;
    wire N__10911;
    wire N__10910;
    wire N__10909;
    wire N__10908;
    wire N__10907;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10873;
    wire N__10872;
    wire N__10871;
    wire N__10870;
    wire N__10867;
    wire N__10864;
    wire N__10861;
    wire N__10858;
    wire N__10855;
    wire N__10854;
    wire N__10853;
    wire N__10852;
    wire N__10851;
    wire N__10850;
    wire N__10849;
    wire N__10848;
    wire N__10847;
    wire N__10846;
    wire N__10845;
    wire N__10844;
    wire N__10841;
    wire N__10840;
    wire N__10839;
    wire N__10838;
    wire N__10837;
    wire N__10836;
    wire N__10833;
    wire N__10832;
    wire N__10831;
    wire N__10830;
    wire N__10829;
    wire N__10828;
    wire N__10825;
    wire N__10824;
    wire N__10823;
    wire N__10822;
    wire N__10821;
    wire N__10820;
    wire N__10819;
    wire N__10816;
    wire N__10815;
    wire N__10814;
    wire N__10813;
    wire N__10812;
    wire N__10811;
    wire N__10810;
    wire N__10809;
    wire N__10808;
    wire N__10807;
    wire N__10806;
    wire N__10803;
    wire N__10802;
    wire N__10801;
    wire N__10800;
    wire N__10799;
    wire N__10798;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10693;
    wire N__10690;
    wire N__10687;
    wire N__10686;
    wire N__10685;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10639;
    wire N__10636;
    wire N__10633;
    wire N__10628;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10600;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10586;
    wire N__10581;
    wire N__10578;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10558;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10528;
    wire N__10527;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10503;
    wire N__10500;
    wire N__10495;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10483;
    wire N__10478;
    wire N__10477;
    wire N__10476;
    wire N__10473;
    wire N__10470;
    wire N__10467;
    wire N__10460;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10411;
    wire N__10410;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10363;
    wire N__10360;
    wire N__10355;
    wire N__10354;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10311;
    wire N__10306;
    wire N__10303;
    wire N__10302;
    wire N__10301;
    wire N__10296;
    wire N__10295;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10280;
    wire N__10271;
    wire N__10268;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10260;
    wire N__10255;
    wire N__10252;
    wire N__10249;
    wire N__10248;
    wire N__10247;
    wire N__10242;
    wire N__10237;
    wire N__10232;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10224;
    wire N__10221;
    wire N__10218;
    wire N__10217;
    wire N__10216;
    wire N__10215;
    wire N__10212;
    wire N__10211;
    wire N__10206;
    wire N__10203;
    wire N__10200;
    wire N__10197;
    wire N__10194;
    wire N__10191;
    wire N__10186;
    wire N__10181;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10135;
    wire N__10134;
    wire N__10131;
    wire N__10126;
    wire N__10125;
    wire N__10120;
    wire N__10117;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10102;
    wire N__10099;
    wire N__10096;
    wire N__10093;
    wire N__10090;
    wire N__10087;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10054;
    wire N__10053;
    wire N__10052;
    wire N__10051;
    wire N__10050;
    wire N__10045;
    wire N__10040;
    wire N__10037;
    wire N__10036;
    wire N__10033;
    wire N__10028;
    wire N__10025;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__9998;
    wire N__9997;
    wire N__9996;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9988;
    wire N__9987;
    wire N__9984;
    wire N__9981;
    wire N__9978;
    wire N__9975;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9957;
    wire N__9954;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9922;
    wire N__9921;
    wire N__9920;
    wire N__9919;
    wire N__9918;
    wire N__9917;
    wire N__9916;
    wire N__9915;
    wire N__9914;
    wire N__9913;
    wire N__9912;
    wire N__9911;
    wire N__9910;
    wire N__9909;
    wire N__9908;
    wire N__9907;
    wire N__9904;
    wire N__9903;
    wire N__9902;
    wire N__9901;
    wire N__9900;
    wire N__9899;
    wire N__9898;
    wire N__9897;
    wire N__9896;
    wire N__9895;
    wire N__9842;
    wire N__9839;
    wire N__9838;
    wire N__9837;
    wire N__9834;
    wire N__9833;
    wire N__9830;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9801;
    wire N__9798;
    wire N__9793;
    wire N__9792;
    wire N__9787;
    wire N__9784;
    wire N__9779;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9742;
    wire N__9741;
    wire N__9740;
    wire N__9737;
    wire N__9736;
    wire N__9735;
    wire N__9732;
    wire N__9731;
    wire N__9728;
    wire N__9727;
    wire N__9726;
    wire N__9725;
    wire N__9724;
    wire N__9723;
    wire N__9720;
    wire N__9719;
    wire N__9718;
    wire N__9717;
    wire N__9716;
    wire N__9715;
    wire N__9714;
    wire N__9711;
    wire N__9710;
    wire N__9709;
    wire N__9704;
    wire N__9703;
    wire N__9702;
    wire N__9699;
    wire N__9696;
    wire N__9693;
    wire N__9690;
    wire N__9681;
    wire N__9678;
    wire N__9671;
    wire N__9666;
    wire N__9665;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9653;
    wire N__9650;
    wire N__9645;
    wire N__9640;
    wire N__9633;
    wire N__9626;
    wire N__9621;
    wire N__9602;
    wire N__9599;
    wire N__9598;
    wire N__9597;
    wire N__9594;
    wire N__9593;
    wire N__9592;
    wire N__9591;
    wire N__9590;
    wire N__9589;
    wire N__9588;
    wire N__9585;
    wire N__9584;
    wire N__9583;
    wire N__9582;
    wire N__9581;
    wire N__9578;
    wire N__9577;
    wire N__9576;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9568;
    wire N__9567;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9541;
    wire N__9536;
    wire N__9529;
    wire N__9524;
    wire N__9521;
    wire N__9520;
    wire N__9519;
    wire N__9514;
    wire N__9507;
    wire N__9496;
    wire N__9495;
    wire N__9492;
    wire N__9487;
    wire N__9484;
    wire N__9483;
    wire N__9480;
    wire N__9473;
    wire N__9470;
    wire N__9463;
    wire N__9460;
    wire N__9457;
    wire N__9454;
    wire N__9449;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9414;
    wire N__9413;
    wire N__9408;
    wire N__9405;
    wire N__9402;
    wire N__9395;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9360;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9347;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9283;
    wire N__9282;
    wire N__9275;
    wire N__9274;
    wire N__9273;
    wire N__9272;
    wire N__9271;
    wire N__9268;
    wire N__9265;
    wire N__9262;
    wire N__9261;
    wire N__9260;
    wire N__9255;
    wire N__9250;
    wire N__9247;
    wire N__9246;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9210;
    wire N__9205;
    wire N__9200;
    wire N__9197;
    wire N__9190;
    wire N__9185;
    wire N__9184;
    wire N__9181;
    wire N__9180;
    wire N__9179;
    wire N__9178;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9167;
    wire N__9160;
    wire N__9157;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9134;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9118;
    wire N__9113;
    wire N__9110;
    wire N__9109;
    wire N__9108;
    wire N__9105;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9094;
    wire N__9093;
    wire N__9092;
    wire N__9085;
    wire N__9084;
    wire N__9081;
    wire N__9078;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9039;
    wire N__9034;
    wire N__9031;
    wire N__9026;
    wire N__9023;
    wire N__9022;
    wire N__9021;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9007;
    wire N__9006;
    wire N__9003;
    wire N__8998;
    wire N__8997;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8971;
    wire N__8968;
    wire N__8965;
    wire N__8962;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8878;
    wire N__8875;
    wire N__8872;
    wire N__8871;
    wire N__8870;
    wire N__8869;
    wire N__8866;
    wire N__8865;
    wire N__8864;
    wire N__8863;
    wire N__8862;
    wire N__8861;
    wire N__8858;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8820;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8808;
    wire N__8805;
    wire N__8802;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8764;
    wire N__8761;
    wire N__8758;
    wire N__8755;
    wire N__8754;
    wire N__8751;
    wire N__8748;
    wire N__8745;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8635;
    wire N__8634;
    wire N__8631;
    wire N__8630;
    wire N__8629;
    wire N__8628;
    wire N__8625;
    wire N__8624;
    wire N__8623;
    wire N__8620;
    wire N__8617;
    wire N__8608;
    wire N__8601;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8581;
    wire N__8580;
    wire N__8579;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8569;
    wire N__8566;
    wire N__8563;
    wire N__8562;
    wire N__8561;
    wire N__8560;
    wire N__8559;
    wire N__8558;
    wire N__8557;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8534;
    wire N__8529;
    wire N__8526;
    wire N__8513;
    wire N__8510;
    wire N__8509;
    wire N__8506;
    wire N__8503;
    wire N__8498;
    wire N__8497;
    wire N__8494;
    wire N__8493;
    wire N__8492;
    wire N__8489;
    wire N__8488;
    wire N__8485;
    wire N__8480;
    wire N__8479;
    wire N__8476;
    wire N__8473;
    wire N__8470;
    wire N__8467;
    wire N__8464;
    wire N__8463;
    wire N__8462;
    wire N__8461;
    wire N__8460;
    wire N__8459;
    wire N__8458;
    wire N__8457;
    wire N__8456;
    wire N__8455;
    wire N__8450;
    wire N__8443;
    wire N__8438;
    wire N__8433;
    wire N__8432;
    wire N__8429;
    wire N__8420;
    wire N__8417;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8401;
    wire N__8392;
    wire N__8389;
    wire N__8386;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8363;
    wire N__8362;
    wire N__8359;
    wire N__8358;
    wire N__8355;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8339;
    wire N__8336;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8328;
    wire N__8325;
    wire N__8322;
    wire N__8319;
    wire N__8316;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8304;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8288;
    wire N__8285;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8257;
    wire N__8256;
    wire N__8253;
    wire N__8250;
    wire N__8249;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8233;
    wire N__8228;
    wire N__8225;
    wire N__8216;
    wire N__8213;
    wire N__8212;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8195;
    wire N__8194;
    wire N__8191;
    wire N__8186;
    wire N__8183;
    wire N__8180;
    wire N__8171;
    wire N__8170;
    wire N__8169;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8155;
    wire N__8154;
    wire N__8153;
    wire N__8148;
    wire N__8147;
    wire N__8142;
    wire N__8139;
    wire N__8136;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8122;
    wire N__8119;
    wire N__8116;
    wire N__8111;
    wire N__8108;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8098;
    wire N__8095;
    wire N__8094;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8060;
    wire N__8057;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8049;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8039;
    wire N__8034;
    wire N__8031;
    wire N__8028;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8005;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7954;
    wire N__7953;
    wire N__7952;
    wire N__7949;
    wire N__7948;
    wire N__7947;
    wire N__7946;
    wire N__7943;
    wire N__7942;
    wire N__7941;
    wire N__7940;
    wire N__7939;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7927;
    wire N__7924;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7908;
    wire N__7905;
    wire N__7886;
    wire N__7883;
    wire N__7882;
    wire N__7881;
    wire N__7878;
    wire N__7877;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7869;
    wire N__7868;
    wire N__7867;
    wire N__7864;
    wire N__7861;
    wire N__7858;
    wire N__7857;
    wire N__7856;
    wire N__7855;
    wire N__7854;
    wire N__7853;
    wire N__7852;
    wire N__7847;
    wire N__7840;
    wire N__7839;
    wire N__7832;
    wire N__7829;
    wire N__7828;
    wire N__7823;
    wire N__7816;
    wire N__7811;
    wire N__7808;
    wire N__7803;
    wire N__7800;
    wire N__7787;
    wire N__7784;
    wire N__7781;
    wire N__7778;
    wire N__7777;
    wire N__7776;
    wire N__7775;
    wire N__7772;
    wire N__7767;
    wire N__7764;
    wire N__7757;
    wire N__7754;
    wire N__7751;
    wire N__7748;
    wire N__7747;
    wire N__7746;
    wire N__7745;
    wire N__7742;
    wire N__7737;
    wire N__7734;
    wire N__7727;
    wire N__7724;
    wire N__7721;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7711;
    wire N__7708;
    wire N__7707;
    wire N__7704;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7685;
    wire N__7684;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7664;
    wire N__7661;
    wire N__7660;
    wire N__7659;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7651;
    wire N__7648;
    wire N__7645;
    wire N__7644;
    wire N__7643;
    wire N__7642;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7632;
    wire N__7629;
    wire N__7626;
    wire N__7621;
    wire N__7616;
    wire N__7601;
    wire N__7598;
    wire N__7595;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7585;
    wire N__7582;
    wire N__7581;
    wire N__7580;
    wire N__7579;
    wire N__7578;
    wire N__7577;
    wire N__7576;
    wire N__7575;
    wire N__7574;
    wire N__7573;
    wire N__7570;
    wire N__7567;
    wire N__7564;
    wire N__7561;
    wire N__7558;
    wire N__7555;
    wire N__7550;
    wire N__7543;
    wire N__7540;
    wire N__7523;
    wire N__7520;
    wire N__7519;
    wire N__7516;
    wire N__7515;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7507;
    wire N__7506;
    wire N__7505;
    wire N__7504;
    wire N__7501;
    wire N__7498;
    wire N__7495;
    wire N__7492;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7466;
    wire N__7465;
    wire N__7464;
    wire N__7463;
    wire N__7462;
    wire N__7461;
    wire N__7460;
    wire N__7457;
    wire N__7456;
    wire N__7455;
    wire N__7454;
    wire N__7451;
    wire N__7446;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7428;
    wire N__7425;
    wire N__7420;
    wire N__7417;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7381;
    wire N__7376;
    wire N__7373;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7342;
    wire N__7341;
    wire N__7338;
    wire N__7335;
    wire N__7332;
    wire N__7331;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7323;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7309;
    wire N__7306;
    wire N__7301;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7273;
    wire N__7272;
    wire N__7271;
    wire N__7270;
    wire N__7267;
    wire N__7262;
    wire N__7259;
    wire N__7256;
    wire N__7247;
    wire N__7246;
    wire N__7245;
    wire N__7242;
    wire N__7241;
    wire N__7238;
    wire N__7237;
    wire N__7236;
    wire N__7233;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7222;
    wire N__7219;
    wire N__7216;
    wire N__7215;
    wire N__7214;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7191;
    wire N__7188;
    wire N__7185;
    wire N__7182;
    wire N__7179;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7143;
    wire N__7140;
    wire N__7137;
    wire N__7134;
    wire N__7127;
    wire N__7124;
    wire N__7123;
    wire N__7120;
    wire N__7119;
    wire N__7118;
    wire N__7117;
    wire N__7114;
    wire N__7111;
    wire N__7108;
    wire N__7103;
    wire N__7094;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7084;
    wire N__7081;
    wire N__7080;
    wire N__7079;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7067;
    wire N__7066;
    wire N__7063;
    wire N__7062;
    wire N__7057;
    wire N__7054;
    wire N__7049;
    wire N__7046;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6974;
    wire N__6971;
    wire N__6968;
    wire N__6965;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6953;
    wire N__6950;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6942;
    wire N__6941;
    wire N__6938;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6920;
    wire N__6919;
    wire N__6914;
    wire N__6911;
    wire N__6908;
    wire N__6905;
    wire N__6902;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6710;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6661;
    wire N__6660;
    wire N__6657;
    wire N__6656;
    wire N__6655;
    wire N__6654;
    wire N__6653;
    wire N__6650;
    wire N__6649;
    wire N__6648;
    wire N__6645;
    wire N__6642;
    wire N__6635;
    wire N__6632;
    wire N__6627;
    wire N__6624;
    wire N__6611;
    wire N__6608;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6582;
    wire N__6579;
    wire N__6576;
    wire N__6573;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6548;
    wire N__6545;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6527;
    wire N__6524;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6512;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6499;
    wire N__6494;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6452;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6440;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6400;
    wire N__6399;
    wire N__6398;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6386;
    wire N__6383;
    wire N__6374;
    wire N__6371;
    wire N__6370;
    wire N__6369;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6357;
    wire N__6352;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6286;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6230;
    wire N__6227;
    wire N__6224;
    wire N__6223;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6206;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6191;
    wire N__6190;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6176;
    wire N__6173;
    wire N__6172;
    wire N__6169;
    wire N__6166;
    wire N__6163;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6148;
    wire N__6147;
    wire N__6144;
    wire N__6143;
    wire N__6140;
    wire N__6137;
    wire N__6134;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6126;
    wire N__6123;
    wire N__6120;
    wire N__6117;
    wire N__6112;
    wire N__6109;
    wire N__6106;
    wire N__6101;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6082;
    wire N__6079;
    wire N__6076;
    wire N__6071;
    wire N__6068;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6056;
    wire N__6053;
    wire N__6050;
    wire N__6049;
    wire N__6048;
    wire N__6047;
    wire N__6044;
    wire N__6041;
    wire N__6038;
    wire N__6035;
    wire N__6026;
    wire N__6025;
    wire N__6024;
    wire N__6023;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6012;
    wire N__6011;
    wire N__6008;
    wire N__6005;
    wire N__6000;
    wire N__5999;
    wire N__5998;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5983;
    wire N__5980;
    wire N__5973;
    wire N__5960;
    wire N__5959;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5942;
    wire N__5939;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5931;
    wire N__5926;
    wire N__5923;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5894;
    wire N__5893;
    wire N__5892;
    wire N__5891;
    wire N__5890;
    wire N__5889;
    wire N__5886;
    wire N__5881;
    wire N__5874;
    wire N__5867;
    wire N__5864;
    wire N__5863;
    wire N__5860;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5848;
    wire N__5845;
    wire N__5842;
    wire N__5839;
    wire N__5836;
    wire N__5833;
    wire N__5830;
    wire N__5827;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5804;
    wire N__5801;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5758;
    wire N__5757;
    wire N__5756;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5727;
    wire N__5724;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5644;
    wire N__5641;
    wire N__5636;
    wire N__5633;
    wire N__5630;
    wire N__5627;
    wire N__5624;
    wire N__5623;
    wire N__5622;
    wire N__5621;
    wire N__5620;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5602;
    wire N__5599;
    wire N__5588;
    wire N__5587;
    wire N__5584;
    wire N__5583;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5536;
    wire N__5535;
    wire N__5532;
    wire N__5529;
    wire N__5526;
    wire N__5519;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5459;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5387;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5254;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5237;
    wire N__5234;
    wire N__5233;
    wire N__5232;
    wire N__5231;
    wire N__5228;
    wire N__5221;
    wire N__5216;
    wire N__5213;
    wire N__5212;
    wire N__5209;
    wire N__5208;
    wire N__5207;
    wire N__5206;
    wire N__5203;
    wire N__5202;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5171;
    wire N__5170;
    wire N__5167;
    wire N__5166;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5154;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5125;
    wire N__5124;
    wire N__5123;
    wire N__5120;
    wire N__5119;
    wire N__5118;
    wire N__5115;
    wire N__5114;
    wire N__5113;
    wire N__5112;
    wire N__5109;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5094;
    wire N__5091;
    wire N__5084;
    wire N__5081;
    wire N__5066;
    wire N__5065;
    wire N__5064;
    wire N__5063;
    wire N__5062;
    wire N__5059;
    wire N__5058;
    wire N__5055;
    wire N__5054;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5046;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5020;
    wire N__5017;
    wire N__5000;
    wire N__4999;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4982;
    wire N__4981;
    wire N__4980;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4968;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4954;
    wire N__4951;
    wire N__4948;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4889;
    wire N__4888;
    wire N__4887;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4865;
    wire N__4864;
    wire N__4863;
    wire N__4862;
    wire N__4861;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4825;
    wire N__4822;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4787;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4748;
    wire N__4745;
    wire N__4742;
    wire N__4739;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4727;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4715;
    wire N__4712;
    wire N__4709;
    wire N__4706;
    wire N__4703;
    wire N__4700;
    wire N__4697;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4672;
    wire N__4669;
    wire N__4666;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4589;
    wire N__4588;
    wire N__4585;
    wire N__4582;
    wire N__4577;
    wire N__4576;
    wire N__4573;
    wire N__4570;
    wire N__4567;
    wire N__4562;
    wire N__4561;
    wire N__4558;
    wire N__4555;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4508;
    wire N__4507;
    wire N__4506;
    wire N__4505;
    wire N__4502;
    wire N__4497;
    wire N__4494;
    wire N__4487;
    wire N__4486;
    wire N__4485;
    wire N__4484;
    wire N__4483;
    wire N__4482;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4462;
    wire N__4457;
    wire N__4448;
    wire N__4447;
    wire N__4446;
    wire N__4443;
    wire N__4438;
    wire N__4433;
    wire N__4430;
    wire N__4427;
    wire N__4426;
    wire N__4423;
    wire N__4420;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4384;
    wire N__4381;
    wire N__4378;
    wire N__4375;
    wire N__4372;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4345;
    wire N__4342;
    wire N__4339;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4324;
    wire N__4323;
    wire N__4318;
    wire N__4315;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4294;
    wire N__4291;
    wire N__4288;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4267;
    wire N__4266;
    wire N__4263;
    wire N__4260;
    wire N__4257;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4231;
    wire N__4230;
    wire N__4229;
    wire N__4228;
    wire N__4227;
    wire N__4226;
    wire N__4225;
    wire N__4224;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4139;
    wire N__4136;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_PLL_i_i;
    wire N_882_i;
    wire \U712_REG_SM.N_71_i_cascade_ ;
    wire TACK_EN_i_ess;
    wire \U712_REG_SM.N_265_cascade_ ;
    wire ASn_c;
    wire \INVU712_REG_SM.STATE_COUNTER_9C_net ;
    wire REGENn_c;
    wire \INVU712_REG_SM.REGENnC_net ;
    wire VBENn_c;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_8_10_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_REG_SM.N_330_cascade_ ;
    wire \INVU712_REG_SM.LDSnC_net ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0 ;
    wire TACK_OUTn;
    wire \U712_REG_SM.N_295_cascade_ ;
    wire \U712_REG_SM.LDSn_6_iv_i_0_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_REG_SM.N_332 ;
    wire \U712_REG_SM.UDSn_6_iv_i_0_0 ;
    wire \U712_REG_SM.STATE_COUNTER_RNI7KTS1Z0Z_9 ;
    wire UDSn_c;
    wire \U712_REG_SM.N_266 ;
    wire \U712_REG_SM.STATE_COUNTER_srsts_i_i_i_a3_3_0_cascade_ ;
    wire REGSPACEn_c;
    wire \U712_REG_SM.CYCLE_RUNZ0 ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \INVU712_REG_SM.UDSnC_net ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_9 ;
    wire \U712_REG_SM.N_71_i ;
    wire REG_CPU_CYCLE;
    wire \INVU712_REG_SM.LATCH_REGC_net ;
    wire C3_c;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \INVU712_REG_SM.C3_SYNC_0C_net ;
    wire A_c_3;
    wire \U712_CHIP_RAM.N_241_cascade_ ;
    wire \U712_BYTE_ENABLE.N_276 ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0_cascade_ ;
    wire N_47_i;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire A_c_14;
    wire A_c_7;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5_cascade_ ;
    wire DBRn_c_i_0;
    wire A_c_20;
    wire \U712_CHIP_RAM.N_361_cascade_ ;
    wire BANK0_c;
    wire \U712_CHIP_RAM.N_452 ;
    wire \U712_CHIP_RAM.N_452_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0 ;
    wire LDSn_c;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_0 ;
    wire \U712_REG_SM.N_309 ;
    wire \U712_REG_SM.STATE_COUNTER_srsts_i_i_i_a3_2_0 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_5 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_7 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_3 ;
    wire \U712_REG_SM.un18_0_i_0_0_1_cascade_ ;
    wire \INVU712_REG_SM.STATE_COUNTER_5C_net ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_8 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_4 ;
    wire \U712_REG_SM.N_442_cascade_ ;
    wire \U712_REG_SM.REG_CPU_CYCLE_e_1 ;
    wire \U712_REG_SM.N_84 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_447 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_6 ;
    wire \U712_REG_SM.N_288 ;
    wire LATCH_REG;
    wire LATCH_CLK_0_i;
    wire A_c_8;
    wire A_c_15;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ;
    wire A_c_13;
    wire A_c_6;
    wire A_c_16;
    wire A_c_18;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.un1_CMA28_0_i ;
    wire A_c_11;
    wire A_c_4;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_1 ;
    wire \U712_CHIP_RAM.N_325_cascade_ ;
    wire \U712_CHIP_RAM.N_301 ;
    wire \U712_CHIP_RAM.N_392_cascade_ ;
    wire \U712_CHIP_RAM.N_449 ;
    wire \U712_CHIP_RAM.N_376_cascade_ ;
    wire \U712_CHIP_RAM.N_45_i_cascade_ ;
    wire \U712_CHIP_RAM.N_324_2 ;
    wire \U712_CHIP_RAM.N_324_2_cascade_ ;
    wire \U712_CHIP_RAM.N_450 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVCZ0Z_4 ;
    wire \U712_CHIP_RAM.N_252 ;
    wire \U712_CHIP_RAM.N_252_cascade_ ;
    wire \U712_CHIP_RAM.N_365_1_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0 ;
    wire RnW_c;
    wire CLK_EN_c;
    wire RAMSPACEn_c;
    wire TSn_c;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire DBR_SYNCZ0Z_1;
    wire DBR_SYNCZ0Z_0;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ;
    wire LATCH_RAM;
    wire \U712_REG_SM.N_265 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTERZ0Z_2 ;
    wire \U712_REG_SM.DBR_SYNCZ0Z_1 ;
    wire DBRn_c;
    wire \U712_REG_SM.DBR_SYNCZ0Z_0 ;
    wire \INVU712_REG_SM.STATE_COUNTER_2C_net ;
    wire REG_WRITE_CYCLE;
    wire N_289;
    wire A_c_5;
    wire A_c_12;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ;
    wire \U712_CHIP_RAM.CMA_5_0_8_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ;
    wire A_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire AWEn_c;
    wire DBDIR_c;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH5lt7 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.N_324 ;
    wire \U712_CHIP_RAM.N_456_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1 ;
    wire bfn_11_11_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.N_363 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.N_384_cascade_ ;
    wire \U712_CHIP_RAM.N_448_cascade_ ;
    wire \U712_CHIP_RAM.N_255 ;
    wire \U712_CHIP_RAM.N_255_cascade_ ;
    wire \U712_CHIP_RAM.N_269 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0_0 ;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_444 ;
    wire \U712_CHIP_RAM.N_392 ;
    wire \U712_CHIP_RAM.N_444_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0 ;
    wire \U712_CHIP_RAM.N_334 ;
    wire \U712_CHIP_RAM.N_334_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0 ;
    wire \U712_CHIP_RAM.N_448 ;
    wire \U712_CHIP_RAM.N_323 ;
    wire \U712_CHIP_RAM.N_323_cascade_ ;
    wire \U712_CHIP_RAM.un3_DMA_CYCLE_START ;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire CMA_c_2;
    wire N_46_i;
    wire \U712_BYTE_ENABLE.UUBE_cascade_ ;
    wire N_48_i;
    wire \U712_BYTE_ENABLE.N_278 ;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0 ;
    wire N_49_i;
    wire \U712_BYTE_ENABLE.N_277 ;
    wire DBENn_c;
    wire \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0Z0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_2_0 ;
    wire \U712_CHIP_RAM.N_325_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ;
    wire \U712_CHIP_RAM.N_365_1 ;
    wire \U712_CHIP_RAM.N_294 ;
    wire DMA_CYCLE;
    wire \U712_CHIP_RAM.N_305_cascade_ ;
    wire \U712_CHIP_RAM.N_388 ;
    wire \U712_CHIP_RAM.N_45_i ;
    wire \U712_CHIP_RAM.N_346_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_2 ;
    wire \U712_CHIP_RAM.N_407 ;
    wire \U712_CHIP_RAM.N_407_cascade_ ;
    wire \U712_CHIP_RAM.N_400 ;
    wire WRITE_CYCLE;
    wire \U712_CHIP_RAM.N_257_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_396_cascade_ ;
    wire \U712_CHIP_RAM.N_436 ;
    wire \U712_CHIP_RAM.N_436_cascade_ ;
    wire \U712_CHIP_RAM.N_257 ;
    wire \U712_CHIP_RAM.N_357 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_1 ;
    wire \U712_CHIP_RAM.N_396 ;
    wire \U712_CHIP_RAM.N_384 ;
    wire \U712_CHIP_RAM.N_351 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_cascade_ ;
    wire \U712_CHIP_RAM.N_117 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_0_a2_0_2 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.N_274_i_0_0_cascade_ ;
    wire \U712_CYCLE_TERM.N_274_i_0_en_cascade_ ;
    wire \U712_CYCLE_TERM.N_274_i_0_en_0 ;
    wire \U712_CHIP_RAM.N_456 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire \U712_CHIP_RAM.N_202 ;
    wire \U712_CHIP_RAM.N_359 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire RESETn_c;
    wire RESETn_c_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire CLK40_PLL;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_2 ;
    wire \U712_CYCLE_TERM.N_8 ;
    wire REG_TACK;
    wire CPU_TACK;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire CASLn_c;
    wire CASUn_c;
    wire REG_CYCLE;
    wire DRDENn_c;
    wire CLK40_PLL_g;
    wire CLK40_PLL_iso_i;
    wire U712_BYTE_ENABLE_UUBE_i;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire A_c_17;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ;
    wire N_276_i;
    wire N_278_i;
    wire A_c_0;
    wire SIZ_c_0;
    wire A_c_1;
    wire SIZ_c_1;
    wire N_277_i;
    wire CRCSn_c;
    wire RASn_c;
    wire CASn_c;
    wire WEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire RAS0n_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire \U712_CHIP_RAM.CMA_5_sn_N_5_mux ;
    wire \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ;
    wire CMA_c_0;
    wire CLK80_PLL;
    wire \U712_CHIP_RAM.un1_CMA28_0_i_0 ;
    wire A_c_9;
    wire A_c_2;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CPU_CYCLE;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_AZ0Z20 ;
    wire \INVU712_CHIP_RAM.DMA_A20C_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire DRA_c_7;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire AGNUS_REV_c;
    wire DRA_c_0;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire _gnd_net_;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL),
            .REFERENCECLK(N__4061),
            .RESETB(N__6878),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__12003),
            .DIN(N__12002),
            .DOUT(N__12001),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__12003),
            .PADOUT(N__12002),
            .PADIN(N__12001),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6959),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__11994),
            .DIN(N__11993),
            .DOUT(N__11992),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__11994),
            .PADOUT(N__11993),
            .PADIN(N__11992),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__11985),
            .DIN(N__11984),
            .DOUT(N__11983),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__11985),
            .PADOUT(N__11984),
            .PADIN(N__11983),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8897),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__11976),
            .DIN(N__11975),
            .DOUT(N__11974),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__11976),
            .PADOUT(N__11975),
            .PADIN(N__11974),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5867),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__11967),
            .DIN(N__11966),
            .DOUT(N__11965),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__11967),
            .PADOUT(N__11966),
            .PADIN(N__11965),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__11958),
            .DIN(N__11957),
            .DOUT(N__11956),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__11958),
            .PADOUT(N__11957),
            .PADIN(N__11956),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__11949),
            .DIN(N__11948),
            .DOUT(N__11947),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__11949),
            .PADOUT(N__11948),
            .PADIN(N__11947),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__11940),
            .DIN(N__11939),
            .DOUT(N__11938),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__11940),
            .PADOUT(N__11939),
            .PADIN(N__11938),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__11931),
            .DIN(N__11930),
            .DOUT(N__11929),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__11931),
            .PADOUT(N__11930),
            .PADIN(N__11929),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__11922),
            .DIN(N__11921),
            .DOUT(N__11920),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__11922),
            .PADOUT(N__11921),
            .PADIN(N__11920),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__11913),
            .DIN(N__11912),
            .DOUT(N__11911),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__11913),
            .PADOUT(N__11912),
            .PADIN(N__11911),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6857),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__11904),
            .DIN(N__11903),
            .DOUT(N__11902),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__11904),
            .PADOUT(N__11903),
            .PADIN(N__11902),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8780),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__11895),
            .DIN(N__11894),
            .DOUT(N__11893),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__11895),
            .PADOUT(N__11894),
            .PADIN(N__11893),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__11886),
            .DIN(N__11885),
            .DOUT(N__11884),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__11886),
            .PADOUT(N__11885),
            .PADIN(N__11884),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__11877),
            .DIN(N__11876),
            .DOUT(N__11875),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__11877),
            .PADOUT(N__11876),
            .PADIN(N__11875),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__11868),
            .DIN(N__11867),
            .DOUT(N__11866),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__11868),
            .PADOUT(N__11867),
            .PADIN(N__11866),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4139),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__11859),
            .DIN(N__11858),
            .DOUT(N__11857),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__11859),
            .PADOUT(N__11858),
            .PADIN(N__11857),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__11850),
            .DIN(N__11849),
            .DOUT(N__11848),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__11850),
            .PADOUT(N__11849),
            .PADIN(N__11848),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__11841),
            .DIN(N__11840),
            .DOUT(N__11839),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__11841),
            .PADOUT(N__11840),
            .PADIN(N__11839),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9947),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__11832),
            .DIN(N__11831),
            .DOUT(N__11830),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__11832),
            .PADOUT(N__11831),
            .PADIN(N__11830),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__11823),
            .DIN(N__11822),
            .DOUT(N__11821),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__11823),
            .PADOUT(N__11822),
            .PADIN(N__11821),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8936),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__11814),
            .DIN(N__11813),
            .DOUT(N__11812),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__11814),
            .PADOUT(N__11813),
            .PADIN(N__11812),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__11805),
            .DIN(N__11804),
            .DOUT(N__11803),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__11805),
            .PADOUT(N__11804),
            .PADIN(N__11803),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9314),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__11796),
            .DIN(N__11795),
            .DOUT(N__11794),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__11796),
            .PADOUT(N__11795),
            .PADIN(N__11794),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__11787),
            .DIN(N__11786),
            .DOUT(N__11785),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__11787),
            .PADOUT(N__11786),
            .PADIN(N__11785),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__11778),
            .DIN(N__11777),
            .DOUT(N__11776),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__11778),
            .PADOUT(N__11777),
            .PADIN(N__11776),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__11769),
            .DIN(N__11768),
            .DOUT(N__11767),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__11769),
            .PADOUT(N__11768),
            .PADIN(N__11767),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__11760),
            .DIN(N__11759),
            .DOUT(N__11758),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__11760),
            .PADOUT(N__11759),
            .PADIN(N__11758),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__11751),
            .DIN(N__11750),
            .DOUT(N__11749),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__11751),
            .PADOUT(N__11750),
            .PADIN(N__11749),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5863),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__11742),
            .DIN(N__11741),
            .DOUT(N__11740),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__11742),
            .PADOUT(N__11741),
            .PADIN(N__11740),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__11733),
            .DIN(N__11732),
            .DOUT(N__11731),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__11733),
            .PADOUT(N__11732),
            .PADIN(N__11731),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__11724),
            .DIN(N__11723),
            .DOUT(N__11722),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__11724),
            .PADOUT(N__11723),
            .PADIN(N__11722),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__11715),
            .DIN(N__11714),
            .DOUT(N__11713),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__11715),
            .PADOUT(N__11714),
            .PADIN(N__11713),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__11706),
            .DIN(N__11705),
            .DOUT(N__11704),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__11706),
            .PADOUT(N__11705),
            .PADIN(N__11704),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__11697),
            .DIN(N__11696),
            .DOUT(N__11695),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__11697),
            .PADOUT(N__11696),
            .PADIN(N__11695),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8918),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__11688),
            .DIN(N__11687),
            .DOUT(N__11686),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__11688),
            .PADOUT(N__11687),
            .PADIN(N__11686),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4733),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11679),
            .DIN(N__11678),
            .DOUT(N__11677),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11679),
            .PADOUT(N__11678),
            .PADIN(N__11677),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8827),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11670),
            .DIN(N__11669),
            .DOUT(N__11668),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11670),
            .PADOUT(N__11669),
            .PADIN(N__11668),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4115),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__11661),
            .DIN(N__11660),
            .DOUT(N__11659),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__11661),
            .PADOUT(N__11660),
            .PADIN(N__11659),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__11652),
            .DIN(N__11651),
            .DOUT(N__11650),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__11652),
            .PADOUT(N__11651),
            .PADIN(N__11650),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4196),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11643),
            .DIN(N__11642),
            .DOUT(N__11641),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11643),
            .PADOUT(N__11642),
            .PADIN(N__11641),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6803),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11634),
            .DIN(N__11633),
            .DOUT(N__11632),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11634),
            .PADOUT(N__11633),
            .PADIN(N__11632),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11625),
            .DIN(N__11624),
            .DOUT(N__11623),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11625),
            .PADOUT(N__11624),
            .PADIN(N__11623),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11616),
            .DIN(N__11615),
            .DOUT(N__11614),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11616),
            .PADOUT(N__11615),
            .PADIN(N__11614),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__11607),
            .DIN(N__11606),
            .DOUT(N__11605),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__11607),
            .PADOUT(N__11606),
            .PADIN(N__11605),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__11598),
            .DIN(N__11597),
            .DOUT(N__11596),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__11598),
            .PADOUT(N__11597),
            .PADIN(N__11596),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10172),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11589),
            .DIN(N__11588),
            .DOUT(N__11587),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11589),
            .PADOUT(N__11588),
            .PADIN(N__11587),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11580),
            .DIN(N__11579),
            .DOUT(N__11578),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11580),
            .PADOUT(N__11579),
            .PADIN(N__11578),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8820),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__11571),
            .DIN(N__11570),
            .DOUT(N__11569),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__11571),
            .PADOUT(N__11570),
            .PADIN(N__11569),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6830),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11562),
            .DIN(N__11561),
            .DOUT(N__11560),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11562),
            .PADOUT(N__11561),
            .PADIN(N__11560),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7976),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11553),
            .DIN(N__11552),
            .DOUT(N__11551),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11553),
            .PADOUT(N__11552),
            .PADIN(N__11551),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4622),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11544),
            .DIN(N__11543),
            .DOUT(N__11542),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11544),
            .PADOUT(N__11543),
            .PADIN(N__11542),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6734),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__11535),
            .DIN(N__11534),
            .DOUT(N__11533),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__11535),
            .PADOUT(N__11534),
            .PADIN(N__11533),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4166),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__11526),
            .DIN(N__11525),
            .DOUT(N__11524),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__11526),
            .PADOUT(N__11525),
            .PADIN(N__11524),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__11517),
            .DIN(N__11516),
            .DOUT(N__11515),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__11517),
            .PADOUT(N__11516),
            .PADIN(N__11515),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__11508),
            .DIN(N__11507),
            .DOUT(N__11506),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__11508),
            .PADOUT(N__11507),
            .PADIN(N__11506),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6986),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__11499),
            .DIN(N__11498),
            .DOUT(N__11497),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__11499),
            .PADOUT(N__11498),
            .PADIN(N__11497),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10340),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__11490),
            .DIN(N__11489),
            .DOUT(N__11488),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__11490),
            .PADOUT(N__11489),
            .PADIN(N__11488),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6233),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__11481),
            .DIN(N__11480),
            .DOUT(N__11479),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__11481),
            .PADOUT(N__11480),
            .PADIN(N__11479),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6692),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__11472),
            .DIN(N__11471),
            .DOUT(N__11470),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__11472),
            .PADOUT(N__11471),
            .PADIN(N__11470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__11463),
            .DIN(N__11462),
            .DOUT(N__11461),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__11463),
            .PADOUT(N__11462),
            .PADIN(N__11461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__11454),
            .DIN(N__11453),
            .DOUT(N__11452),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__11454),
            .PADOUT(N__11453),
            .PADIN(N__11452),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__11445),
            .DIN(N__11444),
            .DOUT(N__11443),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__11445),
            .PADOUT(N__11444),
            .PADIN(N__11443),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__11436),
            .DIN(N__11435),
            .DOUT(N__11434),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__11436),
            .PADOUT(N__11435),
            .PADIN(N__11434),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5315),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__11427),
            .DIN(N__11426),
            .DOUT(N__11425),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__11427),
            .PADOUT(N__11426),
            .PADIN(N__11425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9299),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__11418),
            .DIN(N__11417),
            .DOUT(N__11416),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__11418),
            .PADOUT(N__11417),
            .PADIN(N__11416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__11409),
            .DIN(N__11408),
            .DOUT(N__11407),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__11409),
            .PADOUT(N__11408),
            .PADIN(N__11407),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7031),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__11400),
            .DIN(N__11399),
            .DOUT(N__11398),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__11400),
            .PADOUT(N__11399),
            .PADIN(N__11398),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4100),
            .DIN0(),
            .DOUT0(N__4361),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__11391),
            .DIN(N__11390),
            .DOUT(N__11389),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__11391),
            .PADOUT(N__11390),
            .PADIN(N__11389),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6713),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__11382),
            .DIN(N__11381),
            .DOUT(N__11380),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__11382),
            .PADOUT(N__11381),
            .PADIN(N__11380),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__11373),
            .DIN(N__11372),
            .DOUT(N__11371),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__11373),
            .PADOUT(N__11372),
            .PADIN(N__11371),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__11364),
            .DIN(N__11363),
            .DOUT(N__11362),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__11364),
            .PADOUT(N__11363),
            .PADIN(N__11362),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8717),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__11355),
            .DIN(N__11354),
            .DOUT(N__11353),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__11355),
            .PADOUT(N__11354),
            .PADIN(N__11353),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__11346),
            .DIN(N__11345),
            .DOUT(N__11344),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__11346),
            .PADOUT(N__11345),
            .PADIN(N__11344),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11337),
            .DIN(N__11336),
            .DOUT(N__11335),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11337),
            .PADOUT(N__11336),
            .PADIN(N__11335),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11328),
            .DIN(N__11327),
            .DOUT(N__11326),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11328),
            .PADOUT(N__11327),
            .PADIN(N__11326),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__11319),
            .DIN(N__11318),
            .DOUT(N__11317),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__11319),
            .PADOUT(N__11318),
            .PADIN(N__11317),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5342),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__11310),
            .DIN(N__11309),
            .DOUT(N__11308),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__11310),
            .PADOUT(N__11309),
            .PADIN(N__11308),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4283),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__11301),
            .DIN(N__11300),
            .DOUT(N__11299),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__11301),
            .PADOUT(N__11300),
            .PADIN(N__11299),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8954),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__11292),
            .DIN(N__11291),
            .DOUT(N__11290),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__11292),
            .PADOUT(N__11291),
            .PADIN(N__11290),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5702),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__11283),
            .DIN(N__11282),
            .DOUT(N__11281),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__11283),
            .PADOUT(N__11282),
            .PADIN(N__11281),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11274),
            .DIN(N__11273),
            .DOUT(N__11272),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11274),
            .PADOUT(N__11273),
            .PADIN(N__11272),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__11265),
            .DIN(N__11264),
            .DOUT(N__11263),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__11265),
            .PADOUT(N__11264),
            .PADIN(N__11263),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6773),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__11256),
            .DIN(N__11255),
            .DOUT(N__11254),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__11256),
            .PADOUT(N__11255),
            .PADIN(N__11254),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__11247),
            .DIN(N__11246),
            .DOUT(N__11245),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__11247),
            .PADOUT(N__11246),
            .PADIN(N__11245),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__11238),
            .DIN(N__11237),
            .DOUT(N__11236),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__11238),
            .PADOUT(N__11237),
            .PADIN(N__11236),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4943),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__11229),
            .DIN(N__11228),
            .DOUT(N__11227),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__11229),
            .PADOUT(N__11228),
            .PADIN(N__11227),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4907),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11220),
            .DIN(N__11219),
            .DOUT(N__11218),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11220),
            .PADOUT(N__11219),
            .PADIN(N__11218),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8831),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11211),
            .DIN(N__11210),
            .DOUT(N__11209),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11211),
            .PADOUT(N__11210),
            .PADIN(N__11209),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__2739 (
            .O(N__11192),
            .I(N__11189));
    InMux I__2738 (
            .O(N__11189),
            .I(N__11185));
    CascadeMux I__2737 (
            .O(N__11188),
            .I(N__11178));
    LocalMux I__2736 (
            .O(N__11185),
            .I(N__11174));
    InMux I__2735 (
            .O(N__11184),
            .I(N__11169));
    InMux I__2734 (
            .O(N__11183),
            .I(N__11169));
    InMux I__2733 (
            .O(N__11182),
            .I(N__11164));
    InMux I__2732 (
            .O(N__11181),
            .I(N__11164));
    InMux I__2731 (
            .O(N__11178),
            .I(N__11158));
    InMux I__2730 (
            .O(N__11177),
            .I(N__11158));
    Span4Mux_v I__2729 (
            .O(N__11174),
            .I(N__11147));
    LocalMux I__2728 (
            .O(N__11169),
            .I(N__11142));
    LocalMux I__2727 (
            .O(N__11164),
            .I(N__11142));
    InMux I__2726 (
            .O(N__11163),
            .I(N__11139));
    LocalMux I__2725 (
            .O(N__11158),
            .I(N__11136));
    InMux I__2724 (
            .O(N__11157),
            .I(N__11133));
    InMux I__2723 (
            .O(N__11156),
            .I(N__11126));
    InMux I__2722 (
            .O(N__11155),
            .I(N__11126));
    InMux I__2721 (
            .O(N__11154),
            .I(N__11126));
    InMux I__2720 (
            .O(N__11153),
            .I(N__11123));
    InMux I__2719 (
            .O(N__11152),
            .I(N__11120));
    InMux I__2718 (
            .O(N__11151),
            .I(N__11117));
    InMux I__2717 (
            .O(N__11150),
            .I(N__11114));
    Span4Mux_h I__2716 (
            .O(N__11147),
            .I(N__11105));
    Span4Mux_v I__2715 (
            .O(N__11142),
            .I(N__11105));
    LocalMux I__2714 (
            .O(N__11139),
            .I(N__11105));
    Span4Mux_h I__2713 (
            .O(N__11136),
            .I(N__11100));
    LocalMux I__2712 (
            .O(N__11133),
            .I(N__11100));
    LocalMux I__2711 (
            .O(N__11126),
            .I(N__11088));
    LocalMux I__2710 (
            .O(N__11123),
            .I(N__11088));
    LocalMux I__2709 (
            .O(N__11120),
            .I(N__11088));
    LocalMux I__2708 (
            .O(N__11117),
            .I(N__11088));
    LocalMux I__2707 (
            .O(N__11114),
            .I(N__11088));
    InMux I__2706 (
            .O(N__11113),
            .I(N__11084));
    InMux I__2705 (
            .O(N__11112),
            .I(N__11080));
    Span4Mux_h I__2704 (
            .O(N__11105),
            .I(N__11075));
    Span4Mux_v I__2703 (
            .O(N__11100),
            .I(N__11075));
    InMux I__2702 (
            .O(N__11099),
            .I(N__11072));
    Span4Mux_v I__2701 (
            .O(N__11088),
            .I(N__11069));
    InMux I__2700 (
            .O(N__11087),
            .I(N__11066));
    LocalMux I__2699 (
            .O(N__11084),
            .I(N__11063));
    InMux I__2698 (
            .O(N__11083),
            .I(N__11060));
    LocalMux I__2697 (
            .O(N__11080),
            .I(N__11057));
    Sp12to4 I__2696 (
            .O(N__11075),
            .I(N__11048));
    LocalMux I__2695 (
            .O(N__11072),
            .I(N__11048));
    Sp12to4 I__2694 (
            .O(N__11069),
            .I(N__11048));
    LocalMux I__2693 (
            .O(N__11066),
            .I(N__11048));
    Sp12to4 I__2692 (
            .O(N__11063),
            .I(N__11043));
    LocalMux I__2691 (
            .O(N__11060),
            .I(N__11043));
    Span12Mux_h I__2690 (
            .O(N__11057),
            .I(N__11040));
    Span12Mux_h I__2689 (
            .O(N__11048),
            .I(N__11037));
    Span12Mux_v I__2688 (
            .O(N__11043),
            .I(N__11034));
    Span12Mux_v I__2687 (
            .O(N__11040),
            .I(N__11031));
    Span12Mux_v I__2686 (
            .O(N__11037),
            .I(N__11026));
    Span12Mux_h I__2685 (
            .O(N__11034),
            .I(N__11026));
    Odrv12 I__2684 (
            .O(N__11031),
            .I(AGNUS_REV_c));
    Odrv12 I__2683 (
            .O(N__11026),
            .I(AGNUS_REV_c));
    InMux I__2682 (
            .O(N__11021),
            .I(N__11017));
    InMux I__2681 (
            .O(N__11020),
            .I(N__11014));
    LocalMux I__2680 (
            .O(N__11017),
            .I(N__11009));
    LocalMux I__2679 (
            .O(N__11014),
            .I(N__11009));
    Sp12to4 I__2678 (
            .O(N__11009),
            .I(N__11006));
    Span12Mux_v I__2677 (
            .O(N__11006),
            .I(N__11003));
    Span12Mux_h I__2676 (
            .O(N__11003),
            .I(N__11000));
    Odrv12 I__2675 (
            .O(N__11000),
            .I(DRA_c_0));
    InMux I__2674 (
            .O(N__10997),
            .I(N__10992));
    InMux I__2673 (
            .O(N__10996),
            .I(N__10988));
    InMux I__2672 (
            .O(N__10995),
            .I(N__10985));
    LocalMux I__2671 (
            .O(N__10992),
            .I(N__10982));
    InMux I__2670 (
            .O(N__10991),
            .I(N__10979));
    LocalMux I__2669 (
            .O(N__10988),
            .I(N__10972));
    LocalMux I__2668 (
            .O(N__10985),
            .I(N__10972));
    Span4Mux_v I__2667 (
            .O(N__10982),
            .I(N__10972));
    LocalMux I__2666 (
            .O(N__10979),
            .I(N__10969));
    Sp12to4 I__2665 (
            .O(N__10972),
            .I(N__10966));
    Span4Mux_h I__2664 (
            .O(N__10969),
            .I(N__10963));
    Span12Mux_h I__2663 (
            .O(N__10966),
            .I(N__10958));
    Sp12to4 I__2662 (
            .O(N__10963),
            .I(N__10958));
    Span12Mux_v I__2661 (
            .O(N__10958),
            .I(N__10955));
    Odrv12 I__2660 (
            .O(N__10955),
            .I(DRA_c_1));
    InMux I__2659 (
            .O(N__10952),
            .I(N__10949));
    LocalMux I__2658 (
            .O(N__10949),
            .I(N__10946));
    Odrv4 I__2657 (
            .O(N__10946),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    ClkMux I__2656 (
            .O(N__10943),
            .I(N__10925));
    ClkMux I__2655 (
            .O(N__10942),
            .I(N__10925));
    ClkMux I__2654 (
            .O(N__10941),
            .I(N__10925));
    ClkMux I__2653 (
            .O(N__10940),
            .I(N__10925));
    ClkMux I__2652 (
            .O(N__10939),
            .I(N__10925));
    ClkMux I__2651 (
            .O(N__10938),
            .I(N__10925));
    GlobalMux I__2650 (
            .O(N__10925),
            .I(N__10922));
    gio2CtrlBuf I__2649 (
            .O(N__10922),
            .I(C3_c_g));
    CEMux I__2648 (
            .O(N__10919),
            .I(N__10880));
    CEMux I__2647 (
            .O(N__10918),
            .I(N__10880));
    CEMux I__2646 (
            .O(N__10917),
            .I(N__10880));
    CEMux I__2645 (
            .O(N__10916),
            .I(N__10880));
    CEMux I__2644 (
            .O(N__10915),
            .I(N__10880));
    CEMux I__2643 (
            .O(N__10914),
            .I(N__10880));
    CEMux I__2642 (
            .O(N__10913),
            .I(N__10880));
    CEMux I__2641 (
            .O(N__10912),
            .I(N__10880));
    CEMux I__2640 (
            .O(N__10911),
            .I(N__10880));
    CEMux I__2639 (
            .O(N__10910),
            .I(N__10880));
    CEMux I__2638 (
            .O(N__10909),
            .I(N__10880));
    CEMux I__2637 (
            .O(N__10908),
            .I(N__10880));
    CEMux I__2636 (
            .O(N__10907),
            .I(N__10880));
    GlobalMux I__2635 (
            .O(N__10880),
            .I(N__10877));
    gio2CtrlBuf I__2634 (
            .O(N__10877),
            .I(DBRn_c_i_0_g));
    InMux I__2633 (
            .O(N__10874),
            .I(N__10867));
    InMux I__2632 (
            .O(N__10873),
            .I(N__10864));
    InMux I__2631 (
            .O(N__10872),
            .I(N__10861));
    InMux I__2630 (
            .O(N__10871),
            .I(N__10858));
    InMux I__2629 (
            .O(N__10870),
            .I(N__10855));
    LocalMux I__2628 (
            .O(N__10867),
            .I(N__10841));
    LocalMux I__2627 (
            .O(N__10864),
            .I(N__10833));
    LocalMux I__2626 (
            .O(N__10861),
            .I(N__10825));
    LocalMux I__2625 (
            .O(N__10858),
            .I(N__10816));
    LocalMux I__2624 (
            .O(N__10855),
            .I(N__10803));
    SRMux I__2623 (
            .O(N__10854),
            .I(N__10703));
    SRMux I__2622 (
            .O(N__10853),
            .I(N__10703));
    SRMux I__2621 (
            .O(N__10852),
            .I(N__10703));
    SRMux I__2620 (
            .O(N__10851),
            .I(N__10703));
    SRMux I__2619 (
            .O(N__10850),
            .I(N__10703));
    SRMux I__2618 (
            .O(N__10849),
            .I(N__10703));
    SRMux I__2617 (
            .O(N__10848),
            .I(N__10703));
    SRMux I__2616 (
            .O(N__10847),
            .I(N__10703));
    SRMux I__2615 (
            .O(N__10846),
            .I(N__10703));
    SRMux I__2614 (
            .O(N__10845),
            .I(N__10703));
    SRMux I__2613 (
            .O(N__10844),
            .I(N__10703));
    Glb2LocalMux I__2612 (
            .O(N__10841),
            .I(N__10703));
    SRMux I__2611 (
            .O(N__10840),
            .I(N__10703));
    SRMux I__2610 (
            .O(N__10839),
            .I(N__10703));
    SRMux I__2609 (
            .O(N__10838),
            .I(N__10703));
    SRMux I__2608 (
            .O(N__10837),
            .I(N__10703));
    SRMux I__2607 (
            .O(N__10836),
            .I(N__10703));
    Glb2LocalMux I__2606 (
            .O(N__10833),
            .I(N__10703));
    SRMux I__2605 (
            .O(N__10832),
            .I(N__10703));
    SRMux I__2604 (
            .O(N__10831),
            .I(N__10703));
    SRMux I__2603 (
            .O(N__10830),
            .I(N__10703));
    SRMux I__2602 (
            .O(N__10829),
            .I(N__10703));
    SRMux I__2601 (
            .O(N__10828),
            .I(N__10703));
    Glb2LocalMux I__2600 (
            .O(N__10825),
            .I(N__10703));
    SRMux I__2599 (
            .O(N__10824),
            .I(N__10703));
    SRMux I__2598 (
            .O(N__10823),
            .I(N__10703));
    SRMux I__2597 (
            .O(N__10822),
            .I(N__10703));
    SRMux I__2596 (
            .O(N__10821),
            .I(N__10703));
    SRMux I__2595 (
            .O(N__10820),
            .I(N__10703));
    SRMux I__2594 (
            .O(N__10819),
            .I(N__10703));
    Glb2LocalMux I__2593 (
            .O(N__10816),
            .I(N__10703));
    SRMux I__2592 (
            .O(N__10815),
            .I(N__10703));
    SRMux I__2591 (
            .O(N__10814),
            .I(N__10703));
    SRMux I__2590 (
            .O(N__10813),
            .I(N__10703));
    SRMux I__2589 (
            .O(N__10812),
            .I(N__10703));
    SRMux I__2588 (
            .O(N__10811),
            .I(N__10703));
    SRMux I__2587 (
            .O(N__10810),
            .I(N__10703));
    SRMux I__2586 (
            .O(N__10809),
            .I(N__10703));
    SRMux I__2585 (
            .O(N__10808),
            .I(N__10703));
    SRMux I__2584 (
            .O(N__10807),
            .I(N__10703));
    SRMux I__2583 (
            .O(N__10806),
            .I(N__10703));
    Glb2LocalMux I__2582 (
            .O(N__10803),
            .I(N__10703));
    SRMux I__2581 (
            .O(N__10802),
            .I(N__10703));
    SRMux I__2580 (
            .O(N__10801),
            .I(N__10703));
    SRMux I__2579 (
            .O(N__10800),
            .I(N__10703));
    SRMux I__2578 (
            .O(N__10799),
            .I(N__10703));
    SRMux I__2577 (
            .O(N__10798),
            .I(N__10703));
    GlobalMux I__2576 (
            .O(N__10703),
            .I(N__10700));
    gio2CtrlBuf I__2575 (
            .O(N__10700),
            .I(RESETn_c_i_g));
    CascadeMux I__2574 (
            .O(N__10697),
            .I(N__10694));
    InMux I__2573 (
            .O(N__10694),
            .I(N__10690));
    InMux I__2572 (
            .O(N__10693),
            .I(N__10687));
    LocalMux I__2571 (
            .O(N__10690),
            .I(N__10680));
    LocalMux I__2570 (
            .O(N__10687),
            .I(N__10680));
    InMux I__2569 (
            .O(N__10686),
            .I(N__10677));
    InMux I__2568 (
            .O(N__10685),
            .I(N__10674));
    Sp12to4 I__2567 (
            .O(N__10680),
            .I(N__10667));
    LocalMux I__2566 (
            .O(N__10677),
            .I(N__10667));
    LocalMux I__2565 (
            .O(N__10674),
            .I(N__10667));
    Span12Mux_v I__2564 (
            .O(N__10667),
            .I(N__10664));
    Span12Mux_h I__2563 (
            .O(N__10664),
            .I(N__10661));
    Odrv12 I__2562 (
            .O(N__10661),
            .I(DRA_c_6));
    InMux I__2561 (
            .O(N__10658),
            .I(N__10655));
    LocalMux I__2560 (
            .O(N__10655),
            .I(N__10652));
    Span4Mux_h I__2559 (
            .O(N__10652),
            .I(N__10649));
    Odrv4 I__2558 (
            .O(N__10649),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__2557 (
            .O(N__10646),
            .I(N__10643));
    LocalMux I__2556 (
            .O(N__10643),
            .I(N__10640));
    Span4Mux_h I__2555 (
            .O(N__10640),
            .I(N__10636));
    InMux I__2554 (
            .O(N__10639),
            .I(N__10633));
    Odrv4 I__2553 (
            .O(N__10636),
            .I(DBRn_c_i));
    LocalMux I__2552 (
            .O(N__10633),
            .I(DBRn_c_i));
    InMux I__2551 (
            .O(N__10628),
            .I(N__10624));
    InMux I__2550 (
            .O(N__10627),
            .I(N__10621));
    LocalMux I__2549 (
            .O(N__10624),
            .I(N__10618));
    LocalMux I__2548 (
            .O(N__10621),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    Odrv12 I__2547 (
            .O(N__10618),
            .I(\U712_CHIP_RAM.DMA_AZ0Z20 ));
    InMux I__2546 (
            .O(N__10613),
            .I(N__10610));
    LocalMux I__2545 (
            .O(N__10610),
            .I(N__10607));
    Span4Mux_h I__2544 (
            .O(N__10607),
            .I(N__10604));
    Odrv4 I__2543 (
            .O(N__10604),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__2542 (
            .O(N__10601),
            .I(N__10596));
    InMux I__2541 (
            .O(N__10600),
            .I(N__10593));
    InMux I__2540 (
            .O(N__10599),
            .I(N__10590));
    LocalMux I__2539 (
            .O(N__10596),
            .I(N__10587));
    LocalMux I__2538 (
            .O(N__10593),
            .I(N__10581));
    LocalMux I__2537 (
            .O(N__10590),
            .I(N__10581));
    Span4Mux_v I__2536 (
            .O(N__10587),
            .I(N__10578));
    CascadeMux I__2535 (
            .O(N__10586),
            .I(N__10575));
    Span4Mux_h I__2534 (
            .O(N__10581),
            .I(N__10572));
    Span4Mux_v I__2533 (
            .O(N__10578),
            .I(N__10569));
    InMux I__2532 (
            .O(N__10575),
            .I(N__10566));
    Span4Mux_v I__2531 (
            .O(N__10572),
            .I(N__10563));
    Sp12to4 I__2530 (
            .O(N__10569),
            .I(N__10558));
    LocalMux I__2529 (
            .O(N__10566),
            .I(N__10558));
    Sp12to4 I__2528 (
            .O(N__10563),
            .I(N__10555));
    Span12Mux_h I__2527 (
            .O(N__10558),
            .I(N__10552));
    Span12Mux_v I__2526 (
            .O(N__10555),
            .I(N__10549));
    Span12Mux_v I__2525 (
            .O(N__10552),
            .I(N__10546));
    Odrv12 I__2524 (
            .O(N__10549),
            .I(DRA_c_9));
    Odrv12 I__2523 (
            .O(N__10546),
            .I(DRA_c_9));
    InMux I__2522 (
            .O(N__10541),
            .I(N__10538));
    LocalMux I__2521 (
            .O(N__10538),
            .I(N__10535));
    Span4Mux_h I__2520 (
            .O(N__10535),
            .I(N__10532));
    Odrv4 I__2519 (
            .O(N__10532),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__2518 (
            .O(N__10529),
            .I(N__10523));
    InMux I__2517 (
            .O(N__10528),
            .I(N__10520));
    InMux I__2516 (
            .O(N__10527),
            .I(N__10517));
    InMux I__2515 (
            .O(N__10526),
            .I(N__10514));
    LocalMux I__2514 (
            .O(N__10523),
            .I(N__10511));
    LocalMux I__2513 (
            .O(N__10520),
            .I(N__10508));
    LocalMux I__2512 (
            .O(N__10517),
            .I(N__10503));
    LocalMux I__2511 (
            .O(N__10514),
            .I(N__10503));
    Span4Mux_v I__2510 (
            .O(N__10511),
            .I(N__10500));
    Span4Mux_v I__2509 (
            .O(N__10508),
            .I(N__10495));
    Span4Mux_v I__2508 (
            .O(N__10503),
            .I(N__10495));
    Sp12to4 I__2507 (
            .O(N__10500),
            .I(N__10492));
    Sp12to4 I__2506 (
            .O(N__10495),
            .I(N__10489));
    Span12Mux_h I__2505 (
            .O(N__10492),
            .I(N__10486));
    Span12Mux_h I__2504 (
            .O(N__10489),
            .I(N__10483));
    Odrv12 I__2503 (
            .O(N__10486),
            .I(DRA_c_7));
    Odrv12 I__2502 (
            .O(N__10483),
            .I(DRA_c_7));
    InMux I__2501 (
            .O(N__10478),
            .I(N__10473));
    InMux I__2500 (
            .O(N__10477),
            .I(N__10470));
    InMux I__2499 (
            .O(N__10476),
            .I(N__10467));
    LocalMux I__2498 (
            .O(N__10473),
            .I(N__10460));
    LocalMux I__2497 (
            .O(N__10470),
            .I(N__10460));
    LocalMux I__2496 (
            .O(N__10467),
            .I(N__10460));
    Span4Mux_v I__2495 (
            .O(N__10460),
            .I(N__10456));
    InMux I__2494 (
            .O(N__10459),
            .I(N__10453));
    Sp12to4 I__2493 (
            .O(N__10456),
            .I(N__10448));
    LocalMux I__2492 (
            .O(N__10453),
            .I(N__10448));
    Span12Mux_h I__2491 (
            .O(N__10448),
            .I(N__10445));
    Odrv12 I__2490 (
            .O(N__10445),
            .I(DRA_c_8));
    InMux I__2489 (
            .O(N__10442),
            .I(N__10439));
    LocalMux I__2488 (
            .O(N__10439),
            .I(N__10436));
    Span4Mux_h I__2487 (
            .O(N__10436),
            .I(N__10433));
    Span4Mux_h I__2486 (
            .O(N__10433),
            .I(N__10430));
    Odrv4 I__2485 (
            .O(N__10430),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__2484 (
            .O(N__10427),
            .I(N__10424));
    LocalMux I__2483 (
            .O(N__10424),
            .I(N__10421));
    Odrv12 I__2482 (
            .O(N__10421),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__2481 (
            .O(N__10418),
            .I(N__10415));
    LocalMux I__2480 (
            .O(N__10415),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__2479 (
            .O(N__10412),
            .I(N__10407));
    InMux I__2478 (
            .O(N__10411),
            .I(N__10404));
    InMux I__2477 (
            .O(N__10410),
            .I(N__10401));
    LocalMux I__2476 (
            .O(N__10407),
            .I(N__10397));
    LocalMux I__2475 (
            .O(N__10404),
            .I(N__10394));
    LocalMux I__2474 (
            .O(N__10401),
            .I(N__10391));
    InMux I__2473 (
            .O(N__10400),
            .I(N__10388));
    Span4Mux_v I__2472 (
            .O(N__10397),
            .I(N__10385));
    Span4Mux_v I__2471 (
            .O(N__10394),
            .I(N__10378));
    Span4Mux_h I__2470 (
            .O(N__10391),
            .I(N__10378));
    LocalMux I__2469 (
            .O(N__10388),
            .I(N__10378));
    Span4Mux_v I__2468 (
            .O(N__10385),
            .I(N__10375));
    Span4Mux_h I__2467 (
            .O(N__10378),
            .I(N__10372));
    Sp12to4 I__2466 (
            .O(N__10375),
            .I(N__10369));
    Sp12to4 I__2465 (
            .O(N__10372),
            .I(N__10366));
    Span12Mux_h I__2464 (
            .O(N__10369),
            .I(N__10363));
    Span12Mux_v I__2463 (
            .O(N__10366),
            .I(N__10360));
    Odrv12 I__2462 (
            .O(N__10363),
            .I(DRA_c_2));
    Odrv12 I__2461 (
            .O(N__10360),
            .I(DRA_c_2));
    InMux I__2460 (
            .O(N__10355),
            .I(N__10349));
    InMux I__2459 (
            .O(N__10354),
            .I(N__10349));
    LocalMux I__2458 (
            .O(N__10349),
            .I(N__10346));
    Span4Mux_h I__2457 (
            .O(N__10346),
            .I(N__10343));
    Odrv4 I__2456 (
            .O(N__10343),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    IoInMux I__2455 (
            .O(N__10340),
            .I(N__10337));
    LocalMux I__2454 (
            .O(N__10337),
            .I(N__10334));
    Span4Mux_s2_h I__2453 (
            .O(N__10334),
            .I(N__10331));
    Sp12to4 I__2452 (
            .O(N__10331),
            .I(N__10328));
    Span12Mux_s10_v I__2451 (
            .O(N__10328),
            .I(N__10325));
    Odrv12 I__2450 (
            .O(N__10325),
            .I(WEn_c));
    InMux I__2449 (
            .O(N__10322),
            .I(N__10318));
    InMux I__2448 (
            .O(N__10321),
            .I(N__10315));
    LocalMux I__2447 (
            .O(N__10318),
            .I(N__10312));
    LocalMux I__2446 (
            .O(N__10315),
            .I(N__10306));
    Span4Mux_h I__2445 (
            .O(N__10312),
            .I(N__10306));
    InMux I__2444 (
            .O(N__10311),
            .I(N__10303));
    Span4Mux_v I__2443 (
            .O(N__10306),
            .I(N__10296));
    LocalMux I__2442 (
            .O(N__10303),
            .I(N__10296));
    InMux I__2441 (
            .O(N__10302),
            .I(N__10291));
    InMux I__2440 (
            .O(N__10301),
            .I(N__10288));
    Span4Mux_h I__2439 (
            .O(N__10296),
            .I(N__10285));
    InMux I__2438 (
            .O(N__10295),
            .I(N__10280));
    InMux I__2437 (
            .O(N__10294),
            .I(N__10280));
    LocalMux I__2436 (
            .O(N__10291),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    LocalMux I__2435 (
            .O(N__10288),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv4 I__2434 (
            .O(N__10285),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    LocalMux I__2433 (
            .O(N__10280),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    CascadeMux I__2432 (
            .O(N__10271),
            .I(N__10268));
    InMux I__2431 (
            .O(N__10268),
            .I(N__10264));
    InMux I__2430 (
            .O(N__10267),
            .I(N__10261));
    LocalMux I__2429 (
            .O(N__10264),
            .I(N__10255));
    LocalMux I__2428 (
            .O(N__10261),
            .I(N__10255));
    InMux I__2427 (
            .O(N__10260),
            .I(N__10252));
    Span4Mux_v I__2426 (
            .O(N__10255),
            .I(N__10249));
    LocalMux I__2425 (
            .O(N__10252),
            .I(N__10242));
    Span4Mux_h I__2424 (
            .O(N__10249),
            .I(N__10242));
    InMux I__2423 (
            .O(N__10248),
            .I(N__10237));
    InMux I__2422 (
            .O(N__10247),
            .I(N__10237));
    Odrv4 I__2421 (
            .O(N__10242),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__2420 (
            .O(N__10237),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    InMux I__2419 (
            .O(N__10232),
            .I(N__10228));
    InMux I__2418 (
            .O(N__10231),
            .I(N__10225));
    LocalMux I__2417 (
            .O(N__10228),
            .I(N__10221));
    LocalMux I__2416 (
            .O(N__10225),
            .I(N__10218));
    CascadeMux I__2415 (
            .O(N__10224),
            .I(N__10212));
    Span4Mux_v I__2414 (
            .O(N__10221),
            .I(N__10206));
    Span4Mux_v I__2413 (
            .O(N__10218),
            .I(N__10206));
    InMux I__2412 (
            .O(N__10217),
            .I(N__10203));
    CascadeMux I__2411 (
            .O(N__10216),
            .I(N__10200));
    CascadeMux I__2410 (
            .O(N__10215),
            .I(N__10197));
    InMux I__2409 (
            .O(N__10212),
            .I(N__10194));
    InMux I__2408 (
            .O(N__10211),
            .I(N__10191));
    Span4Mux_h I__2407 (
            .O(N__10206),
            .I(N__10186));
    LocalMux I__2406 (
            .O(N__10203),
            .I(N__10186));
    InMux I__2405 (
            .O(N__10200),
            .I(N__10181));
    InMux I__2404 (
            .O(N__10197),
            .I(N__10181));
    LocalMux I__2403 (
            .O(N__10194),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    LocalMux I__2402 (
            .O(N__10191),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    Odrv4 I__2401 (
            .O(N__10186),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    LocalMux I__2400 (
            .O(N__10181),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    IoInMux I__2399 (
            .O(N__10172),
            .I(N__10169));
    LocalMux I__2398 (
            .O(N__10169),
            .I(N__10166));
    IoSpan4Mux I__2397 (
            .O(N__10166),
            .I(N__10163));
    Span4Mux_s1_v I__2396 (
            .O(N__10163),
            .I(N__10160));
    Sp12to4 I__2395 (
            .O(N__10160),
            .I(N__10157));
    Span12Mux_v I__2394 (
            .O(N__10157),
            .I(N__10154));
    Odrv12 I__2393 (
            .O(N__10154),
            .I(CMA_c_10));
    CascadeMux I__2392 (
            .O(N__10151),
            .I(N__10148));
    InMux I__2391 (
            .O(N__10148),
            .I(N__10145));
    LocalMux I__2390 (
            .O(N__10145),
            .I(N__10142));
    Span4Mux_v I__2389 (
            .O(N__10142),
            .I(N__10139));
    Odrv4 I__2388 (
            .O(N__10139),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__2387 (
            .O(N__10136),
            .I(N__10131));
    InMux I__2386 (
            .O(N__10135),
            .I(N__10126));
    InMux I__2385 (
            .O(N__10134),
            .I(N__10126));
    LocalMux I__2384 (
            .O(N__10131),
            .I(N__10120));
    LocalMux I__2383 (
            .O(N__10126),
            .I(N__10120));
    InMux I__2382 (
            .O(N__10125),
            .I(N__10117));
    Sp12to4 I__2381 (
            .O(N__10120),
            .I(N__10112));
    LocalMux I__2380 (
            .O(N__10117),
            .I(N__10112));
    Span12Mux_v I__2379 (
            .O(N__10112),
            .I(N__10109));
    Span12Mux_h I__2378 (
            .O(N__10109),
            .I(N__10106));
    Odrv12 I__2377 (
            .O(N__10106),
            .I(DRA_c_5));
    InMux I__2376 (
            .O(N__10103),
            .I(N__10099));
    InMux I__2375 (
            .O(N__10102),
            .I(N__10096));
    LocalMux I__2374 (
            .O(N__10099),
            .I(N__10093));
    LocalMux I__2373 (
            .O(N__10096),
            .I(N__10090));
    Span4Mux_h I__2372 (
            .O(N__10093),
            .I(N__10087));
    Odrv12 I__2371 (
            .O(N__10090),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    Odrv4 I__2370 (
            .O(N__10087),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__2369 (
            .O(N__10082),
            .I(N__10079));
    LocalMux I__2368 (
            .O(N__10079),
            .I(N__10076));
    Span12Mux_h I__2367 (
            .O(N__10076),
            .I(N__10073));
    Odrv12 I__2366 (
            .O(N__10073),
            .I(RAS0n_c));
    InMux I__2365 (
            .O(N__10070),
            .I(N__10067));
    LocalMux I__2364 (
            .O(N__10067),
            .I(N__10064));
    Span4Mux_h I__2363 (
            .O(N__10064),
            .I(N__10061));
    Odrv4 I__2362 (
            .O(N__10061),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    CascadeMux I__2361 (
            .O(N__10058),
            .I(N__10055));
    InMux I__2360 (
            .O(N__10055),
            .I(N__10045));
    InMux I__2359 (
            .O(N__10054),
            .I(N__10045));
    InMux I__2358 (
            .O(N__10053),
            .I(N__10040));
    InMux I__2357 (
            .O(N__10052),
            .I(N__10040));
    InMux I__2356 (
            .O(N__10051),
            .I(N__10037));
    InMux I__2355 (
            .O(N__10050),
            .I(N__10033));
    LocalMux I__2354 (
            .O(N__10045),
            .I(N__10028));
    LocalMux I__2353 (
            .O(N__10040),
            .I(N__10028));
    LocalMux I__2352 (
            .O(N__10037),
            .I(N__10025));
    InMux I__2351 (
            .O(N__10036),
            .I(N__10021));
    LocalMux I__2350 (
            .O(N__10033),
            .I(N__10018));
    Span4Mux_h I__2349 (
            .O(N__10028),
            .I(N__10015));
    Span4Mux_h I__2348 (
            .O(N__10025),
            .I(N__10012));
    InMux I__2347 (
            .O(N__10024),
            .I(N__10009));
    LocalMux I__2346 (
            .O(N__10021),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv12 I__2345 (
            .O(N__10018),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__2344 (
            .O(N__10015),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    Odrv4 I__2343 (
            .O(N__10012),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    LocalMux I__2342 (
            .O(N__10009),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ));
    CascadeMux I__2341 (
            .O(N__9998),
            .I(N__9992));
    CascadeMux I__2340 (
            .O(N__9997),
            .I(N__9989));
    CascadeMux I__2339 (
            .O(N__9996),
            .I(N__9984));
    CascadeMux I__2338 (
            .O(N__9995),
            .I(N__9981));
    InMux I__2337 (
            .O(N__9992),
            .I(N__9978));
    InMux I__2336 (
            .O(N__9989),
            .I(N__9975));
    InMux I__2335 (
            .O(N__9988),
            .I(N__9966));
    InMux I__2334 (
            .O(N__9987),
            .I(N__9966));
    InMux I__2333 (
            .O(N__9984),
            .I(N__9966));
    InMux I__2332 (
            .O(N__9981),
            .I(N__9966));
    LocalMux I__2331 (
            .O(N__9978),
            .I(N__9963));
    LocalMux I__2330 (
            .O(N__9975),
            .I(N__9960));
    LocalMux I__2329 (
            .O(N__9966),
            .I(N__9957));
    Span4Mux_h I__2328 (
            .O(N__9963),
            .I(N__9954));
    Odrv4 I__2327 (
            .O(N__9960),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    Odrv12 I__2326 (
            .O(N__9957),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    Odrv4 I__2325 (
            .O(N__9954),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    IoInMux I__2324 (
            .O(N__9947),
            .I(N__9944));
    LocalMux I__2323 (
            .O(N__9944),
            .I(N__9941));
    Span4Mux_s2_v I__2322 (
            .O(N__9941),
            .I(N__9938));
    Span4Mux_v I__2321 (
            .O(N__9938),
            .I(N__9935));
    Span4Mux_v I__2320 (
            .O(N__9935),
            .I(N__9932));
    Span4Mux_h I__2319 (
            .O(N__9932),
            .I(N__9929));
    Odrv4 I__2318 (
            .O(N__9929),
            .I(CMA_c_0));
    InMux I__2317 (
            .O(N__9926),
            .I(N__9923));
    LocalMux I__2316 (
            .O(N__9923),
            .I(N__9904));
    ClkMux I__2315 (
            .O(N__9922),
            .I(N__9842));
    ClkMux I__2314 (
            .O(N__9921),
            .I(N__9842));
    ClkMux I__2313 (
            .O(N__9920),
            .I(N__9842));
    ClkMux I__2312 (
            .O(N__9919),
            .I(N__9842));
    ClkMux I__2311 (
            .O(N__9918),
            .I(N__9842));
    ClkMux I__2310 (
            .O(N__9917),
            .I(N__9842));
    ClkMux I__2309 (
            .O(N__9916),
            .I(N__9842));
    ClkMux I__2308 (
            .O(N__9915),
            .I(N__9842));
    ClkMux I__2307 (
            .O(N__9914),
            .I(N__9842));
    ClkMux I__2306 (
            .O(N__9913),
            .I(N__9842));
    ClkMux I__2305 (
            .O(N__9912),
            .I(N__9842));
    ClkMux I__2304 (
            .O(N__9911),
            .I(N__9842));
    ClkMux I__2303 (
            .O(N__9910),
            .I(N__9842));
    ClkMux I__2302 (
            .O(N__9909),
            .I(N__9842));
    ClkMux I__2301 (
            .O(N__9908),
            .I(N__9842));
    ClkMux I__2300 (
            .O(N__9907),
            .I(N__9842));
    Glb2LocalMux I__2299 (
            .O(N__9904),
            .I(N__9842));
    ClkMux I__2298 (
            .O(N__9903),
            .I(N__9842));
    ClkMux I__2297 (
            .O(N__9902),
            .I(N__9842));
    ClkMux I__2296 (
            .O(N__9901),
            .I(N__9842));
    ClkMux I__2295 (
            .O(N__9900),
            .I(N__9842));
    ClkMux I__2294 (
            .O(N__9899),
            .I(N__9842));
    ClkMux I__2293 (
            .O(N__9898),
            .I(N__9842));
    ClkMux I__2292 (
            .O(N__9897),
            .I(N__9842));
    ClkMux I__2291 (
            .O(N__9896),
            .I(N__9842));
    ClkMux I__2290 (
            .O(N__9895),
            .I(N__9842));
    GlobalMux I__2289 (
            .O(N__9842),
            .I(CLK80_PLL));
    CEMux I__2288 (
            .O(N__9839),
            .I(N__9834));
    CEMux I__2287 (
            .O(N__9838),
            .I(N__9830));
    CEMux I__2286 (
            .O(N__9837),
            .I(N__9826));
    LocalMux I__2285 (
            .O(N__9834),
            .I(N__9823));
    CEMux I__2284 (
            .O(N__9833),
            .I(N__9820));
    LocalMux I__2283 (
            .O(N__9830),
            .I(N__9817));
    CEMux I__2282 (
            .O(N__9829),
            .I(N__9814));
    LocalMux I__2281 (
            .O(N__9826),
            .I(N__9811));
    Span4Mux_v I__2280 (
            .O(N__9823),
            .I(N__9808));
    LocalMux I__2279 (
            .O(N__9820),
            .I(N__9801));
    Span4Mux_h I__2278 (
            .O(N__9817),
            .I(N__9801));
    LocalMux I__2277 (
            .O(N__9814),
            .I(N__9801));
    Span4Mux_v I__2276 (
            .O(N__9811),
            .I(N__9798));
    Span4Mux_h I__2275 (
            .O(N__9808),
            .I(N__9793));
    Span4Mux_v I__2274 (
            .O(N__9801),
            .I(N__9793));
    Sp12to4 I__2273 (
            .O(N__9798),
            .I(N__9787));
    Sp12to4 I__2272 (
            .O(N__9793),
            .I(N__9787));
    CEMux I__2271 (
            .O(N__9792),
            .I(N__9784));
    Span12Mux_h I__2270 (
            .O(N__9787),
            .I(N__9779));
    LocalMux I__2269 (
            .O(N__9784),
            .I(N__9779));
    Odrv12 I__2268 (
            .O(N__9779),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i_0 ));
    InMux I__2267 (
            .O(N__9776),
            .I(N__9773));
    LocalMux I__2266 (
            .O(N__9773),
            .I(N__9770));
    Span12Mux_h I__2265 (
            .O(N__9770),
            .I(N__9767));
    Odrv12 I__2264 (
            .O(N__9767),
            .I(A_c_9));
    InMux I__2263 (
            .O(N__9764),
            .I(N__9761));
    LocalMux I__2262 (
            .O(N__9761),
            .I(N__9758));
    Span4Mux_v I__2261 (
            .O(N__9758),
            .I(N__9755));
    Sp12to4 I__2260 (
            .O(N__9755),
            .I(N__9752));
    Span12Mux_h I__2259 (
            .O(N__9752),
            .I(N__9749));
    Span12Mux_v I__2258 (
            .O(N__9749),
            .I(N__9746));
    Odrv12 I__2257 (
            .O(N__9746),
            .I(A_c_2));
    InMux I__2256 (
            .O(N__9743),
            .I(N__9737));
    InMux I__2255 (
            .O(N__9742),
            .I(N__9732));
    CascadeMux I__2254 (
            .O(N__9741),
            .I(N__9728));
    CascadeMux I__2253 (
            .O(N__9740),
            .I(N__9720));
    LocalMux I__2252 (
            .O(N__9737),
            .I(N__9711));
    InMux I__2251 (
            .O(N__9736),
            .I(N__9704));
    InMux I__2250 (
            .O(N__9735),
            .I(N__9704));
    LocalMux I__2249 (
            .O(N__9732),
            .I(N__9699));
    InMux I__2248 (
            .O(N__9731),
            .I(N__9696));
    InMux I__2247 (
            .O(N__9728),
            .I(N__9693));
    InMux I__2246 (
            .O(N__9727),
            .I(N__9690));
    InMux I__2245 (
            .O(N__9726),
            .I(N__9681));
    InMux I__2244 (
            .O(N__9725),
            .I(N__9681));
    InMux I__2243 (
            .O(N__9724),
            .I(N__9681));
    InMux I__2242 (
            .O(N__9723),
            .I(N__9681));
    InMux I__2241 (
            .O(N__9720),
            .I(N__9678));
    InMux I__2240 (
            .O(N__9719),
            .I(N__9671));
    InMux I__2239 (
            .O(N__9718),
            .I(N__9671));
    InMux I__2238 (
            .O(N__9717),
            .I(N__9671));
    InMux I__2237 (
            .O(N__9716),
            .I(N__9666));
    InMux I__2236 (
            .O(N__9715),
            .I(N__9666));
    InMux I__2235 (
            .O(N__9714),
            .I(N__9661));
    Span12Mux_v I__2234 (
            .O(N__9711),
            .I(N__9658));
    InMux I__2233 (
            .O(N__9710),
            .I(N__9653));
    InMux I__2232 (
            .O(N__9709),
            .I(N__9653));
    LocalMux I__2231 (
            .O(N__9704),
            .I(N__9650));
    InMux I__2230 (
            .O(N__9703),
            .I(N__9645));
    InMux I__2229 (
            .O(N__9702),
            .I(N__9645));
    Span4Mux_v I__2228 (
            .O(N__9699),
            .I(N__9640));
    LocalMux I__2227 (
            .O(N__9696),
            .I(N__9640));
    LocalMux I__2226 (
            .O(N__9693),
            .I(N__9633));
    LocalMux I__2225 (
            .O(N__9690),
            .I(N__9633));
    LocalMux I__2224 (
            .O(N__9681),
            .I(N__9633));
    LocalMux I__2223 (
            .O(N__9678),
            .I(N__9626));
    LocalMux I__2222 (
            .O(N__9671),
            .I(N__9626));
    LocalMux I__2221 (
            .O(N__9666),
            .I(N__9626));
    InMux I__2220 (
            .O(N__9665),
            .I(N__9621));
    InMux I__2219 (
            .O(N__9664),
            .I(N__9621));
    LocalMux I__2218 (
            .O(N__9661),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__2217 (
            .O(N__9658),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2216 (
            .O(N__9653),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv12 I__2215 (
            .O(N__9650),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2214 (
            .O(N__9645),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2213 (
            .O(N__9640),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2212 (
            .O(N__9633),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__2211 (
            .O(N__9626),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__2210 (
            .O(N__9621),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    CascadeMux I__2209 (
            .O(N__9602),
            .I(N__9599));
    InMux I__2208 (
            .O(N__9599),
            .I(N__9594));
    CascadeMux I__2207 (
            .O(N__9598),
            .I(N__9585));
    CascadeMux I__2206 (
            .O(N__9597),
            .I(N__9578));
    LocalMux I__2205 (
            .O(N__9594),
            .I(N__9572));
    InMux I__2204 (
            .O(N__9593),
            .I(N__9569));
    InMux I__2203 (
            .O(N__9592),
            .I(N__9563));
    InMux I__2202 (
            .O(N__9591),
            .I(N__9560));
    InMux I__2201 (
            .O(N__9590),
            .I(N__9557));
    InMux I__2200 (
            .O(N__9589),
            .I(N__9554));
    InMux I__2199 (
            .O(N__9588),
            .I(N__9551));
    InMux I__2198 (
            .O(N__9585),
            .I(N__9548));
    InMux I__2197 (
            .O(N__9584),
            .I(N__9541));
    InMux I__2196 (
            .O(N__9583),
            .I(N__9541));
    InMux I__2195 (
            .O(N__9582),
            .I(N__9541));
    InMux I__2194 (
            .O(N__9581),
            .I(N__9536));
    InMux I__2193 (
            .O(N__9578),
            .I(N__9536));
    InMux I__2192 (
            .O(N__9577),
            .I(N__9529));
    InMux I__2191 (
            .O(N__9576),
            .I(N__9529));
    InMux I__2190 (
            .O(N__9575),
            .I(N__9529));
    Span4Mux_h I__2189 (
            .O(N__9572),
            .I(N__9524));
    LocalMux I__2188 (
            .O(N__9569),
            .I(N__9524));
    InMux I__2187 (
            .O(N__9568),
            .I(N__9521));
    InMux I__2186 (
            .O(N__9567),
            .I(N__9514));
    InMux I__2185 (
            .O(N__9566),
            .I(N__9514));
    LocalMux I__2184 (
            .O(N__9563),
            .I(N__9507));
    LocalMux I__2183 (
            .O(N__9560),
            .I(N__9507));
    LocalMux I__2182 (
            .O(N__9557),
            .I(N__9507));
    LocalMux I__2181 (
            .O(N__9554),
            .I(N__9496));
    LocalMux I__2180 (
            .O(N__9551),
            .I(N__9496));
    LocalMux I__2179 (
            .O(N__9548),
            .I(N__9496));
    LocalMux I__2178 (
            .O(N__9541),
            .I(N__9496));
    LocalMux I__2177 (
            .O(N__9536),
            .I(N__9496));
    LocalMux I__2176 (
            .O(N__9529),
            .I(N__9492));
    Span4Mux_v I__2175 (
            .O(N__9524),
            .I(N__9487));
    LocalMux I__2174 (
            .O(N__9521),
            .I(N__9487));
    InMux I__2173 (
            .O(N__9520),
            .I(N__9484));
    InMux I__2172 (
            .O(N__9519),
            .I(N__9480));
    LocalMux I__2171 (
            .O(N__9514),
            .I(N__9473));
    Span4Mux_h I__2170 (
            .O(N__9507),
            .I(N__9473));
    Span4Mux_v I__2169 (
            .O(N__9496),
            .I(N__9473));
    InMux I__2168 (
            .O(N__9495),
            .I(N__9470));
    Span4Mux_v I__2167 (
            .O(N__9492),
            .I(N__9463));
    Span4Mux_h I__2166 (
            .O(N__9487),
            .I(N__9463));
    LocalMux I__2165 (
            .O(N__9484),
            .I(N__9463));
    InMux I__2164 (
            .O(N__9483),
            .I(N__9460));
    LocalMux I__2163 (
            .O(N__9480),
            .I(N__9457));
    Span4Mux_v I__2162 (
            .O(N__9473),
            .I(N__9454));
    LocalMux I__2161 (
            .O(N__9470),
            .I(N__9449));
    Span4Mux_h I__2160 (
            .O(N__9463),
            .I(N__9449));
    LocalMux I__2159 (
            .O(N__9460),
            .I(CPU_CYCLE));
    Odrv12 I__2158 (
            .O(N__9457),
            .I(CPU_CYCLE));
    Odrv4 I__2157 (
            .O(N__9454),
            .I(CPU_CYCLE));
    Odrv4 I__2156 (
            .O(N__9449),
            .I(CPU_CYCLE));
    CascadeMux I__2155 (
            .O(N__9440),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ));
    InMux I__2154 (
            .O(N__9437),
            .I(N__9434));
    LocalMux I__2153 (
            .O(N__9434),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    InMux I__2152 (
            .O(N__9431),
            .I(N__9428));
    LocalMux I__2151 (
            .O(N__9428),
            .I(N__9425));
    Odrv4 I__2150 (
            .O(N__9425),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2149 (
            .O(N__9422),
            .I(N__9418));
    InMux I__2148 (
            .O(N__9421),
            .I(N__9415));
    LocalMux I__2147 (
            .O(N__9418),
            .I(N__9408));
    LocalMux I__2146 (
            .O(N__9415),
            .I(N__9408));
    InMux I__2145 (
            .O(N__9414),
            .I(N__9405));
    InMux I__2144 (
            .O(N__9413),
            .I(N__9402));
    Span4Mux_h I__2143 (
            .O(N__9408),
            .I(N__9395));
    LocalMux I__2142 (
            .O(N__9405),
            .I(N__9395));
    LocalMux I__2141 (
            .O(N__9402),
            .I(N__9395));
    Span4Mux_v I__2140 (
            .O(N__9395),
            .I(N__9392));
    Span4Mux_v I__2139 (
            .O(N__9392),
            .I(N__9389));
    Sp12to4 I__2138 (
            .O(N__9389),
            .I(N__9386));
    Span12Mux_h I__2137 (
            .O(N__9386),
            .I(N__9383));
    Odrv12 I__2136 (
            .O(N__9383),
            .I(DRA_c_4));
    InMux I__2135 (
            .O(N__9380),
            .I(N__9377));
    LocalMux I__2134 (
            .O(N__9377),
            .I(N__9374));
    Span4Mux_v I__2133 (
            .O(N__9374),
            .I(N__9371));
    Odrv4 I__2132 (
            .O(N__9371),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2131 (
            .O(N__9368),
            .I(N__9364));
    InMux I__2130 (
            .O(N__9367),
            .I(N__9361));
    LocalMux I__2129 (
            .O(N__9364),
            .I(N__9356));
    LocalMux I__2128 (
            .O(N__9361),
            .I(N__9353));
    InMux I__2127 (
            .O(N__9360),
            .I(N__9350));
    InMux I__2126 (
            .O(N__9359),
            .I(N__9347));
    Span4Mux_v I__2125 (
            .O(N__9356),
            .I(N__9338));
    Span4Mux_h I__2124 (
            .O(N__9353),
            .I(N__9338));
    LocalMux I__2123 (
            .O(N__9350),
            .I(N__9338));
    LocalMux I__2122 (
            .O(N__9347),
            .I(N__9338));
    Sp12to4 I__2121 (
            .O(N__9338),
            .I(N__9335));
    Span12Mux_v I__2120 (
            .O(N__9335),
            .I(N__9332));
    Span12Mux_h I__2119 (
            .O(N__9332),
            .I(N__9329));
    Odrv12 I__2118 (
            .O(N__9329),
            .I(DRA_c_3));
    InMux I__2117 (
            .O(N__9326),
            .I(N__9323));
    LocalMux I__2116 (
            .O(N__9323),
            .I(N__9320));
    Span4Mux_v I__2115 (
            .O(N__9320),
            .I(N__9317));
    Odrv4 I__2114 (
            .O(N__9317),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    IoInMux I__2113 (
            .O(N__9314),
            .I(N__9311));
    LocalMux I__2112 (
            .O(N__9311),
            .I(N__9308));
    Span4Mux_s2_v I__2111 (
            .O(N__9308),
            .I(N__9305));
    Span4Mux_v I__2110 (
            .O(N__9305),
            .I(N__9302));
    Odrv4 I__2109 (
            .O(N__9302),
            .I(N_276_i));
    IoInMux I__2108 (
            .O(N__9299),
            .I(N__9296));
    LocalMux I__2107 (
            .O(N__9296),
            .I(N__9293));
    Span4Mux_s2_v I__2106 (
            .O(N__9293),
            .I(N__9290));
    Span4Mux_v I__2105 (
            .O(N__9290),
            .I(N__9287));
    Odrv4 I__2104 (
            .O(N__9287),
            .I(N_278_i));
    InMux I__2103 (
            .O(N__9284),
            .I(N__9275));
    InMux I__2102 (
            .O(N__9283),
            .I(N__9275));
    InMux I__2101 (
            .O(N__9282),
            .I(N__9275));
    LocalMux I__2100 (
            .O(N__9275),
            .I(N__9268));
    InMux I__2099 (
            .O(N__9274),
            .I(N__9265));
    InMux I__2098 (
            .O(N__9273),
            .I(N__9262));
    InMux I__2097 (
            .O(N__9272),
            .I(N__9255));
    InMux I__2096 (
            .O(N__9271),
            .I(N__9255));
    Span4Mux_v I__2095 (
            .O(N__9268),
            .I(N__9250));
    LocalMux I__2094 (
            .O(N__9265),
            .I(N__9250));
    LocalMux I__2093 (
            .O(N__9262),
            .I(N__9247));
    InMux I__2092 (
            .O(N__9261),
            .I(N__9242));
    InMux I__2091 (
            .O(N__9260),
            .I(N__9239));
    LocalMux I__2090 (
            .O(N__9255),
            .I(N__9236));
    Span4Mux_h I__2089 (
            .O(N__9250),
            .I(N__9233));
    Span4Mux_v I__2088 (
            .O(N__9247),
            .I(N__9230));
    InMux I__2087 (
            .O(N__9246),
            .I(N__9227));
    InMux I__2086 (
            .O(N__9245),
            .I(N__9224));
    LocalMux I__2085 (
            .O(N__9242),
            .I(N__9221));
    LocalMux I__2084 (
            .O(N__9239),
            .I(N__9218));
    Span12Mux_v I__2083 (
            .O(N__9236),
            .I(N__9215));
    Span4Mux_v I__2082 (
            .O(N__9233),
            .I(N__9210));
    Span4Mux_v I__2081 (
            .O(N__9230),
            .I(N__9210));
    LocalMux I__2080 (
            .O(N__9227),
            .I(N__9205));
    LocalMux I__2079 (
            .O(N__9224),
            .I(N__9205));
    Span4Mux_v I__2078 (
            .O(N__9221),
            .I(N__9200));
    Span4Mux_v I__2077 (
            .O(N__9218),
            .I(N__9200));
    Span12Mux_h I__2076 (
            .O(N__9215),
            .I(N__9197));
    Sp12to4 I__2075 (
            .O(N__9210),
            .I(N__9190));
    Span12Mux_v I__2074 (
            .O(N__9205),
            .I(N__9190));
    Sp12to4 I__2073 (
            .O(N__9200),
            .I(N__9190));
    Odrv12 I__2072 (
            .O(N__9197),
            .I(A_c_0));
    Odrv12 I__2071 (
            .O(N__9190),
            .I(A_c_0));
    CascadeMux I__2070 (
            .O(N__9185),
            .I(N__9181));
    InMux I__2069 (
            .O(N__9184),
            .I(N__9174));
    InMux I__2068 (
            .O(N__9181),
            .I(N__9171));
    InMux I__2067 (
            .O(N__9180),
            .I(N__9168));
    InMux I__2066 (
            .O(N__9179),
            .I(N__9160));
    InMux I__2065 (
            .O(N__9178),
            .I(N__9160));
    InMux I__2064 (
            .O(N__9177),
            .I(N__9160));
    LocalMux I__2063 (
            .O(N__9174),
            .I(N__9157));
    LocalMux I__2062 (
            .O(N__9171),
            .I(N__9152));
    LocalMux I__2061 (
            .O(N__9168),
            .I(N__9152));
    CascadeMux I__2060 (
            .O(N__9167),
            .I(N__9149));
    LocalMux I__2059 (
            .O(N__9160),
            .I(N__9146));
    Span4Mux_v I__2058 (
            .O(N__9157),
            .I(N__9143));
    Span4Mux_v I__2057 (
            .O(N__9152),
            .I(N__9140));
    InMux I__2056 (
            .O(N__9149),
            .I(N__9137));
    Span4Mux_h I__2055 (
            .O(N__9146),
            .I(N__9134));
    Sp12to4 I__2054 (
            .O(N__9143),
            .I(N__9127));
    Sp12to4 I__2053 (
            .O(N__9140),
            .I(N__9127));
    LocalMux I__2052 (
            .O(N__9137),
            .I(N__9127));
    Span4Mux_v I__2051 (
            .O(N__9134),
            .I(N__9124));
    Span12Mux_h I__2050 (
            .O(N__9127),
            .I(N__9121));
    Sp12to4 I__2049 (
            .O(N__9124),
            .I(N__9118));
    Span12Mux_v I__2048 (
            .O(N__9121),
            .I(N__9113));
    Span12Mux_h I__2047 (
            .O(N__9118),
            .I(N__9113));
    Odrv12 I__2046 (
            .O(N__9113),
            .I(SIZ_c_0));
    InMux I__2045 (
            .O(N__9110),
            .I(N__9105));
    CascadeMux I__2044 (
            .O(N__9109),
            .I(N__9101));
    CascadeMux I__2043 (
            .O(N__9108),
            .I(N__9098));
    LocalMux I__2042 (
            .O(N__9105),
            .I(N__9095));
    InMux I__2041 (
            .O(N__9104),
            .I(N__9085));
    InMux I__2040 (
            .O(N__9101),
            .I(N__9085));
    InMux I__2039 (
            .O(N__9098),
            .I(N__9085));
    Span4Mux_v I__2038 (
            .O(N__9095),
            .I(N__9081));
    CascadeMux I__2037 (
            .O(N__9094),
            .I(N__9078));
    InMux I__2036 (
            .O(N__9093),
            .I(N__9073));
    InMux I__2035 (
            .O(N__9092),
            .I(N__9073));
    LocalMux I__2034 (
            .O(N__9085),
            .I(N__9070));
    InMux I__2033 (
            .O(N__9084),
            .I(N__9067));
    Span4Mux_v I__2032 (
            .O(N__9081),
            .I(N__9064));
    InMux I__2031 (
            .O(N__9078),
            .I(N__9061));
    LocalMux I__2030 (
            .O(N__9073),
            .I(N__9058));
    Span4Mux_v I__2029 (
            .O(N__9070),
            .I(N__9055));
    LocalMux I__2028 (
            .O(N__9067),
            .I(N__9052));
    Span4Mux_v I__2027 (
            .O(N__9064),
            .I(N__9049));
    LocalMux I__2026 (
            .O(N__9061),
            .I(N__9046));
    Span12Mux_v I__2025 (
            .O(N__9058),
            .I(N__9039));
    Sp12to4 I__2024 (
            .O(N__9055),
            .I(N__9039));
    Span12Mux_s7_v I__2023 (
            .O(N__9052),
            .I(N__9039));
    Sp12to4 I__2022 (
            .O(N__9049),
            .I(N__9034));
    Span12Mux_v I__2021 (
            .O(N__9046),
            .I(N__9034));
    Span12Mux_h I__2020 (
            .O(N__9039),
            .I(N__9031));
    Odrv12 I__2019 (
            .O(N__9034),
            .I(A_c_1));
    Odrv12 I__2018 (
            .O(N__9031),
            .I(A_c_1));
    CascadeMux I__2017 (
            .O(N__9026),
            .I(N__9023));
    InMux I__2016 (
            .O(N__9023),
            .I(N__9017));
    InMux I__2015 (
            .O(N__9022),
            .I(N__9014));
    InMux I__2014 (
            .O(N__9021),
            .I(N__9011));
    CascadeMux I__2013 (
            .O(N__9020),
            .I(N__9008));
    LocalMux I__2012 (
            .O(N__9017),
            .I(N__9003));
    LocalMux I__2011 (
            .O(N__9014),
            .I(N__8998));
    LocalMux I__2010 (
            .O(N__9011),
            .I(N__8998));
    InMux I__2009 (
            .O(N__9008),
            .I(N__8990));
    InMux I__2008 (
            .O(N__9007),
            .I(N__8990));
    InMux I__2007 (
            .O(N__9006),
            .I(N__8990));
    Span4Mux_v I__2006 (
            .O(N__9003),
            .I(N__8987));
    Span4Mux_v I__2005 (
            .O(N__8998),
            .I(N__8984));
    InMux I__2004 (
            .O(N__8997),
            .I(N__8981));
    LocalMux I__2003 (
            .O(N__8990),
            .I(N__8978));
    Sp12to4 I__2002 (
            .O(N__8987),
            .I(N__8971));
    Sp12to4 I__2001 (
            .O(N__8984),
            .I(N__8971));
    LocalMux I__2000 (
            .O(N__8981),
            .I(N__8971));
    Sp12to4 I__1999 (
            .O(N__8978),
            .I(N__8968));
    Span12Mux_h I__1998 (
            .O(N__8971),
            .I(N__8965));
    Span12Mux_v I__1997 (
            .O(N__8968),
            .I(N__8962));
    Span12Mux_v I__1996 (
            .O(N__8965),
            .I(N__8957));
    Span12Mux_h I__1995 (
            .O(N__8962),
            .I(N__8957));
    Odrv12 I__1994 (
            .O(N__8957),
            .I(SIZ_c_1));
    IoInMux I__1993 (
            .O(N__8954),
            .I(N__8951));
    LocalMux I__1992 (
            .O(N__8951),
            .I(N__8948));
    Span4Mux_s2_v I__1991 (
            .O(N__8948),
            .I(N__8945));
    Span4Mux_h I__1990 (
            .O(N__8945),
            .I(N__8942));
    Span4Mux_v I__1989 (
            .O(N__8942),
            .I(N__8939));
    Odrv4 I__1988 (
            .O(N__8939),
            .I(N_277_i));
    IoInMux I__1987 (
            .O(N__8936),
            .I(N__8933));
    LocalMux I__1986 (
            .O(N__8933),
            .I(N__8930));
    IoSpan4Mux I__1985 (
            .O(N__8930),
            .I(N__8927));
    Sp12to4 I__1984 (
            .O(N__8927),
            .I(N__8924));
    Span12Mux_s9_v I__1983 (
            .O(N__8924),
            .I(N__8921));
    Odrv12 I__1982 (
            .O(N__8921),
            .I(CRCSn_c));
    IoInMux I__1981 (
            .O(N__8918),
            .I(N__8915));
    LocalMux I__1980 (
            .O(N__8915),
            .I(N__8912));
    Span4Mux_s1_v I__1979 (
            .O(N__8912),
            .I(N__8909));
    Span4Mux_v I__1978 (
            .O(N__8909),
            .I(N__8906));
    Span4Mux_v I__1977 (
            .O(N__8906),
            .I(N__8903));
    Sp12to4 I__1976 (
            .O(N__8903),
            .I(N__8900));
    Odrv12 I__1975 (
            .O(N__8900),
            .I(RASn_c));
    IoInMux I__1974 (
            .O(N__8897),
            .I(N__8894));
    LocalMux I__1973 (
            .O(N__8894),
            .I(N__8891));
    Span4Mux_s1_v I__1972 (
            .O(N__8891),
            .I(N__8888));
    Sp12to4 I__1971 (
            .O(N__8888),
            .I(N__8885));
    Span12Mux_h I__1970 (
            .O(N__8885),
            .I(N__8882));
    Odrv12 I__1969 (
            .O(N__8882),
            .I(CASn_c));
    InMux I__1968 (
            .O(N__8879),
            .I(N__8875));
    InMux I__1967 (
            .O(N__8878),
            .I(N__8872));
    LocalMux I__1966 (
            .O(N__8875),
            .I(N__8866));
    LocalMux I__1965 (
            .O(N__8872),
            .I(N__8858));
    ClkMux I__1964 (
            .O(N__8871),
            .I(N__8837));
    ClkMux I__1963 (
            .O(N__8870),
            .I(N__8837));
    ClkMux I__1962 (
            .O(N__8869),
            .I(N__8837));
    Glb2LocalMux I__1961 (
            .O(N__8866),
            .I(N__8837));
    ClkMux I__1960 (
            .O(N__8865),
            .I(N__8837));
    ClkMux I__1959 (
            .O(N__8864),
            .I(N__8837));
    ClkMux I__1958 (
            .O(N__8863),
            .I(N__8837));
    ClkMux I__1957 (
            .O(N__8862),
            .I(N__8837));
    ClkMux I__1956 (
            .O(N__8861),
            .I(N__8837));
    Glb2LocalMux I__1955 (
            .O(N__8858),
            .I(N__8837));
    GlobalMux I__1954 (
            .O(N__8837),
            .I(N__8834));
    gio2CtrlBuf I__1953 (
            .O(N__8834),
            .I(CLK40_PLL_g));
    IoInMux I__1952 (
            .O(N__8831),
            .I(N__8828));
    LocalMux I__1951 (
            .O(N__8828),
            .I(N__8824));
    IoInMux I__1950 (
            .O(N__8827),
            .I(N__8821));
    IoSpan4Mux I__1949 (
            .O(N__8824),
            .I(N__8817));
    LocalMux I__1948 (
            .O(N__8821),
            .I(N__8814));
    IoInMux I__1947 (
            .O(N__8820),
            .I(N__8811));
    IoSpan4Mux I__1946 (
            .O(N__8817),
            .I(N__8808));
    Span4Mux_s3_v I__1945 (
            .O(N__8814),
            .I(N__8805));
    LocalMux I__1944 (
            .O(N__8811),
            .I(N__8802));
    Span4Mux_s3_v I__1943 (
            .O(N__8808),
            .I(N__8797));
    Span4Mux_h I__1942 (
            .O(N__8805),
            .I(N__8797));
    Span12Mux_s3_h I__1941 (
            .O(N__8802),
            .I(N__8794));
    Span4Mux_h I__1940 (
            .O(N__8797),
            .I(N__8791));
    Span12Mux_h I__1939 (
            .O(N__8794),
            .I(N__8788));
    Span4Mux_h I__1938 (
            .O(N__8791),
            .I(N__8785));
    Odrv12 I__1937 (
            .O(N__8788),
            .I(CLK40_PLL_iso_i));
    Odrv4 I__1936 (
            .O(N__8785),
            .I(CLK40_PLL_iso_i));
    IoInMux I__1935 (
            .O(N__8780),
            .I(N__8777));
    LocalMux I__1934 (
            .O(N__8777),
            .I(N__8774));
    IoSpan4Mux I__1933 (
            .O(N__8774),
            .I(N__8771));
    Span4Mux_s3_v I__1932 (
            .O(N__8771),
            .I(N__8768));
    Odrv4 I__1931 (
            .O(N__8768),
            .I(U712_BYTE_ENABLE_UUBE_i));
    InMux I__1930 (
            .O(N__8765),
            .I(N__8761));
    CascadeMux I__1929 (
            .O(N__8764),
            .I(N__8758));
    LocalMux I__1928 (
            .O(N__8761),
            .I(N__8755));
    InMux I__1927 (
            .O(N__8758),
            .I(N__8751));
    Span4Mux_h I__1926 (
            .O(N__8755),
            .I(N__8748));
    InMux I__1925 (
            .O(N__8754),
            .I(N__8745));
    LocalMux I__1924 (
            .O(N__8751),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    Odrv4 I__1923 (
            .O(N__8748),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    LocalMux I__1922 (
            .O(N__8745),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    InMux I__1921 (
            .O(N__8738),
            .I(N__8735));
    LocalMux I__1920 (
            .O(N__8735),
            .I(N__8732));
    Span4Mux_v I__1919 (
            .O(N__8732),
            .I(N__8729));
    Span4Mux_v I__1918 (
            .O(N__8729),
            .I(N__8726));
    Sp12to4 I__1917 (
            .O(N__8726),
            .I(N__8723));
    Span12Mux_h I__1916 (
            .O(N__8723),
            .I(N__8720));
    Odrv12 I__1915 (
            .O(N__8720),
            .I(A_c_17));
    IoInMux I__1914 (
            .O(N__8717),
            .I(N__8714));
    LocalMux I__1913 (
            .O(N__8714),
            .I(N__8711));
    Span12Mux_s3_h I__1912 (
            .O(N__8711),
            .I(N__8708));
    Span12Mux_h I__1911 (
            .O(N__8708),
            .I(N__8705));
    Odrv12 I__1910 (
            .O(N__8705),
            .I(CMA_c_8));
    InMux I__1909 (
            .O(N__8702),
            .I(N__8699));
    LocalMux I__1908 (
            .O(N__8699),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__1907 (
            .O(N__8696),
            .I(N__8693));
    LocalMux I__1906 (
            .O(N__8693),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__1905 (
            .O(N__8690),
            .I(N__8687));
    LocalMux I__1904 (
            .O(N__8687),
            .I(N__8684));
    Span4Mux_v I__1903 (
            .O(N__8684),
            .I(N__8681));
    Odrv4 I__1902 (
            .O(N__8681),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1901 (
            .O(N__8678),
            .I(N__8675));
    LocalMux I__1900 (
            .O(N__8675),
            .I(N__8672));
    Span4Mux_v I__1899 (
            .O(N__8672),
            .I(N__8669));
    Odrv4 I__1898 (
            .O(N__8669),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__1897 (
            .O(N__8666),
            .I(N__8663));
    LocalMux I__1896 (
            .O(N__8663),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__1895 (
            .O(N__8660),
            .I(N__8657));
    LocalMux I__1894 (
            .O(N__8657),
            .I(N__8654));
    Span4Mux_h I__1893 (
            .O(N__8654),
            .I(N__8651));
    Odrv4 I__1892 (
            .O(N__8651),
            .I(\U712_CHIP_RAM.N_456 ));
    InMux I__1891 (
            .O(N__8648),
            .I(N__8645));
    LocalMux I__1890 (
            .O(N__8645),
            .I(N__8642));
    Odrv4 I__1889 (
            .O(N__8642),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    CascadeMux I__1888 (
            .O(N__8639),
            .I(N__8636));
    InMux I__1887 (
            .O(N__8636),
            .I(N__8631));
    CascadeMux I__1886 (
            .O(N__8635),
            .I(N__8625));
    CascadeMux I__1885 (
            .O(N__8634),
            .I(N__8620));
    LocalMux I__1884 (
            .O(N__8631),
            .I(N__8617));
    InMux I__1883 (
            .O(N__8630),
            .I(N__8608));
    InMux I__1882 (
            .O(N__8629),
            .I(N__8608));
    InMux I__1881 (
            .O(N__8628),
            .I(N__8608));
    InMux I__1880 (
            .O(N__8625),
            .I(N__8608));
    InMux I__1879 (
            .O(N__8624),
            .I(N__8601));
    InMux I__1878 (
            .O(N__8623),
            .I(N__8601));
    InMux I__1877 (
            .O(N__8620),
            .I(N__8601));
    Odrv4 I__1876 (
            .O(N__8617),
            .I(\U712_CHIP_RAM.N_202 ));
    LocalMux I__1875 (
            .O(N__8608),
            .I(\U712_CHIP_RAM.N_202 ));
    LocalMux I__1874 (
            .O(N__8601),
            .I(\U712_CHIP_RAM.N_202 ));
    InMux I__1873 (
            .O(N__8594),
            .I(N__8591));
    LocalMux I__1872 (
            .O(N__8591),
            .I(N__8588));
    Span4Mux_h I__1871 (
            .O(N__8588),
            .I(N__8585));
    Odrv4 I__1870 (
            .O(N__8585),
            .I(\U712_CHIP_RAM.N_359 ));
    InMux I__1869 (
            .O(N__8582),
            .I(N__8575));
    InMux I__1868 (
            .O(N__8581),
            .I(N__8572));
    InMux I__1867 (
            .O(N__8580),
            .I(N__8569));
    InMux I__1866 (
            .O(N__8579),
            .I(N__8566));
    InMux I__1865 (
            .O(N__8578),
            .I(N__8563));
    LocalMux I__1864 (
            .O(N__8575),
            .I(N__8548));
    LocalMux I__1863 (
            .O(N__8572),
            .I(N__8548));
    LocalMux I__1862 (
            .O(N__8569),
            .I(N__8548));
    LocalMux I__1861 (
            .O(N__8566),
            .I(N__8548));
    LocalMux I__1860 (
            .O(N__8563),
            .I(N__8545));
    InMux I__1859 (
            .O(N__8562),
            .I(N__8542));
    InMux I__1858 (
            .O(N__8561),
            .I(N__8539));
    InMux I__1857 (
            .O(N__8560),
            .I(N__8534));
    InMux I__1856 (
            .O(N__8559),
            .I(N__8534));
    InMux I__1855 (
            .O(N__8558),
            .I(N__8529));
    InMux I__1854 (
            .O(N__8557),
            .I(N__8529));
    Span4Mux_h I__1853 (
            .O(N__8548),
            .I(N__8526));
    Odrv4 I__1852 (
            .O(N__8545),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1851 (
            .O(N__8542),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1850 (
            .O(N__8539),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1849 (
            .O(N__8534),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1848 (
            .O(N__8529),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1847 (
            .O(N__8526),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    CEMux I__1846 (
            .O(N__8513),
            .I(N__8510));
    LocalMux I__1845 (
            .O(N__8510),
            .I(N__8506));
    CEMux I__1844 (
            .O(N__8509),
            .I(N__8503));
    Odrv4 I__1843 (
            .O(N__8506),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    LocalMux I__1842 (
            .O(N__8503),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__1841 (
            .O(N__8498),
            .I(N__8494));
    InMux I__1840 (
            .O(N__8497),
            .I(N__8489));
    LocalMux I__1839 (
            .O(N__8494),
            .I(N__8485));
    InMux I__1838 (
            .O(N__8493),
            .I(N__8480));
    InMux I__1837 (
            .O(N__8492),
            .I(N__8480));
    LocalMux I__1836 (
            .O(N__8489),
            .I(N__8476));
    InMux I__1835 (
            .O(N__8488),
            .I(N__8473));
    Span4Mux_v I__1834 (
            .O(N__8485),
            .I(N__8470));
    LocalMux I__1833 (
            .O(N__8480),
            .I(N__8467));
    InMux I__1832 (
            .O(N__8479),
            .I(N__8464));
    Span4Mux_v I__1831 (
            .O(N__8476),
            .I(N__8450));
    LocalMux I__1830 (
            .O(N__8473),
            .I(N__8450));
    Span4Mux_h I__1829 (
            .O(N__8470),
            .I(N__8443));
    Span4Mux_v I__1828 (
            .O(N__8467),
            .I(N__8443));
    LocalMux I__1827 (
            .O(N__8464),
            .I(N__8443));
    InMux I__1826 (
            .O(N__8463),
            .I(N__8438));
    InMux I__1825 (
            .O(N__8462),
            .I(N__8438));
    InMux I__1824 (
            .O(N__8461),
            .I(N__8433));
    InMux I__1823 (
            .O(N__8460),
            .I(N__8433));
    InMux I__1822 (
            .O(N__8459),
            .I(N__8429));
    InMux I__1821 (
            .O(N__8458),
            .I(N__8420));
    InMux I__1820 (
            .O(N__8457),
            .I(N__8420));
    InMux I__1819 (
            .O(N__8456),
            .I(N__8420));
    InMux I__1818 (
            .O(N__8455),
            .I(N__8420));
    Span4Mux_v I__1817 (
            .O(N__8450),
            .I(N__8417));
    Sp12to4 I__1816 (
            .O(N__8443),
            .I(N__8412));
    LocalMux I__1815 (
            .O(N__8438),
            .I(N__8412));
    LocalMux I__1814 (
            .O(N__8433),
            .I(N__8409));
    InMux I__1813 (
            .O(N__8432),
            .I(N__8406));
    LocalMux I__1812 (
            .O(N__8429),
            .I(N__8401));
    LocalMux I__1811 (
            .O(N__8420),
            .I(N__8401));
    Sp12to4 I__1810 (
            .O(N__8417),
            .I(N__8392));
    Span12Mux_v I__1809 (
            .O(N__8412),
            .I(N__8392));
    Span12Mux_v I__1808 (
            .O(N__8409),
            .I(N__8392));
    LocalMux I__1807 (
            .O(N__8406),
            .I(N__8392));
    Span12Mux_h I__1806 (
            .O(N__8401),
            .I(N__8389));
    Span12Mux_h I__1805 (
            .O(N__8392),
            .I(N__8386));
    Odrv12 I__1804 (
            .O(N__8389),
            .I(RESETn_c));
    Odrv12 I__1803 (
            .O(N__8386),
            .I(RESETn_c));
    IoInMux I__1802 (
            .O(N__8381),
            .I(N__8378));
    LocalMux I__1801 (
            .O(N__8378),
            .I(N__8375));
    Span12Mux_s8_v I__1800 (
            .O(N__8375),
            .I(N__8371));
    InMux I__1799 (
            .O(N__8374),
            .I(N__8368));
    Odrv12 I__1798 (
            .O(N__8371),
            .I(RESETn_c_i));
    LocalMux I__1797 (
            .O(N__8368),
            .I(RESETn_c_i));
    CascadeMux I__1796 (
            .O(N__8363),
            .I(N__8359));
    CascadeMux I__1795 (
            .O(N__8362),
            .I(N__8355));
    InMux I__1794 (
            .O(N__8359),
            .I(N__8350));
    InMux I__1793 (
            .O(N__8358),
            .I(N__8350));
    InMux I__1792 (
            .O(N__8355),
            .I(N__8347));
    LocalMux I__1791 (
            .O(N__8350),
            .I(N__8344));
    LocalMux I__1790 (
            .O(N__8347),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    Odrv12 I__1789 (
            .O(N__8344),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    CascadeMux I__1788 (
            .O(N__8339),
            .I(N__8336));
    InMux I__1787 (
            .O(N__8336),
            .I(N__8332));
    IoInMux I__1786 (
            .O(N__8335),
            .I(N__8329));
    LocalMux I__1785 (
            .O(N__8332),
            .I(N__8325));
    LocalMux I__1784 (
            .O(N__8329),
            .I(N__8322));
    InMux I__1783 (
            .O(N__8328),
            .I(N__8319));
    Span4Mux_h I__1782 (
            .O(N__8325),
            .I(N__8316));
    Span12Mux_s3_h I__1781 (
            .O(N__8322),
            .I(N__8313));
    LocalMux I__1780 (
            .O(N__8319),
            .I(N__8310));
    Span4Mux_h I__1779 (
            .O(N__8316),
            .I(N__8307));
    Span12Mux_v I__1778 (
            .O(N__8313),
            .I(N__8304));
    Sp12to4 I__1777 (
            .O(N__8310),
            .I(N__8299));
    Sp12to4 I__1776 (
            .O(N__8307),
            .I(N__8299));
    Span12Mux_h I__1775 (
            .O(N__8304),
            .I(N__8296));
    Span12Mux_v I__1774 (
            .O(N__8299),
            .I(N__8293));
    Odrv12 I__1773 (
            .O(N__8296),
            .I(CLK40_PLL));
    Odrv12 I__1772 (
            .O(N__8293),
            .I(CLK40_PLL));
    InMux I__1771 (
            .O(N__8288),
            .I(N__8285));
    LocalMux I__1770 (
            .O(N__8285),
            .I(N__8281));
    InMux I__1769 (
            .O(N__8284),
            .I(N__8278));
    Span4Mux_v I__1768 (
            .O(N__8281),
            .I(N__8275));
    LocalMux I__1767 (
            .O(N__8278),
            .I(N__8272));
    Sp12to4 I__1766 (
            .O(N__8275),
            .I(N__8267));
    Span12Mux_v I__1765 (
            .O(N__8272),
            .I(N__8267));
    Odrv12 I__1764 (
            .O(N__8267),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ));
    InMux I__1763 (
            .O(N__8264),
            .I(N__8261));
    LocalMux I__1762 (
            .O(N__8261),
            .I(\U712_CYCLE_TERM.N_8 ));
    CascadeMux I__1761 (
            .O(N__8258),
            .I(N__8253));
    InMux I__1760 (
            .O(N__8257),
            .I(N__8250));
    InMux I__1759 (
            .O(N__8256),
            .I(N__8245));
    InMux I__1758 (
            .O(N__8253),
            .I(N__8242));
    LocalMux I__1757 (
            .O(N__8250),
            .I(N__8239));
    InMux I__1756 (
            .O(N__8249),
            .I(N__8236));
    InMux I__1755 (
            .O(N__8248),
            .I(N__8233));
    LocalMux I__1754 (
            .O(N__8245),
            .I(N__8228));
    LocalMux I__1753 (
            .O(N__8242),
            .I(N__8228));
    Span4Mux_h I__1752 (
            .O(N__8239),
            .I(N__8225));
    LocalMux I__1751 (
            .O(N__8236),
            .I(REG_TACK));
    LocalMux I__1750 (
            .O(N__8233),
            .I(REG_TACK));
    Odrv12 I__1749 (
            .O(N__8228),
            .I(REG_TACK));
    Odrv4 I__1748 (
            .O(N__8225),
            .I(REG_TACK));
    InMux I__1747 (
            .O(N__8216),
            .I(N__8213));
    LocalMux I__1746 (
            .O(N__8213),
            .I(N__8208));
    CascadeMux I__1745 (
            .O(N__8212),
            .I(N__8205));
    InMux I__1744 (
            .O(N__8211),
            .I(N__8201));
    Span4Mux_h I__1743 (
            .O(N__8208),
            .I(N__8198));
    InMux I__1742 (
            .O(N__8205),
            .I(N__8195));
    InMux I__1741 (
            .O(N__8204),
            .I(N__8191));
    LocalMux I__1740 (
            .O(N__8201),
            .I(N__8186));
    Span4Mux_h I__1739 (
            .O(N__8198),
            .I(N__8186));
    LocalMux I__1738 (
            .O(N__8195),
            .I(N__8183));
    InMux I__1737 (
            .O(N__8194),
            .I(N__8180));
    LocalMux I__1736 (
            .O(N__8191),
            .I(CPU_TACK));
    Odrv4 I__1735 (
            .O(N__8186),
            .I(CPU_TACK));
    Odrv12 I__1734 (
            .O(N__8183),
            .I(CPU_TACK));
    LocalMux I__1733 (
            .O(N__8180),
            .I(CPU_TACK));
    InMux I__1732 (
            .O(N__8171),
            .I(N__8164));
    InMux I__1731 (
            .O(N__8170),
            .I(N__8164));
    InMux I__1730 (
            .O(N__8169),
            .I(N__8161));
    LocalMux I__1729 (
            .O(N__8164),
            .I(N__8158));
    LocalMux I__1728 (
            .O(N__8161),
            .I(N__8155));
    Span4Mux_v I__1727 (
            .O(N__8158),
            .I(N__8148));
    Span4Mux_h I__1726 (
            .O(N__8155),
            .I(N__8148));
    InMux I__1725 (
            .O(N__8154),
            .I(N__8142));
    InMux I__1724 (
            .O(N__8153),
            .I(N__8142));
    Span4Mux_h I__1723 (
            .O(N__8148),
            .I(N__8139));
    InMux I__1722 (
            .O(N__8147),
            .I(N__8136));
    LocalMux I__1721 (
            .O(N__8142),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    Odrv4 I__1720 (
            .O(N__8139),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1719 (
            .O(N__8136),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    InMux I__1718 (
            .O(N__8129),
            .I(N__8126));
    LocalMux I__1717 (
            .O(N__8126),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1716 (
            .O(N__8123),
            .I(N__8119));
    InMux I__1715 (
            .O(N__8122),
            .I(N__8116));
    LocalMux I__1714 (
            .O(N__8119),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__1713 (
            .O(N__8116),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__1712 (
            .O(N__8111),
            .I(N__8108));
    LocalMux I__1711 (
            .O(N__8108),
            .I(N__8104));
    InMux I__1710 (
            .O(N__8107),
            .I(N__8101));
    Span4Mux_v I__1709 (
            .O(N__8104),
            .I(N__8098));
    LocalMux I__1708 (
            .O(N__8101),
            .I(N__8095));
    Span4Mux_h I__1707 (
            .O(N__8098),
            .I(N__8090));
    Span4Mux_v I__1706 (
            .O(N__8095),
            .I(N__8087));
    InMux I__1705 (
            .O(N__8094),
            .I(N__8084));
    InMux I__1704 (
            .O(N__8093),
            .I(N__8081));
    Sp12to4 I__1703 (
            .O(N__8090),
            .I(N__8078));
    Sp12to4 I__1702 (
            .O(N__8087),
            .I(N__8071));
    LocalMux I__1701 (
            .O(N__8084),
            .I(N__8071));
    LocalMux I__1700 (
            .O(N__8081),
            .I(N__8071));
    Span12Mux_h I__1699 (
            .O(N__8078),
            .I(N__8068));
    Span12Mux_v I__1698 (
            .O(N__8071),
            .I(N__8065));
    Span12Mux_v I__1697 (
            .O(N__8068),
            .I(N__8060));
    Span12Mux_h I__1696 (
            .O(N__8065),
            .I(N__8060));
    Odrv12 I__1695 (
            .O(N__8060),
            .I(CASLn_c));
    InMux I__1694 (
            .O(N__8057),
            .I(N__8053));
    InMux I__1693 (
            .O(N__8056),
            .I(N__8050));
    LocalMux I__1692 (
            .O(N__8053),
            .I(N__8046));
    LocalMux I__1691 (
            .O(N__8050),
            .I(N__8043));
    InMux I__1690 (
            .O(N__8049),
            .I(N__8040));
    Span4Mux_v I__1689 (
            .O(N__8046),
            .I(N__8034));
    Span4Mux_v I__1688 (
            .O(N__8043),
            .I(N__8034));
    LocalMux I__1687 (
            .O(N__8040),
            .I(N__8031));
    InMux I__1686 (
            .O(N__8039),
            .I(N__8028));
    Span4Mux_v I__1685 (
            .O(N__8034),
            .I(N__8021));
    Span4Mux_h I__1684 (
            .O(N__8031),
            .I(N__8021));
    LocalMux I__1683 (
            .O(N__8028),
            .I(N__8021));
    Span4Mux_v I__1682 (
            .O(N__8021),
            .I(N__8018));
    Span4Mux_v I__1681 (
            .O(N__8018),
            .I(N__8015));
    Sp12to4 I__1680 (
            .O(N__8015),
            .I(N__8012));
    Span12Mux_h I__1679 (
            .O(N__8012),
            .I(N__8009));
    Odrv12 I__1678 (
            .O(N__8009),
            .I(CASUn_c));
    InMux I__1677 (
            .O(N__8006),
            .I(N__8002));
    InMux I__1676 (
            .O(N__8005),
            .I(N__7999));
    LocalMux I__1675 (
            .O(N__8002),
            .I(N__7996));
    LocalMux I__1674 (
            .O(N__7999),
            .I(N__7993));
    Span4Mux_v I__1673 (
            .O(N__7996),
            .I(N__7989));
    Span4Mux_v I__1672 (
            .O(N__7993),
            .I(N__7986));
    InMux I__1671 (
            .O(N__7992),
            .I(N__7983));
    Odrv4 I__1670 (
            .O(N__7989),
            .I(REG_CYCLE));
    Odrv4 I__1669 (
            .O(N__7986),
            .I(REG_CYCLE));
    LocalMux I__1668 (
            .O(N__7983),
            .I(REG_CYCLE));
    IoInMux I__1667 (
            .O(N__7976),
            .I(N__7973));
    LocalMux I__1666 (
            .O(N__7973),
            .I(N__7970));
    IoSpan4Mux I__1665 (
            .O(N__7970),
            .I(N__7967));
    Span4Mux_s1_v I__1664 (
            .O(N__7967),
            .I(N__7964));
    Sp12to4 I__1663 (
            .O(N__7964),
            .I(N__7961));
    Span12Mux_h I__1662 (
            .O(N__7961),
            .I(N__7958));
    Odrv12 I__1661 (
            .O(N__7958),
            .I(DRDENn_c));
    CascadeMux I__1660 (
            .O(N__7955),
            .I(N__7949));
    CascadeMux I__1659 (
            .O(N__7954),
            .I(N__7943));
    InMux I__1658 (
            .O(N__7953),
            .I(N__7935));
    InMux I__1657 (
            .O(N__7952),
            .I(N__7932));
    InMux I__1656 (
            .O(N__7949),
            .I(N__7927));
    InMux I__1655 (
            .O(N__7948),
            .I(N__7927));
    InMux I__1654 (
            .O(N__7947),
            .I(N__7924));
    InMux I__1653 (
            .O(N__7946),
            .I(N__7919));
    InMux I__1652 (
            .O(N__7943),
            .I(N__7919));
    InMux I__1651 (
            .O(N__7942),
            .I(N__7916));
    InMux I__1650 (
            .O(N__7941),
            .I(N__7913));
    InMux I__1649 (
            .O(N__7940),
            .I(N__7908));
    InMux I__1648 (
            .O(N__7939),
            .I(N__7908));
    InMux I__1647 (
            .O(N__7938),
            .I(N__7905));
    LocalMux I__1646 (
            .O(N__7935),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1645 (
            .O(N__7932),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1644 (
            .O(N__7927),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1643 (
            .O(N__7924),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1642 (
            .O(N__7919),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1641 (
            .O(N__7916),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1640 (
            .O(N__7913),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1639 (
            .O(N__7908),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1638 (
            .O(N__7905),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    CascadeMux I__1637 (
            .O(N__7886),
            .I(N__7883));
    InMux I__1636 (
            .O(N__7883),
            .I(N__7878));
    InMux I__1635 (
            .O(N__7882),
            .I(N__7873));
    InMux I__1634 (
            .O(N__7881),
            .I(N__7870));
    LocalMux I__1633 (
            .O(N__7878),
            .I(N__7864));
    InMux I__1632 (
            .O(N__7877),
            .I(N__7861));
    InMux I__1631 (
            .O(N__7876),
            .I(N__7858));
    LocalMux I__1630 (
            .O(N__7873),
            .I(N__7847));
    LocalMux I__1629 (
            .O(N__7870),
            .I(N__7847));
    InMux I__1628 (
            .O(N__7869),
            .I(N__7840));
    InMux I__1627 (
            .O(N__7868),
            .I(N__7840));
    InMux I__1626 (
            .O(N__7867),
            .I(N__7840));
    Span4Mux_v I__1625 (
            .O(N__7864),
            .I(N__7832));
    LocalMux I__1624 (
            .O(N__7861),
            .I(N__7832));
    LocalMux I__1623 (
            .O(N__7858),
            .I(N__7832));
    InMux I__1622 (
            .O(N__7857),
            .I(N__7829));
    InMux I__1621 (
            .O(N__7856),
            .I(N__7823));
    InMux I__1620 (
            .O(N__7855),
            .I(N__7823));
    InMux I__1619 (
            .O(N__7854),
            .I(N__7816));
    InMux I__1618 (
            .O(N__7853),
            .I(N__7816));
    InMux I__1617 (
            .O(N__7852),
            .I(N__7816));
    Span4Mux_v I__1616 (
            .O(N__7847),
            .I(N__7811));
    LocalMux I__1615 (
            .O(N__7840),
            .I(N__7811));
    InMux I__1614 (
            .O(N__7839),
            .I(N__7808));
    Span4Mux_h I__1613 (
            .O(N__7832),
            .I(N__7803));
    LocalMux I__1612 (
            .O(N__7829),
            .I(N__7803));
    InMux I__1611 (
            .O(N__7828),
            .I(N__7800));
    LocalMux I__1610 (
            .O(N__7823),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1609 (
            .O(N__7816),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1608 (
            .O(N__7811),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1607 (
            .O(N__7808),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1606 (
            .O(N__7803),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1605 (
            .O(N__7800),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    CascadeMux I__1604 (
            .O(N__7787),
            .I(\U712_CHIP_RAM.N_396_cascade_ ));
    InMux I__1603 (
            .O(N__7784),
            .I(N__7781));
    LocalMux I__1602 (
            .O(N__7781),
            .I(N__7778));
    Span4Mux_v I__1601 (
            .O(N__7778),
            .I(N__7772));
    InMux I__1600 (
            .O(N__7777),
            .I(N__7767));
    InMux I__1599 (
            .O(N__7776),
            .I(N__7767));
    InMux I__1598 (
            .O(N__7775),
            .I(N__7764));
    Odrv4 I__1597 (
            .O(N__7772),
            .I(\U712_CHIP_RAM.N_436 ));
    LocalMux I__1596 (
            .O(N__7767),
            .I(\U712_CHIP_RAM.N_436 ));
    LocalMux I__1595 (
            .O(N__7764),
            .I(\U712_CHIP_RAM.N_436 ));
    CascadeMux I__1594 (
            .O(N__7757),
            .I(\U712_CHIP_RAM.N_436_cascade_ ));
    InMux I__1593 (
            .O(N__7754),
            .I(N__7751));
    LocalMux I__1592 (
            .O(N__7751),
            .I(N__7748));
    Span4Mux_h I__1591 (
            .O(N__7748),
            .I(N__7742));
    InMux I__1590 (
            .O(N__7747),
            .I(N__7737));
    InMux I__1589 (
            .O(N__7746),
            .I(N__7737));
    InMux I__1588 (
            .O(N__7745),
            .I(N__7734));
    Odrv4 I__1587 (
            .O(N__7742),
            .I(\U712_CHIP_RAM.N_257 ));
    LocalMux I__1586 (
            .O(N__7737),
            .I(\U712_CHIP_RAM.N_257 ));
    LocalMux I__1585 (
            .O(N__7734),
            .I(\U712_CHIP_RAM.N_257 ));
    InMux I__1584 (
            .O(N__7727),
            .I(N__7724));
    LocalMux I__1583 (
            .O(N__7724),
            .I(N__7721));
    Odrv4 I__1582 (
            .O(N__7721),
            .I(\U712_CHIP_RAM.N_357 ));
    InMux I__1581 (
            .O(N__7718),
            .I(N__7715));
    LocalMux I__1580 (
            .O(N__7715),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_1 ));
    CascadeMux I__1579 (
            .O(N__7712),
            .I(N__7708));
    InMux I__1578 (
            .O(N__7711),
            .I(N__7704));
    InMux I__1577 (
            .O(N__7708),
            .I(N__7700));
    CascadeMux I__1576 (
            .O(N__7707),
            .I(N__7697));
    LocalMux I__1575 (
            .O(N__7704),
            .I(N__7694));
    InMux I__1574 (
            .O(N__7703),
            .I(N__7691));
    LocalMux I__1573 (
            .O(N__7700),
            .I(N__7688));
    InMux I__1572 (
            .O(N__7697),
            .I(N__7685));
    Span4Mux_v I__1571 (
            .O(N__7694),
            .I(N__7677));
    LocalMux I__1570 (
            .O(N__7691),
            .I(N__7677));
    Span4Mux_v I__1569 (
            .O(N__7688),
            .I(N__7677));
    LocalMux I__1568 (
            .O(N__7685),
            .I(N__7674));
    InMux I__1567 (
            .O(N__7684),
            .I(N__7671));
    Odrv4 I__1566 (
            .O(N__7677),
            .I(\U712_CHIP_RAM.N_396 ));
    Odrv4 I__1565 (
            .O(N__7674),
            .I(\U712_CHIP_RAM.N_396 ));
    LocalMux I__1564 (
            .O(N__7671),
            .I(\U712_CHIP_RAM.N_396 ));
    InMux I__1563 (
            .O(N__7664),
            .I(N__7661));
    LocalMux I__1562 (
            .O(N__7661),
            .I(N__7655));
    InMux I__1561 (
            .O(N__7660),
            .I(N__7652));
    InMux I__1560 (
            .O(N__7659),
            .I(N__7648));
    CascadeMux I__1559 (
            .O(N__7658),
            .I(N__7645));
    Span4Mux_h I__1558 (
            .O(N__7655),
            .I(N__7638));
    LocalMux I__1557 (
            .O(N__7652),
            .I(N__7635));
    InMux I__1556 (
            .O(N__7651),
            .I(N__7632));
    LocalMux I__1555 (
            .O(N__7648),
            .I(N__7629));
    InMux I__1554 (
            .O(N__7645),
            .I(N__7626));
    InMux I__1553 (
            .O(N__7644),
            .I(N__7621));
    InMux I__1552 (
            .O(N__7643),
            .I(N__7621));
    InMux I__1551 (
            .O(N__7642),
            .I(N__7616));
    InMux I__1550 (
            .O(N__7641),
            .I(N__7616));
    Odrv4 I__1549 (
            .O(N__7638),
            .I(\U712_CHIP_RAM.N_384 ));
    Odrv4 I__1548 (
            .O(N__7635),
            .I(\U712_CHIP_RAM.N_384 ));
    LocalMux I__1547 (
            .O(N__7632),
            .I(\U712_CHIP_RAM.N_384 ));
    Odrv4 I__1546 (
            .O(N__7629),
            .I(\U712_CHIP_RAM.N_384 ));
    LocalMux I__1545 (
            .O(N__7626),
            .I(\U712_CHIP_RAM.N_384 ));
    LocalMux I__1544 (
            .O(N__7621),
            .I(\U712_CHIP_RAM.N_384 ));
    LocalMux I__1543 (
            .O(N__7616),
            .I(\U712_CHIP_RAM.N_384 ));
    InMux I__1542 (
            .O(N__7601),
            .I(N__7598));
    LocalMux I__1541 (
            .O(N__7598),
            .I(\U712_CHIP_RAM.N_351 ));
    CascadeMux I__1540 (
            .O(N__7595),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_cascade_ ));
    InMux I__1539 (
            .O(N__7592),
            .I(N__7589));
    LocalMux I__1538 (
            .O(N__7589),
            .I(\U712_CHIP_RAM.N_117 ));
    InMux I__1537 (
            .O(N__7586),
            .I(N__7582));
    InMux I__1536 (
            .O(N__7585),
            .I(N__7570));
    LocalMux I__1535 (
            .O(N__7582),
            .I(N__7567));
    InMux I__1534 (
            .O(N__7581),
            .I(N__7564));
    InMux I__1533 (
            .O(N__7580),
            .I(N__7561));
    InMux I__1532 (
            .O(N__7579),
            .I(N__7558));
    InMux I__1531 (
            .O(N__7578),
            .I(N__7555));
    InMux I__1530 (
            .O(N__7577),
            .I(N__7550));
    InMux I__1529 (
            .O(N__7576),
            .I(N__7550));
    InMux I__1528 (
            .O(N__7575),
            .I(N__7543));
    InMux I__1527 (
            .O(N__7574),
            .I(N__7543));
    InMux I__1526 (
            .O(N__7573),
            .I(N__7543));
    LocalMux I__1525 (
            .O(N__7570),
            .I(N__7540));
    Odrv12 I__1524 (
            .O(N__7567),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1523 (
            .O(N__7564),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1522 (
            .O(N__7561),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1521 (
            .O(N__7558),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1520 (
            .O(N__7555),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1519 (
            .O(N__7550),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1518 (
            .O(N__7543),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1517 (
            .O(N__7540),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    CascadeMux I__1516 (
            .O(N__7523),
            .I(N__7520));
    InMux I__1515 (
            .O(N__7520),
            .I(N__7516));
    InMux I__1514 (
            .O(N__7519),
            .I(N__7511));
    LocalMux I__1513 (
            .O(N__7516),
            .I(N__7508));
    InMux I__1512 (
            .O(N__7515),
            .I(N__7501));
    InMux I__1511 (
            .O(N__7514),
            .I(N__7498));
    LocalMux I__1510 (
            .O(N__7511),
            .I(N__7495));
    Span4Mux_v I__1509 (
            .O(N__7508),
            .I(N__7492));
    InMux I__1508 (
            .O(N__7507),
            .I(N__7487));
    InMux I__1507 (
            .O(N__7506),
            .I(N__7487));
    InMux I__1506 (
            .O(N__7505),
            .I(N__7484));
    InMux I__1505 (
            .O(N__7504),
            .I(N__7481));
    LocalMux I__1504 (
            .O(N__7501),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1503 (
            .O(N__7498),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1502 (
            .O(N__7495),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1501 (
            .O(N__7492),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1500 (
            .O(N__7487),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1499 (
            .O(N__7484),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1498 (
            .O(N__7481),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__1497 (
            .O(N__7466),
            .I(N__7457));
    InMux I__1496 (
            .O(N__7465),
            .I(N__7451));
    InMux I__1495 (
            .O(N__7464),
            .I(N__7446));
    InMux I__1494 (
            .O(N__7463),
            .I(N__7446));
    InMux I__1493 (
            .O(N__7462),
            .I(N__7442));
    InMux I__1492 (
            .O(N__7461),
            .I(N__7439));
    InMux I__1491 (
            .O(N__7460),
            .I(N__7436));
    InMux I__1490 (
            .O(N__7457),
            .I(N__7433));
    InMux I__1489 (
            .O(N__7456),
            .I(N__7428));
    InMux I__1488 (
            .O(N__7455),
            .I(N__7428));
    InMux I__1487 (
            .O(N__7454),
            .I(N__7425));
    LocalMux I__1486 (
            .O(N__7451),
            .I(N__7420));
    LocalMux I__1485 (
            .O(N__7446),
            .I(N__7420));
    InMux I__1484 (
            .O(N__7445),
            .I(N__7417));
    LocalMux I__1483 (
            .O(N__7442),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1482 (
            .O(N__7439),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1481 (
            .O(N__7436),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1480 (
            .O(N__7433),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1479 (
            .O(N__7428),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1478 (
            .O(N__7425),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1477 (
            .O(N__7420),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1476 (
            .O(N__7417),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    InMux I__1475 (
            .O(N__7400),
            .I(N__7397));
    LocalMux I__1474 (
            .O(N__7397),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_0_a2_0_2 ));
    CascadeMux I__1473 (
            .O(N__7394),
            .I(N__7390));
    InMux I__1472 (
            .O(N__7393),
            .I(N__7387));
    InMux I__1471 (
            .O(N__7390),
            .I(N__7384));
    LocalMux I__1470 (
            .O(N__7387),
            .I(N__7381));
    LocalMux I__1469 (
            .O(N__7384),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    Odrv12 I__1468 (
            .O(N__7381),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    CascadeMux I__1467 (
            .O(N__7376),
            .I(\U712_CYCLE_TERM.N_274_i_0_0_cascade_ ));
    CascadeMux I__1466 (
            .O(N__7373),
            .I(\U712_CYCLE_TERM.N_274_i_0_en_cascade_ ));
    CEMux I__1465 (
            .O(N__7370),
            .I(N__7367));
    LocalMux I__1464 (
            .O(N__7367),
            .I(N__7364));
    Span4Mux_h I__1463 (
            .O(N__7364),
            .I(N__7361));
    Span4Mux_h I__1462 (
            .O(N__7361),
            .I(N__7358));
    Odrv4 I__1461 (
            .O(N__7358),
            .I(\U712_CYCLE_TERM.N_274_i_0_en_0 ));
    InMux I__1460 (
            .O(N__7355),
            .I(N__7352));
    LocalMux I__1459 (
            .O(N__7352),
            .I(N__7349));
    Span4Mux_h I__1458 (
            .O(N__7349),
            .I(N__7346));
    Odrv4 I__1457 (
            .O(N__7346),
            .I(\U712_CHIP_RAM.N_294 ));
    InMux I__1456 (
            .O(N__7343),
            .I(N__7338));
    CascadeMux I__1455 (
            .O(N__7342),
            .I(N__7335));
    CascadeMux I__1454 (
            .O(N__7341),
            .I(N__7332));
    LocalMux I__1453 (
            .O(N__7338),
            .I(N__7327));
    InMux I__1452 (
            .O(N__7335),
            .I(N__7324));
    InMux I__1451 (
            .O(N__7332),
            .I(N__7320));
    InMux I__1450 (
            .O(N__7331),
            .I(N__7317));
    InMux I__1449 (
            .O(N__7330),
            .I(N__7314));
    Span4Mux_v I__1448 (
            .O(N__7327),
            .I(N__7309));
    LocalMux I__1447 (
            .O(N__7324),
            .I(N__7309));
    InMux I__1446 (
            .O(N__7323),
            .I(N__7306));
    LocalMux I__1445 (
            .O(N__7320),
            .I(N__7301));
    LocalMux I__1444 (
            .O(N__7317),
            .I(N__7301));
    LocalMux I__1443 (
            .O(N__7314),
            .I(N__7298));
    Span4Mux_h I__1442 (
            .O(N__7309),
            .I(N__7295));
    LocalMux I__1441 (
            .O(N__7306),
            .I(N__7292));
    Span4Mux_h I__1440 (
            .O(N__7301),
            .I(N__7289));
    Odrv4 I__1439 (
            .O(N__7298),
            .I(DMA_CYCLE));
    Odrv4 I__1438 (
            .O(N__7295),
            .I(DMA_CYCLE));
    Odrv12 I__1437 (
            .O(N__7292),
            .I(DMA_CYCLE));
    Odrv4 I__1436 (
            .O(N__7289),
            .I(DMA_CYCLE));
    CascadeMux I__1435 (
            .O(N__7280),
            .I(\U712_CHIP_RAM.N_305_cascade_ ));
    InMux I__1434 (
            .O(N__7277),
            .I(N__7274));
    LocalMux I__1433 (
            .O(N__7274),
            .I(N__7267));
    InMux I__1432 (
            .O(N__7273),
            .I(N__7262));
    InMux I__1431 (
            .O(N__7272),
            .I(N__7262));
    InMux I__1430 (
            .O(N__7271),
            .I(N__7259));
    InMux I__1429 (
            .O(N__7270),
            .I(N__7256));
    Odrv4 I__1428 (
            .O(N__7267),
            .I(\U712_CHIP_RAM.N_388 ));
    LocalMux I__1427 (
            .O(N__7262),
            .I(\U712_CHIP_RAM.N_388 ));
    LocalMux I__1426 (
            .O(N__7259),
            .I(\U712_CHIP_RAM.N_388 ));
    LocalMux I__1425 (
            .O(N__7256),
            .I(\U712_CHIP_RAM.N_388 ));
    CascadeMux I__1424 (
            .O(N__7247),
            .I(N__7242));
    CascadeMux I__1423 (
            .O(N__7246),
            .I(N__7238));
    InMux I__1422 (
            .O(N__7245),
            .I(N__7233));
    InMux I__1421 (
            .O(N__7242),
            .I(N__7229));
    InMux I__1420 (
            .O(N__7241),
            .I(N__7226));
    InMux I__1419 (
            .O(N__7238),
            .I(N__7223));
    CascadeMux I__1418 (
            .O(N__7237),
            .I(N__7219));
    CascadeMux I__1417 (
            .O(N__7236),
            .I(N__7216));
    LocalMux I__1416 (
            .O(N__7233),
            .I(N__7210));
    InMux I__1415 (
            .O(N__7232),
            .I(N__7207));
    LocalMux I__1414 (
            .O(N__7229),
            .I(N__7202));
    LocalMux I__1413 (
            .O(N__7226),
            .I(N__7202));
    LocalMux I__1412 (
            .O(N__7223),
            .I(N__7199));
    InMux I__1411 (
            .O(N__7222),
            .I(N__7196));
    InMux I__1410 (
            .O(N__7219),
            .I(N__7191));
    InMux I__1409 (
            .O(N__7216),
            .I(N__7191));
    InMux I__1408 (
            .O(N__7215),
            .I(N__7188));
    InMux I__1407 (
            .O(N__7214),
            .I(N__7185));
    InMux I__1406 (
            .O(N__7213),
            .I(N__7182));
    Span4Mux_h I__1405 (
            .O(N__7210),
            .I(N__7179));
    LocalMux I__1404 (
            .O(N__7207),
            .I(\U712_CHIP_RAM.N_45_i ));
    Odrv4 I__1403 (
            .O(N__7202),
            .I(\U712_CHIP_RAM.N_45_i ));
    Odrv4 I__1402 (
            .O(N__7199),
            .I(\U712_CHIP_RAM.N_45_i ));
    LocalMux I__1401 (
            .O(N__7196),
            .I(\U712_CHIP_RAM.N_45_i ));
    LocalMux I__1400 (
            .O(N__7191),
            .I(\U712_CHIP_RAM.N_45_i ));
    LocalMux I__1399 (
            .O(N__7188),
            .I(\U712_CHIP_RAM.N_45_i ));
    LocalMux I__1398 (
            .O(N__7185),
            .I(\U712_CHIP_RAM.N_45_i ));
    LocalMux I__1397 (
            .O(N__7182),
            .I(\U712_CHIP_RAM.N_45_i ));
    Odrv4 I__1396 (
            .O(N__7179),
            .I(\U712_CHIP_RAM.N_45_i ));
    CascadeMux I__1395 (
            .O(N__7160),
            .I(\U712_CHIP_RAM.N_346_cascade_ ));
    InMux I__1394 (
            .O(N__7157),
            .I(N__7154));
    LocalMux I__1393 (
            .O(N__7154),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_2 ));
    CascadeMux I__1392 (
            .O(N__7151),
            .I(N__7147));
    InMux I__1391 (
            .O(N__7150),
            .I(N__7144));
    InMux I__1390 (
            .O(N__7147),
            .I(N__7140));
    LocalMux I__1389 (
            .O(N__7144),
            .I(N__7137));
    InMux I__1388 (
            .O(N__7143),
            .I(N__7134));
    LocalMux I__1387 (
            .O(N__7140),
            .I(\U712_CHIP_RAM.N_407 ));
    Odrv4 I__1386 (
            .O(N__7137),
            .I(\U712_CHIP_RAM.N_407 ));
    LocalMux I__1385 (
            .O(N__7134),
            .I(\U712_CHIP_RAM.N_407 ));
    CascadeMux I__1384 (
            .O(N__7127),
            .I(\U712_CHIP_RAM.N_407_cascade_ ));
    InMux I__1383 (
            .O(N__7124),
            .I(N__7120));
    InMux I__1382 (
            .O(N__7123),
            .I(N__7114));
    LocalMux I__1381 (
            .O(N__7120),
            .I(N__7111));
    InMux I__1380 (
            .O(N__7119),
            .I(N__7108));
    InMux I__1379 (
            .O(N__7118),
            .I(N__7103));
    InMux I__1378 (
            .O(N__7117),
            .I(N__7103));
    LocalMux I__1377 (
            .O(N__7114),
            .I(\U712_CHIP_RAM.N_400 ));
    Odrv4 I__1376 (
            .O(N__7111),
            .I(\U712_CHIP_RAM.N_400 ));
    LocalMux I__1375 (
            .O(N__7108),
            .I(\U712_CHIP_RAM.N_400 ));
    LocalMux I__1374 (
            .O(N__7103),
            .I(\U712_CHIP_RAM.N_400 ));
    InMux I__1373 (
            .O(N__7094),
            .I(N__7090));
    CascadeMux I__1372 (
            .O(N__7093),
            .I(N__7087));
    LocalMux I__1371 (
            .O(N__7090),
            .I(N__7084));
    InMux I__1370 (
            .O(N__7087),
            .I(N__7081));
    Span4Mux_v I__1369 (
            .O(N__7084),
            .I(N__7075));
    LocalMux I__1368 (
            .O(N__7081),
            .I(N__7072));
    InMux I__1367 (
            .O(N__7080),
            .I(N__7067));
    InMux I__1366 (
            .O(N__7079),
            .I(N__7067));
    CascadeMux I__1365 (
            .O(N__7078),
            .I(N__7063));
    Span4Mux_v I__1364 (
            .O(N__7075),
            .I(N__7057));
    Span4Mux_h I__1363 (
            .O(N__7072),
            .I(N__7057));
    LocalMux I__1362 (
            .O(N__7067),
            .I(N__7054));
    InMux I__1361 (
            .O(N__7066),
            .I(N__7049));
    InMux I__1360 (
            .O(N__7063),
            .I(N__7049));
    InMux I__1359 (
            .O(N__7062),
            .I(N__7046));
    Odrv4 I__1358 (
            .O(N__7057),
            .I(WRITE_CYCLE));
    Odrv4 I__1357 (
            .O(N__7054),
            .I(WRITE_CYCLE));
    LocalMux I__1356 (
            .O(N__7049),
            .I(WRITE_CYCLE));
    LocalMux I__1355 (
            .O(N__7046),
            .I(WRITE_CYCLE));
    CascadeMux I__1354 (
            .O(N__7037),
            .I(\U712_CHIP_RAM.N_257_cascade_ ));
    CascadeMux I__1353 (
            .O(N__7034),
            .I(\U712_BYTE_ENABLE.UUBE_cascade_ ));
    IoInMux I__1352 (
            .O(N__7031),
            .I(N__7028));
    LocalMux I__1351 (
            .O(N__7028),
            .I(N__7025));
    Span4Mux_s3_h I__1350 (
            .O(N__7025),
            .I(N__7022));
    Span4Mux_v I__1349 (
            .O(N__7022),
            .I(N__7019));
    Span4Mux_h I__1348 (
            .O(N__7019),
            .I(N__7016));
    Span4Mux_h I__1347 (
            .O(N__7016),
            .I(N__7013));
    Span4Mux_h I__1346 (
            .O(N__7013),
            .I(N__7010));
    Odrv4 I__1345 (
            .O(N__7010),
            .I(N_48_i));
    CascadeMux I__1344 (
            .O(N__7007),
            .I(N__7004));
    InMux I__1343 (
            .O(N__7004),
            .I(N__7001));
    LocalMux I__1342 (
            .O(N__7001),
            .I(N__6998));
    Odrv12 I__1341 (
            .O(N__6998),
            .I(\U712_BYTE_ENABLE.N_278 ));
    InMux I__1340 (
            .O(N__6995),
            .I(N__6992));
    LocalMux I__1339 (
            .O(N__6992),
            .I(N__6989));
    Odrv4 I__1338 (
            .O(N__6989),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0 ));
    IoInMux I__1337 (
            .O(N__6986),
            .I(N__6983));
    LocalMux I__1336 (
            .O(N__6983),
            .I(N__6980));
    Span12Mux_s4_h I__1335 (
            .O(N__6980),
            .I(N__6977));
    Span12Mux_h I__1334 (
            .O(N__6977),
            .I(N__6974));
    Span12Mux_v I__1333 (
            .O(N__6974),
            .I(N__6971));
    Odrv12 I__1332 (
            .O(N__6971),
            .I(N_49_i));
    CascadeMux I__1331 (
            .O(N__6968),
            .I(N__6965));
    InMux I__1330 (
            .O(N__6965),
            .I(N__6962));
    LocalMux I__1329 (
            .O(N__6962),
            .I(\U712_BYTE_ENABLE.N_277 ));
    IoInMux I__1328 (
            .O(N__6959),
            .I(N__6956));
    LocalMux I__1327 (
            .O(N__6956),
            .I(N__6953));
    Span4Mux_s2_v I__1326 (
            .O(N__6953),
            .I(N__6950));
    Sp12to4 I__1325 (
            .O(N__6950),
            .I(N__6946));
    InMux I__1324 (
            .O(N__6949),
            .I(N__6943));
    Span12Mux_h I__1323 (
            .O(N__6946),
            .I(N__6938));
    LocalMux I__1322 (
            .O(N__6943),
            .I(N__6935));
    InMux I__1321 (
            .O(N__6942),
            .I(N__6932));
    InMux I__1320 (
            .O(N__6941),
            .I(N__6929));
    Odrv12 I__1319 (
            .O(N__6938),
            .I(DBENn_c));
    Odrv4 I__1318 (
            .O(N__6935),
            .I(DBENn_c));
    LocalMux I__1317 (
            .O(N__6932),
            .I(DBENn_c));
    LocalMux I__1316 (
            .O(N__6929),
            .I(DBENn_c));
    InMux I__1315 (
            .O(N__6920),
            .I(N__6914));
    InMux I__1314 (
            .O(N__6919),
            .I(N__6914));
    LocalMux I__1313 (
            .O(N__6914),
            .I(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0Z0Z_0 ));
    InMux I__1312 (
            .O(N__6911),
            .I(N__6908));
    LocalMux I__1311 (
            .O(N__6908),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_2_0 ));
    CascadeMux I__1310 (
            .O(N__6905),
            .I(\U712_CHIP_RAM.N_325_0_cascade_ ));
    InMux I__1309 (
            .O(N__6902),
            .I(N__6899));
    LocalMux I__1308 (
            .O(N__6899),
            .I(N__6896));
    Odrv4 I__1307 (
            .O(N__6896),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ));
    CascadeMux I__1306 (
            .O(N__6893),
            .I(N__6890));
    InMux I__1305 (
            .O(N__6890),
            .I(N__6887));
    LocalMux I__1304 (
            .O(N__6887),
            .I(N__6884));
    Span4Mux_h I__1303 (
            .O(N__6884),
            .I(N__6881));
    Odrv4 I__1302 (
            .O(N__6881),
            .I(\U712_CHIP_RAM.N_365_1 ));
    IoInMux I__1301 (
            .O(N__6878),
            .I(N__6875));
    LocalMux I__1300 (
            .O(N__6875),
            .I(N__6872));
    Span4Mux_s2_v I__1299 (
            .O(N__6872),
            .I(N__6869));
    Span4Mux_v I__1298 (
            .O(N__6869),
            .I(N__6866));
    Odrv4 I__1297 (
            .O(N__6866),
            .I(CONSTANT_ONE_NET));
    InMux I__1296 (
            .O(N__6863),
            .I(N__6860));
    LocalMux I__1295 (
            .O(N__6860),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__1294 (
            .O(N__6857),
            .I(N__6854));
    LocalMux I__1293 (
            .O(N__6854),
            .I(N__6851));
    Span4Mux_s3_h I__1292 (
            .O(N__6851),
            .I(N__6848));
    Span4Mux_v I__1291 (
            .O(N__6848),
            .I(N__6845));
    Sp12to4 I__1290 (
            .O(N__6845),
            .I(N__6842));
    Span12Mux_h I__1289 (
            .O(N__6842),
            .I(N__6839));
    Odrv12 I__1288 (
            .O(N__6839),
            .I(CMA_c_7));
    InMux I__1287 (
            .O(N__6836),
            .I(N__6833));
    LocalMux I__1286 (
            .O(N__6833),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__1285 (
            .O(N__6830),
            .I(N__6827));
    LocalMux I__1284 (
            .O(N__6827),
            .I(N__6824));
    IoSpan4Mux I__1283 (
            .O(N__6824),
            .I(N__6821));
    Sp12to4 I__1282 (
            .O(N__6821),
            .I(N__6818));
    Span12Mux_s9_h I__1281 (
            .O(N__6818),
            .I(N__6815));
    Span12Mux_v I__1280 (
            .O(N__6815),
            .I(N__6812));
    Odrv12 I__1279 (
            .O(N__6812),
            .I(CMA_c_4));
    InMux I__1278 (
            .O(N__6809),
            .I(N__6806));
    LocalMux I__1277 (
            .O(N__6806),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__1276 (
            .O(N__6803),
            .I(N__6800));
    LocalMux I__1275 (
            .O(N__6800),
            .I(N__6797));
    IoSpan4Mux I__1274 (
            .O(N__6797),
            .I(N__6794));
    Span4Mux_s2_h I__1273 (
            .O(N__6794),
            .I(N__6791));
    Sp12to4 I__1272 (
            .O(N__6791),
            .I(N__6788));
    Span12Mux_h I__1271 (
            .O(N__6788),
            .I(N__6785));
    Odrv12 I__1270 (
            .O(N__6785),
            .I(CMA_c_3));
    InMux I__1269 (
            .O(N__6782),
            .I(N__6779));
    LocalMux I__1268 (
            .O(N__6779),
            .I(N__6776));
    Odrv4 I__1267 (
            .O(N__6776),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__1266 (
            .O(N__6773),
            .I(N__6770));
    LocalMux I__1265 (
            .O(N__6770),
            .I(N__6767));
    IoSpan4Mux I__1264 (
            .O(N__6767),
            .I(N__6764));
    Span4Mux_s3_h I__1263 (
            .O(N__6764),
            .I(N__6761));
    Span4Mux_v I__1262 (
            .O(N__6761),
            .I(N__6758));
    Span4Mux_v I__1261 (
            .O(N__6758),
            .I(N__6755));
    Sp12to4 I__1260 (
            .O(N__6755),
            .I(N__6752));
    Odrv12 I__1259 (
            .O(N__6752),
            .I(CMA_c_6));
    InMux I__1258 (
            .O(N__6749),
            .I(N__6746));
    LocalMux I__1257 (
            .O(N__6746),
            .I(N__6743));
    Span12Mux_v I__1256 (
            .O(N__6743),
            .I(N__6740));
    Span12Mux_h I__1255 (
            .O(N__6740),
            .I(N__6737));
    Odrv12 I__1254 (
            .O(N__6737),
            .I(A_c_19));
    IoInMux I__1253 (
            .O(N__6734),
            .I(N__6731));
    LocalMux I__1252 (
            .O(N__6731),
            .I(N__6728));
    Span12Mux_s4_h I__1251 (
            .O(N__6728),
            .I(N__6725));
    Span12Mux_h I__1250 (
            .O(N__6725),
            .I(N__6722));
    Odrv12 I__1249 (
            .O(N__6722),
            .I(CMA_c_9));
    InMux I__1248 (
            .O(N__6719),
            .I(N__6716));
    LocalMux I__1247 (
            .O(N__6716),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    IoInMux I__1246 (
            .O(N__6713),
            .I(N__6710));
    LocalMux I__1245 (
            .O(N__6710),
            .I(N__6707));
    Span4Mux_s1_v I__1244 (
            .O(N__6707),
            .I(N__6704));
    Span4Mux_v I__1243 (
            .O(N__6704),
            .I(N__6701));
    Span4Mux_v I__1242 (
            .O(N__6701),
            .I(N__6698));
    Span4Mux_v I__1241 (
            .O(N__6698),
            .I(N__6695));
    Odrv4 I__1240 (
            .O(N__6695),
            .I(CMA_c_2));
    IoInMux I__1239 (
            .O(N__6692),
            .I(N__6689));
    LocalMux I__1238 (
            .O(N__6689),
            .I(N__6686));
    Span4Mux_s0_h I__1237 (
            .O(N__6686),
            .I(N__6683));
    Span4Mux_h I__1236 (
            .O(N__6683),
            .I(N__6680));
    Sp12to4 I__1235 (
            .O(N__6680),
            .I(N__6677));
    Span12Mux_s10_v I__1234 (
            .O(N__6677),
            .I(N__6674));
    Span12Mux_h I__1233 (
            .O(N__6674),
            .I(N__6671));
    Odrv12 I__1232 (
            .O(N__6671),
            .I(N_46_i));
    InMux I__1231 (
            .O(N__6668),
            .I(N__6665));
    LocalMux I__1230 (
            .O(N__6665),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0_0 ));
    CascadeMux I__1229 (
            .O(N__6662),
            .I(N__6657));
    CascadeMux I__1228 (
            .O(N__6661),
            .I(N__6650));
    InMux I__1227 (
            .O(N__6660),
            .I(N__6645));
    InMux I__1226 (
            .O(N__6657),
            .I(N__6642));
    InMux I__1225 (
            .O(N__6656),
            .I(N__6635));
    InMux I__1224 (
            .O(N__6655),
            .I(N__6635));
    InMux I__1223 (
            .O(N__6654),
            .I(N__6635));
    InMux I__1222 (
            .O(N__6653),
            .I(N__6632));
    InMux I__1221 (
            .O(N__6650),
            .I(N__6627));
    InMux I__1220 (
            .O(N__6649),
            .I(N__6627));
    InMux I__1219 (
            .O(N__6648),
            .I(N__6624));
    LocalMux I__1218 (
            .O(N__6645),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1217 (
            .O(N__6642),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1216 (
            .O(N__6635),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1215 (
            .O(N__6632),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1214 (
            .O(N__6627),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1213 (
            .O(N__6624),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CascadeMux I__1212 (
            .O(N__6611),
            .I(N__6608));
    InMux I__1211 (
            .O(N__6608),
            .I(N__6605));
    LocalMux I__1210 (
            .O(N__6605),
            .I(N__6602));
    Odrv4 I__1209 (
            .O(N__6602),
            .I(\U712_CHIP_RAM.N_444 ));
    CascadeMux I__1208 (
            .O(N__6599),
            .I(N__6596));
    InMux I__1207 (
            .O(N__6596),
            .I(N__6592));
    InMux I__1206 (
            .O(N__6595),
            .I(N__6589));
    LocalMux I__1205 (
            .O(N__6592),
            .I(N__6586));
    LocalMux I__1204 (
            .O(N__6589),
            .I(N__6583));
    Span4Mux_h I__1203 (
            .O(N__6586),
            .I(N__6579));
    Span4Mux_h I__1202 (
            .O(N__6583),
            .I(N__6576));
    InMux I__1201 (
            .O(N__6582),
            .I(N__6573));
    Odrv4 I__1200 (
            .O(N__6579),
            .I(\U712_CHIP_RAM.N_392 ));
    Odrv4 I__1199 (
            .O(N__6576),
            .I(\U712_CHIP_RAM.N_392 ));
    LocalMux I__1198 (
            .O(N__6573),
            .I(\U712_CHIP_RAM.N_392 ));
    CascadeMux I__1197 (
            .O(N__6566),
            .I(\U712_CHIP_RAM.N_444_cascade_ ));
    InMux I__1196 (
            .O(N__6563),
            .I(N__6560));
    LocalMux I__1195 (
            .O(N__6560),
            .I(N__6556));
    InMux I__1194 (
            .O(N__6559),
            .I(N__6553));
    Odrv12 I__1193 (
            .O(N__6556),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0 ));
    LocalMux I__1192 (
            .O(N__6553),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0 ));
    InMux I__1191 (
            .O(N__6548),
            .I(N__6545));
    LocalMux I__1190 (
            .O(N__6545),
            .I(N__6542));
    Odrv4 I__1189 (
            .O(N__6542),
            .I(\U712_CHIP_RAM.N_334 ));
    CascadeMux I__1188 (
            .O(N__6539),
            .I(\U712_CHIP_RAM.N_334_cascade_ ));
    InMux I__1187 (
            .O(N__6536),
            .I(N__6533));
    LocalMux I__1186 (
            .O(N__6533),
            .I(N__6530));
    Odrv12 I__1185 (
            .O(N__6530),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0 ));
    CascadeMux I__1184 (
            .O(N__6527),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_ ));
    CEMux I__1183 (
            .O(N__6524),
            .I(N__6521));
    LocalMux I__1182 (
            .O(N__6521),
            .I(N__6518));
    Span4Mux_h I__1181 (
            .O(N__6518),
            .I(N__6515));
    Odrv4 I__1180 (
            .O(N__6515),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0 ));
    CascadeMux I__1179 (
            .O(N__6512),
            .I(N__6508));
    CascadeMux I__1178 (
            .O(N__6511),
            .I(N__6505));
    InMux I__1177 (
            .O(N__6508),
            .I(N__6502));
    InMux I__1176 (
            .O(N__6505),
            .I(N__6499));
    LocalMux I__1175 (
            .O(N__6502),
            .I(\U712_CHIP_RAM.N_448 ));
    LocalMux I__1174 (
            .O(N__6499),
            .I(\U712_CHIP_RAM.N_448 ));
    InMux I__1173 (
            .O(N__6494),
            .I(N__6491));
    LocalMux I__1172 (
            .O(N__6491),
            .I(\U712_CHIP_RAM.N_323 ));
    CascadeMux I__1171 (
            .O(N__6488),
            .I(\U712_CHIP_RAM.N_323_cascade_ ));
    InMux I__1170 (
            .O(N__6485),
            .I(N__6482));
    LocalMux I__1169 (
            .O(N__6482),
            .I(N__6479));
    Odrv4 I__1168 (
            .O(N__6479),
            .I(\U712_CHIP_RAM.un3_DMA_CYCLE_START ));
    InMux I__1167 (
            .O(N__6476),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    InMux I__1166 (
            .O(N__6473),
            .I(N__6470));
    LocalMux I__1165 (
            .O(N__6470),
            .I(N__6467));
    Odrv4 I__1164 (
            .O(N__6467),
            .I(\U712_CHIP_RAM.N_363 ));
    InMux I__1163 (
            .O(N__6464),
            .I(N__6460));
    InMux I__1162 (
            .O(N__6463),
            .I(N__6457));
    LocalMux I__1161 (
            .O(N__6460),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1160 (
            .O(N__6457),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    InMux I__1159 (
            .O(N__6452),
            .I(N__6448));
    InMux I__1158 (
            .O(N__6451),
            .I(N__6445));
    LocalMux I__1157 (
            .O(N__6448),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__1156 (
            .O(N__6445),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__1155 (
            .O(N__6440),
            .I(N__6436));
    InMux I__1154 (
            .O(N__6439),
            .I(N__6433));
    LocalMux I__1153 (
            .O(N__6436),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__1152 (
            .O(N__6433),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__1151 (
            .O(N__6428),
            .I(\U712_CHIP_RAM.N_384_cascade_ ));
    CascadeMux I__1150 (
            .O(N__6425),
            .I(\U712_CHIP_RAM.N_448_cascade_ ));
    InMux I__1149 (
            .O(N__6422),
            .I(N__6419));
    LocalMux I__1148 (
            .O(N__6419),
            .I(\U712_CHIP_RAM.N_255 ));
    CascadeMux I__1147 (
            .O(N__6416),
            .I(\U712_CHIP_RAM.N_255_cascade_ ));
    InMux I__1146 (
            .O(N__6413),
            .I(N__6410));
    LocalMux I__1145 (
            .O(N__6410),
            .I(\U712_CHIP_RAM.N_269 ));
    CascadeMux I__1144 (
            .O(N__6407),
            .I(N__6404));
    InMux I__1143 (
            .O(N__6404),
            .I(N__6401));
    LocalMux I__1142 (
            .O(N__6401),
            .I(N__6394));
    InMux I__1141 (
            .O(N__6400),
            .I(N__6391));
    InMux I__1140 (
            .O(N__6399),
            .I(N__6386));
    InMux I__1139 (
            .O(N__6398),
            .I(N__6386));
    InMux I__1138 (
            .O(N__6397),
            .I(N__6383));
    Odrv4 I__1137 (
            .O(N__6394),
            .I(\U712_CHIP_RAM.N_324 ));
    LocalMux I__1136 (
            .O(N__6391),
            .I(\U712_CHIP_RAM.N_324 ));
    LocalMux I__1135 (
            .O(N__6386),
            .I(\U712_CHIP_RAM.N_324 ));
    LocalMux I__1134 (
            .O(N__6383),
            .I(\U712_CHIP_RAM.N_324 ));
    CascadeMux I__1133 (
            .O(N__6374),
            .I(\U712_CHIP_RAM.N_456_cascade_ ));
    InMux I__1132 (
            .O(N__6371),
            .I(N__6365));
    InMux I__1131 (
            .O(N__6370),
            .I(N__6362));
    InMux I__1130 (
            .O(N__6369),
            .I(N__6357));
    InMux I__1129 (
            .O(N__6368),
            .I(N__6357));
    LocalMux I__1128 (
            .O(N__6365),
            .I(N__6352));
    LocalMux I__1127 (
            .O(N__6362),
            .I(N__6352));
    LocalMux I__1126 (
            .O(N__6357),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1 ));
    Odrv4 I__1125 (
            .O(N__6352),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1 ));
    InMux I__1124 (
            .O(N__6347),
            .I(bfn_11_11_0_));
    InMux I__1123 (
            .O(N__6344),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    InMux I__1122 (
            .O(N__6341),
            .I(N__6338));
    LocalMux I__1121 (
            .O(N__6338),
            .I(N__6334));
    InMux I__1120 (
            .O(N__6337),
            .I(N__6331));
    Odrv4 I__1119 (
            .O(N__6334),
            .I(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa ));
    LocalMux I__1118 (
            .O(N__6331),
            .I(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa ));
    InMux I__1117 (
            .O(N__6326),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    InMux I__1116 (
            .O(N__6323),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__1115 (
            .O(N__6320),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__1114 (
            .O(N__6317),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__1113 (
            .O(N__6314),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    CascadeMux I__1112 (
            .O(N__6311),
            .I(N__6308));
    InMux I__1111 (
            .O(N__6308),
            .I(N__6305));
    LocalMux I__1110 (
            .O(N__6305),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ));
    CascadeMux I__1109 (
            .O(N__6302),
            .I(\U712_CHIP_RAM.CMA_5_0_8_cascade_ ));
    InMux I__1108 (
            .O(N__6299),
            .I(N__6296));
    LocalMux I__1107 (
            .O(N__6296),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    InMux I__1106 (
            .O(N__6293),
            .I(N__6290));
    LocalMux I__1105 (
            .O(N__6290),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ));
    InMux I__1104 (
            .O(N__6287),
            .I(N__6281));
    InMux I__1103 (
            .O(N__6286),
            .I(N__6281));
    LocalMux I__1102 (
            .O(N__6281),
            .I(N__6278));
    Span4Mux_v I__1101 (
            .O(N__6278),
            .I(N__6275));
    Sp12to4 I__1100 (
            .O(N__6275),
            .I(N__6272));
    Span12Mux_h I__1099 (
            .O(N__6272),
            .I(N__6269));
    Odrv12 I__1098 (
            .O(N__6269),
            .I(A_c_10));
    InMux I__1097 (
            .O(N__6266),
            .I(N__6263));
    LocalMux I__1096 (
            .O(N__6263),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    InMux I__1095 (
            .O(N__6260),
            .I(N__6257));
    LocalMux I__1094 (
            .O(N__6257),
            .I(N__6253));
    InMux I__1093 (
            .O(N__6256),
            .I(N__6250));
    Span4Mux_v I__1092 (
            .O(N__6253),
            .I(N__6245));
    LocalMux I__1091 (
            .O(N__6250),
            .I(N__6245));
    Span4Mux_v I__1090 (
            .O(N__6245),
            .I(N__6242));
    Sp12to4 I__1089 (
            .O(N__6242),
            .I(N__6239));
    Span12Mux_h I__1088 (
            .O(N__6239),
            .I(N__6236));
    Odrv12 I__1087 (
            .O(N__6236),
            .I(AWEn_c));
    IoInMux I__1086 (
            .O(N__6233),
            .I(N__6230));
    LocalMux I__1085 (
            .O(N__6230),
            .I(N__6227));
    Span4Mux_s2_v I__1084 (
            .O(N__6227),
            .I(N__6224));
    Span4Mux_h I__1083 (
            .O(N__6224),
            .I(N__6220));
    CascadeMux I__1082 (
            .O(N__6223),
            .I(N__6217));
    Sp12to4 I__1081 (
            .O(N__6220),
            .I(N__6214));
    InMux I__1080 (
            .O(N__6217),
            .I(N__6211));
    Odrv12 I__1079 (
            .O(N__6214),
            .I(DBDIR_c));
    LocalMux I__1078 (
            .O(N__6211),
            .I(DBDIR_c));
    InMux I__1077 (
            .O(N__6206),
            .I(N__6202));
    InMux I__1076 (
            .O(N__6205),
            .I(N__6199));
    LocalMux I__1075 (
            .O(N__6202),
            .I(N__6196));
    LocalMux I__1074 (
            .O(N__6199),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    Odrv12 I__1073 (
            .O(N__6196),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__1072 (
            .O(N__6191),
            .I(N__6187));
    InMux I__1071 (
            .O(N__6190),
            .I(N__6184));
    LocalMux I__1070 (
            .O(N__6187),
            .I(N__6181));
    LocalMux I__1069 (
            .O(N__6184),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    Odrv4 I__1068 (
            .O(N__6181),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    CascadeMux I__1067 (
            .O(N__6176),
            .I(N__6173));
    InMux I__1066 (
            .O(N__6173),
            .I(N__6169));
    InMux I__1065 (
            .O(N__6172),
            .I(N__6166));
    LocalMux I__1064 (
            .O(N__6169),
            .I(N__6163));
    LocalMux I__1063 (
            .O(N__6166),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv12 I__1062 (
            .O(N__6163),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__1061 (
            .O(N__6158),
            .I(N__6155));
    LocalMux I__1060 (
            .O(N__6155),
            .I(N__6152));
    Odrv4 I__1059 (
            .O(N__6152),
            .I(\U712_CHIP_RAM.REFRESH5lt7 ));
    CascadeMux I__1058 (
            .O(N__6149),
            .I(N__6144));
    InMux I__1057 (
            .O(N__6148),
            .I(N__6140));
    InMux I__1056 (
            .O(N__6147),
            .I(N__6137));
    InMux I__1055 (
            .O(N__6144),
            .I(N__6134));
    InMux I__1054 (
            .O(N__6143),
            .I(N__6130));
    LocalMux I__1053 (
            .O(N__6140),
            .I(N__6127));
    LocalMux I__1052 (
            .O(N__6137),
            .I(N__6123));
    LocalMux I__1051 (
            .O(N__6134),
            .I(N__6120));
    InMux I__1050 (
            .O(N__6133),
            .I(N__6117));
    LocalMux I__1049 (
            .O(N__6130),
            .I(N__6112));
    Span4Mux_v I__1048 (
            .O(N__6127),
            .I(N__6112));
    InMux I__1047 (
            .O(N__6126),
            .I(N__6109));
    Span4Mux_h I__1046 (
            .O(N__6123),
            .I(N__6106));
    Span4Mux_h I__1045 (
            .O(N__6120),
            .I(N__6101));
    LocalMux I__1044 (
            .O(N__6117),
            .I(N__6101));
    Odrv4 I__1043 (
            .O(N__6112),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__1042 (
            .O(N__6109),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__1041 (
            .O(N__6106),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    Odrv4 I__1040 (
            .O(N__6101),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    InMux I__1039 (
            .O(N__6092),
            .I(N__6089));
    LocalMux I__1038 (
            .O(N__6089),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ));
    InMux I__1037 (
            .O(N__6086),
            .I(N__6083));
    LocalMux I__1036 (
            .O(N__6083),
            .I(N__6079));
    InMux I__1035 (
            .O(N__6082),
            .I(N__6076));
    Odrv4 I__1034 (
            .O(N__6079),
            .I(LATCH_RAM));
    LocalMux I__1033 (
            .O(N__6076),
            .I(LATCH_RAM));
    InMux I__1032 (
            .O(N__6071),
            .I(N__6068));
    LocalMux I__1031 (
            .O(N__6068),
            .I(N__6064));
    InMux I__1030 (
            .O(N__6067),
            .I(N__6061));
    Odrv12 I__1029 (
            .O(N__6064),
            .I(\U712_REG_SM.N_265 ));
    LocalMux I__1028 (
            .O(N__6061),
            .I(\U712_REG_SM.N_265 ));
    InMux I__1027 (
            .O(N__6056),
            .I(N__6053));
    LocalMux I__1026 (
            .O(N__6053),
            .I(N__6050));
    Span4Mux_h I__1025 (
            .O(N__6050),
            .I(N__6044));
    InMux I__1024 (
            .O(N__6049),
            .I(N__6041));
    InMux I__1023 (
            .O(N__6048),
            .I(N__6038));
    InMux I__1022 (
            .O(N__6047),
            .I(N__6035));
    Odrv4 I__1021 (
            .O(N__6044),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_1 ));
    LocalMux I__1020 (
            .O(N__6041),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_1 ));
    LocalMux I__1019 (
            .O(N__6038),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_1 ));
    LocalMux I__1018 (
            .O(N__6035),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_1 ));
    InMux I__1017 (
            .O(N__6026),
            .I(N__6019));
    InMux I__1016 (
            .O(N__6025),
            .I(N__6016));
    CascadeMux I__1015 (
            .O(N__6024),
            .I(N__6013));
    InMux I__1014 (
            .O(N__6023),
            .I(N__6008));
    InMux I__1013 (
            .O(N__6022),
            .I(N__6005));
    LocalMux I__1012 (
            .O(N__6019),
            .I(N__6000));
    LocalMux I__1011 (
            .O(N__6016),
            .I(N__6000));
    InMux I__1010 (
            .O(N__6013),
            .I(N__5994));
    InMux I__1009 (
            .O(N__6012),
            .I(N__5991));
    InMux I__1008 (
            .O(N__6011),
            .I(N__5988));
    LocalMux I__1007 (
            .O(N__6008),
            .I(N__5983));
    LocalMux I__1006 (
            .O(N__6005),
            .I(N__5983));
    Span4Mux_h I__1005 (
            .O(N__6000),
            .I(N__5980));
    InMux I__1004 (
            .O(N__5999),
            .I(N__5973));
    InMux I__1003 (
            .O(N__5998),
            .I(N__5973));
    InMux I__1002 (
            .O(N__5997),
            .I(N__5973));
    LocalMux I__1001 (
            .O(N__5994),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    LocalMux I__1000 (
            .O(N__5991),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    LocalMux I__999 (
            .O(N__5988),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    Odrv4 I__998 (
            .O(N__5983),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    Odrv4 I__997 (
            .O(N__5980),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    LocalMux I__996 (
            .O(N__5973),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_2 ));
    InMux I__995 (
            .O(N__5960),
            .I(N__5955));
    InMux I__994 (
            .O(N__5959),
            .I(N__5952));
    InMux I__993 (
            .O(N__5958),
            .I(N__5949));
    LocalMux I__992 (
            .O(N__5955),
            .I(\U712_REG_SM.DBR_SYNCZ0Z_1 ));
    LocalMux I__991 (
            .O(N__5952),
            .I(\U712_REG_SM.DBR_SYNCZ0Z_1 ));
    LocalMux I__990 (
            .O(N__5949),
            .I(\U712_REG_SM.DBR_SYNCZ0Z_1 ));
    InMux I__989 (
            .O(N__5942),
            .I(N__5939));
    LocalMux I__988 (
            .O(N__5939),
            .I(N__5935));
    InMux I__987 (
            .O(N__5938),
            .I(N__5932));
    Span4Mux_v I__986 (
            .O(N__5935),
            .I(N__5926));
    LocalMux I__985 (
            .O(N__5932),
            .I(N__5926));
    InMux I__984 (
            .O(N__5931),
            .I(N__5923));
    Span4Mux_h I__983 (
            .O(N__5926),
            .I(N__5918));
    LocalMux I__982 (
            .O(N__5923),
            .I(N__5918));
    Span4Mux_v I__981 (
            .O(N__5918),
            .I(N__5915));
    Sp12to4 I__980 (
            .O(N__5915),
            .I(N__5912));
    Span12Mux_h I__979 (
            .O(N__5912),
            .I(N__5909));
    Odrv12 I__978 (
            .O(N__5909),
            .I(DBRn_c));
    InMux I__977 (
            .O(N__5906),
            .I(N__5903));
    LocalMux I__976 (
            .O(N__5903),
            .I(\U712_REG_SM.DBR_SYNCZ0Z_0 ));
    InMux I__975 (
            .O(N__5900),
            .I(N__5897));
    LocalMux I__974 (
            .O(N__5897),
            .I(N__5894));
    Span4Mux_v I__973 (
            .O(N__5894),
            .I(N__5886));
    InMux I__972 (
            .O(N__5893),
            .I(N__5881));
    InMux I__971 (
            .O(N__5892),
            .I(N__5881));
    InMux I__970 (
            .O(N__5891),
            .I(N__5874));
    InMux I__969 (
            .O(N__5890),
            .I(N__5874));
    InMux I__968 (
            .O(N__5889),
            .I(N__5874));
    Odrv4 I__967 (
            .O(N__5886),
            .I(REG_WRITE_CYCLE));
    LocalMux I__966 (
            .O(N__5881),
            .I(REG_WRITE_CYCLE));
    LocalMux I__965 (
            .O(N__5874),
            .I(REG_WRITE_CYCLE));
    IoInMux I__964 (
            .O(N__5867),
            .I(N__5864));
    LocalMux I__963 (
            .O(N__5864),
            .I(N__5860));
    IoInMux I__962 (
            .O(N__5863),
            .I(N__5857));
    IoSpan4Mux I__961 (
            .O(N__5860),
            .I(N__5854));
    LocalMux I__960 (
            .O(N__5857),
            .I(N__5851));
    Span4Mux_s3_h I__959 (
            .O(N__5854),
            .I(N__5848));
    IoSpan4Mux I__958 (
            .O(N__5851),
            .I(N__5845));
    Span4Mux_h I__957 (
            .O(N__5848),
            .I(N__5842));
    Span4Mux_s2_v I__956 (
            .O(N__5845),
            .I(N__5839));
    Sp12to4 I__955 (
            .O(N__5842),
            .I(N__5836));
    Sp12to4 I__954 (
            .O(N__5839),
            .I(N__5833));
    Span12Mux_h I__953 (
            .O(N__5836),
            .I(N__5830));
    Span12Mux_s10_v I__952 (
            .O(N__5833),
            .I(N__5827));
    Odrv12 I__951 (
            .O(N__5830),
            .I(N_289));
    Odrv12 I__950 (
            .O(N__5827),
            .I(N_289));
    InMux I__949 (
            .O(N__5822),
            .I(N__5819));
    LocalMux I__948 (
            .O(N__5819),
            .I(N__5816));
    Sp12to4 I__947 (
            .O(N__5816),
            .I(N__5813));
    Span12Mux_v I__946 (
            .O(N__5813),
            .I(N__5810));
    Span12Mux_h I__945 (
            .O(N__5810),
            .I(N__5807));
    Odrv12 I__944 (
            .O(N__5807),
            .I(A_c_5));
    InMux I__943 (
            .O(N__5804),
            .I(N__5801));
    LocalMux I__942 (
            .O(N__5801),
            .I(N__5798));
    Span4Mux_v I__941 (
            .O(N__5798),
            .I(N__5795));
    Sp12to4 I__940 (
            .O(N__5795),
            .I(N__5792));
    Span12Mux_h I__939 (
            .O(N__5792),
            .I(N__5789));
    Odrv12 I__938 (
            .O(N__5789),
            .I(A_c_12));
    CascadeMux I__937 (
            .O(N__5786),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ));
    InMux I__936 (
            .O(N__5783),
            .I(N__5780));
    LocalMux I__935 (
            .O(N__5780),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ));
    CascadeMux I__934 (
            .O(N__5777),
            .I(\U712_CHIP_RAM.N_365_1_cascade_ ));
    CascadeMux I__933 (
            .O(N__5774),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_ ));
    CEMux I__932 (
            .O(N__5771),
            .I(N__5768));
    LocalMux I__931 (
            .O(N__5768),
            .I(N__5765));
    Span4Mux_h I__930 (
            .O(N__5765),
            .I(N__5762));
    Odrv4 I__929 (
            .O(N__5762),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0 ));
    InMux I__928 (
            .O(N__5759),
            .I(N__5753));
    CascadeMux I__927 (
            .O(N__5758),
            .I(N__5750));
    InMux I__926 (
            .O(N__5757),
            .I(N__5747));
    InMux I__925 (
            .O(N__5756),
            .I(N__5744));
    LocalMux I__924 (
            .O(N__5753),
            .I(N__5741));
    InMux I__923 (
            .O(N__5750),
            .I(N__5738));
    LocalMux I__922 (
            .O(N__5747),
            .I(N__5735));
    LocalMux I__921 (
            .O(N__5744),
            .I(N__5732));
    Span4Mux_h I__920 (
            .O(N__5741),
            .I(N__5727));
    LocalMux I__919 (
            .O(N__5738),
            .I(N__5727));
    Sp12to4 I__918 (
            .O(N__5735),
            .I(N__5724));
    Span4Mux_v I__917 (
            .O(N__5732),
            .I(N__5719));
    Span4Mux_v I__916 (
            .O(N__5727),
            .I(N__5719));
    Span12Mux_v I__915 (
            .O(N__5724),
            .I(N__5716));
    Sp12to4 I__914 (
            .O(N__5719),
            .I(N__5713));
    Span12Mux_h I__913 (
            .O(N__5716),
            .I(N__5710));
    Span12Mux_h I__912 (
            .O(N__5713),
            .I(N__5707));
    Odrv12 I__911 (
            .O(N__5710),
            .I(RnW_c));
    Odrv12 I__910 (
            .O(N__5707),
            .I(RnW_c));
    IoInMux I__909 (
            .O(N__5702),
            .I(N__5699));
    LocalMux I__908 (
            .O(N__5699),
            .I(N__5696));
    IoSpan4Mux I__907 (
            .O(N__5696),
            .I(N__5693));
    Span4Mux_s3_h I__906 (
            .O(N__5693),
            .I(N__5690));
    Span4Mux_h I__905 (
            .O(N__5690),
            .I(N__5687));
    Sp12to4 I__904 (
            .O(N__5687),
            .I(N__5684));
    Span12Mux_h I__903 (
            .O(N__5684),
            .I(N__5680));
    InMux I__902 (
            .O(N__5683),
            .I(N__5677));
    Odrv12 I__901 (
            .O(N__5680),
            .I(CLK_EN_c));
    LocalMux I__900 (
            .O(N__5677),
            .I(CLK_EN_c));
    InMux I__899 (
            .O(N__5672),
            .I(N__5669));
    LocalMux I__898 (
            .O(N__5669),
            .I(N__5666));
    Span12Mux_h I__897 (
            .O(N__5666),
            .I(N__5663));
    Span12Mux_v I__896 (
            .O(N__5663),
            .I(N__5660));
    Odrv12 I__895 (
            .O(N__5660),
            .I(RAMSPACEn_c));
    CascadeMux I__894 (
            .O(N__5657),
            .I(N__5654));
    InMux I__893 (
            .O(N__5654),
            .I(N__5650));
    CascadeMux I__892 (
            .O(N__5653),
            .I(N__5647));
    LocalMux I__891 (
            .O(N__5650),
            .I(N__5644));
    InMux I__890 (
            .O(N__5647),
            .I(N__5641));
    Span4Mux_h I__889 (
            .O(N__5644),
            .I(N__5636));
    LocalMux I__888 (
            .O(N__5641),
            .I(N__5636));
    Span4Mux_v I__887 (
            .O(N__5636),
            .I(N__5633));
    Sp12to4 I__886 (
            .O(N__5633),
            .I(N__5630));
    Span12Mux_h I__885 (
            .O(N__5630),
            .I(N__5627));
    Odrv12 I__884 (
            .O(N__5627),
            .I(TSn_c));
    InMux I__883 (
            .O(N__5624),
            .I(N__5617));
    CascadeMux I__882 (
            .O(N__5623),
            .I(N__5614));
    InMux I__881 (
            .O(N__5622),
            .I(N__5611));
    InMux I__880 (
            .O(N__5621),
            .I(N__5608));
    InMux I__879 (
            .O(N__5620),
            .I(N__5605));
    LocalMux I__878 (
            .O(N__5617),
            .I(N__5602));
    InMux I__877 (
            .O(N__5614),
            .I(N__5599));
    LocalMux I__876 (
            .O(N__5611),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__875 (
            .O(N__5608),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__874 (
            .O(N__5605),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv4 I__873 (
            .O(N__5602),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__872 (
            .O(N__5599),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__871 (
            .O(N__5588),
            .I(N__5584));
    InMux I__870 (
            .O(N__5587),
            .I(N__5579));
    LocalMux I__869 (
            .O(N__5584),
            .I(N__5576));
    InMux I__868 (
            .O(N__5583),
            .I(N__5573));
    InMux I__867 (
            .O(N__5582),
            .I(N__5570));
    LocalMux I__866 (
            .O(N__5579),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__865 (
            .O(N__5576),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__864 (
            .O(N__5573),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__863 (
            .O(N__5570),
            .I(DBR_SYNCZ0Z_1));
    InMux I__862 (
            .O(N__5561),
            .I(N__5558));
    LocalMux I__861 (
            .O(N__5558),
            .I(DBR_SYNCZ0Z_0));
    CascadeMux I__860 (
            .O(N__5555),
            .I(\U712_CHIP_RAM.N_376_cascade_ ));
    CascadeMux I__859 (
            .O(N__5552),
            .I(\U712_CHIP_RAM.N_45_i_cascade_ ));
    InMux I__858 (
            .O(N__5549),
            .I(N__5546));
    LocalMux I__857 (
            .O(N__5546),
            .I(\U712_CHIP_RAM.N_324_2 ));
    CascadeMux I__856 (
            .O(N__5543),
            .I(\U712_CHIP_RAM.N_324_2_cascade_ ));
    CascadeMux I__855 (
            .O(N__5540),
            .I(N__5537));
    InMux I__854 (
            .O(N__5537),
            .I(N__5532));
    InMux I__853 (
            .O(N__5536),
            .I(N__5529));
    InMux I__852 (
            .O(N__5535),
            .I(N__5526));
    LocalMux I__851 (
            .O(N__5532),
            .I(\U712_CHIP_RAM.N_450 ));
    LocalMux I__850 (
            .O(N__5529),
            .I(\U712_CHIP_RAM.N_450 ));
    LocalMux I__849 (
            .O(N__5526),
            .I(\U712_CHIP_RAM.N_450 ));
    InMux I__848 (
            .O(N__5519),
            .I(N__5515));
    InMux I__847 (
            .O(N__5518),
            .I(N__5512));
    LocalMux I__846 (
            .O(N__5515),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVCZ0Z_4 ));
    LocalMux I__845 (
            .O(N__5512),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVCZ0Z_4 ));
    InMux I__844 (
            .O(N__5507),
            .I(N__5504));
    LocalMux I__843 (
            .O(N__5504),
            .I(\U712_CHIP_RAM.N_252 ));
    CascadeMux I__842 (
            .O(N__5501),
            .I(\U712_CHIP_RAM.N_252_cascade_ ));
    CascadeMux I__841 (
            .O(N__5498),
            .I(\U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ));
    InMux I__840 (
            .O(N__5495),
            .I(N__5492));
    LocalMux I__839 (
            .O(N__5492),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ));
    InMux I__838 (
            .O(N__5489),
            .I(N__5486));
    LocalMux I__837 (
            .O(N__5486),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_1 ));
    CascadeMux I__836 (
            .O(N__5483),
            .I(\U712_CHIP_RAM.N_325_cascade_ ));
    InMux I__835 (
            .O(N__5480),
            .I(N__5477));
    LocalMux I__834 (
            .O(N__5477),
            .I(N__5474));
    Span4Mux_v I__833 (
            .O(N__5474),
            .I(N__5471));
    Odrv4 I__832 (
            .O(N__5471),
            .I(\U712_CHIP_RAM.N_301 ));
    CascadeMux I__831 (
            .O(N__5468),
            .I(\U712_CHIP_RAM.N_392_cascade_ ));
    InMux I__830 (
            .O(N__5465),
            .I(N__5462));
    LocalMux I__829 (
            .O(N__5462),
            .I(\U712_CHIP_RAM.N_449 ));
    InMux I__828 (
            .O(N__5459),
            .I(N__5456));
    LocalMux I__827 (
            .O(N__5456),
            .I(N__5453));
    Span4Mux_h I__826 (
            .O(N__5453),
            .I(N__5450));
    Span4Mux_v I__825 (
            .O(N__5450),
            .I(N__5447));
    Sp12to4 I__824 (
            .O(N__5447),
            .I(N__5444));
    Odrv12 I__823 (
            .O(N__5444),
            .I(A_c_8));
    InMux I__822 (
            .O(N__5441),
            .I(N__5438));
    LocalMux I__821 (
            .O(N__5438),
            .I(N__5435));
    Span4Mux_v I__820 (
            .O(N__5435),
            .I(N__5432));
    Span4Mux_v I__819 (
            .O(N__5432),
            .I(N__5429));
    Sp12to4 I__818 (
            .O(N__5429),
            .I(N__5426));
    Span12Mux_h I__817 (
            .O(N__5426),
            .I(N__5423));
    Odrv12 I__816 (
            .O(N__5423),
            .I(A_c_15));
    CascadeMux I__815 (
            .O(N__5420),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ));
    InMux I__814 (
            .O(N__5417),
            .I(N__5414));
    LocalMux I__813 (
            .O(N__5414),
            .I(N__5411));
    Span4Mux_v I__812 (
            .O(N__5411),
            .I(N__5408));
    Sp12to4 I__811 (
            .O(N__5408),
            .I(N__5405));
    Span12Mux_h I__810 (
            .O(N__5405),
            .I(N__5402));
    Odrv12 I__809 (
            .O(N__5402),
            .I(A_c_13));
    InMux I__808 (
            .O(N__5399),
            .I(N__5396));
    LocalMux I__807 (
            .O(N__5396),
            .I(N__5393));
    Span12Mux_v I__806 (
            .O(N__5393),
            .I(N__5390));
    Span12Mux_h I__805 (
            .O(N__5390),
            .I(N__5387));
    Odrv12 I__804 (
            .O(N__5387),
            .I(A_c_6));
    InMux I__803 (
            .O(N__5384),
            .I(N__5381));
    LocalMux I__802 (
            .O(N__5381),
            .I(N__5378));
    Span12Mux_v I__801 (
            .O(N__5378),
            .I(N__5375));
    Span12Mux_h I__800 (
            .O(N__5375),
            .I(N__5372));
    Odrv12 I__799 (
            .O(N__5372),
            .I(A_c_16));
    InMux I__798 (
            .O(N__5369),
            .I(N__5366));
    LocalMux I__797 (
            .O(N__5366),
            .I(N__5363));
    Span12Mux_v I__796 (
            .O(N__5363),
            .I(N__5360));
    Span12Mux_h I__795 (
            .O(N__5360),
            .I(N__5357));
    Odrv12 I__794 (
            .O(N__5357),
            .I(A_c_18));
    CascadeMux I__793 (
            .O(N__5354),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5_cascade_ ));
    InMux I__792 (
            .O(N__5351),
            .I(N__5348));
    LocalMux I__791 (
            .O(N__5348),
            .I(N__5345));
    Odrv4 I__790 (
            .O(N__5345),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ));
    IoInMux I__789 (
            .O(N__5342),
            .I(N__5339));
    LocalMux I__788 (
            .O(N__5339),
            .I(N__5336));
    IoSpan4Mux I__787 (
            .O(N__5336),
            .I(N__5333));
    Sp12to4 I__786 (
            .O(N__5333),
            .I(N__5330));
    Span12Mux_s7_h I__785 (
            .O(N__5330),
            .I(N__5327));
    Span12Mux_v I__784 (
            .O(N__5327),
            .I(N__5324));
    Odrv12 I__783 (
            .O(N__5324),
            .I(CMA_c_5));
    InMux I__782 (
            .O(N__5321),
            .I(N__5318));
    LocalMux I__781 (
            .O(N__5318),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    IoInMux I__780 (
            .O(N__5315),
            .I(N__5312));
    LocalMux I__779 (
            .O(N__5312),
            .I(N__5309));
    Span4Mux_s1_v I__778 (
            .O(N__5309),
            .I(N__5306));
    Span4Mux_v I__777 (
            .O(N__5306),
            .I(N__5303));
    Span4Mux_v I__776 (
            .O(N__5303),
            .I(N__5300));
    Span4Mux_v I__775 (
            .O(N__5300),
            .I(N__5297));
    Odrv4 I__774 (
            .O(N__5297),
            .I(CMA_c_1));
    InMux I__773 (
            .O(N__5294),
            .I(N__5291));
    LocalMux I__772 (
            .O(N__5291),
            .I(\U712_CHIP_RAM.un1_CMA28_0_i ));
    InMux I__771 (
            .O(N__5288),
            .I(N__5285));
    LocalMux I__770 (
            .O(N__5285),
            .I(N__5282));
    Span4Mux_v I__769 (
            .O(N__5282),
            .I(N__5279));
    Sp12to4 I__768 (
            .O(N__5279),
            .I(N__5276));
    Span12Mux_h I__767 (
            .O(N__5276),
            .I(N__5273));
    Odrv12 I__766 (
            .O(N__5273),
            .I(A_c_11));
    InMux I__765 (
            .O(N__5270),
            .I(N__5267));
    LocalMux I__764 (
            .O(N__5267),
            .I(N__5264));
    Span12Mux_v I__763 (
            .O(N__5264),
            .I(N__5261));
    Span12Mux_h I__762 (
            .O(N__5261),
            .I(N__5258));
    Odrv12 I__761 (
            .O(N__5258),
            .I(A_c_4));
    InMux I__760 (
            .O(N__5255),
            .I(N__5250));
    InMux I__759 (
            .O(N__5254),
            .I(N__5247));
    InMux I__758 (
            .O(N__5253),
            .I(N__5244));
    LocalMux I__757 (
            .O(N__5250),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_7 ));
    LocalMux I__756 (
            .O(N__5247),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_7 ));
    LocalMux I__755 (
            .O(N__5244),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_7 ));
    CascadeMux I__754 (
            .O(N__5237),
            .I(N__5234));
    InMux I__753 (
            .O(N__5234),
            .I(N__5228));
    InMux I__752 (
            .O(N__5233),
            .I(N__5221));
    InMux I__751 (
            .O(N__5232),
            .I(N__5221));
    InMux I__750 (
            .O(N__5231),
            .I(N__5221));
    LocalMux I__749 (
            .O(N__5228),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_3 ));
    LocalMux I__748 (
            .O(N__5221),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_3 ));
    CascadeMux I__747 (
            .O(N__5216),
            .I(\U712_REG_SM.un18_0_i_0_0_1_cascade_ ));
    CascadeMux I__746 (
            .O(N__5213),
            .I(N__5209));
    CascadeMux I__745 (
            .O(N__5212),
            .I(N__5203));
    InMux I__744 (
            .O(N__5209),
            .I(N__5198));
    InMux I__743 (
            .O(N__5208),
            .I(N__5195));
    InMux I__742 (
            .O(N__5207),
            .I(N__5188));
    InMux I__741 (
            .O(N__5206),
            .I(N__5188));
    InMux I__740 (
            .O(N__5203),
            .I(N__5188));
    InMux I__739 (
            .O(N__5202),
            .I(N__5185));
    InMux I__738 (
            .O(N__5201),
            .I(N__5182));
    LocalMux I__737 (
            .O(N__5198),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_8 ));
    LocalMux I__736 (
            .O(N__5195),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_8 ));
    LocalMux I__735 (
            .O(N__5188),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_8 ));
    LocalMux I__734 (
            .O(N__5185),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_8 ));
    LocalMux I__733 (
            .O(N__5182),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_8 ));
    InMux I__732 (
            .O(N__5171),
            .I(N__5167));
    InMux I__731 (
            .O(N__5170),
            .I(N__5162));
    LocalMux I__730 (
            .O(N__5167),
            .I(N__5159));
    InMux I__729 (
            .O(N__5166),
            .I(N__5154));
    InMux I__728 (
            .O(N__5165),
            .I(N__5154));
    LocalMux I__727 (
            .O(N__5162),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_4 ));
    Odrv4 I__726 (
            .O(N__5159),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_4 ));
    LocalMux I__725 (
            .O(N__5154),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_4 ));
    CascadeMux I__724 (
            .O(N__5147),
            .I(\U712_REG_SM.N_442_cascade_ ));
    CascadeMux I__723 (
            .O(N__5144),
            .I(N__5141));
    InMux I__722 (
            .O(N__5141),
            .I(N__5138));
    LocalMux I__721 (
            .O(N__5138),
            .I(N__5135));
    Odrv4 I__720 (
            .O(N__5135),
            .I(\U712_REG_SM.REG_CPU_CYCLE_e_1 ));
    InMux I__719 (
            .O(N__5132),
            .I(N__5129));
    LocalMux I__718 (
            .O(N__5129),
            .I(\U712_REG_SM.N_84 ));
    CascadeMux I__717 (
            .O(N__5126),
            .I(N__5120));
    CascadeMux I__716 (
            .O(N__5125),
            .I(N__5115));
    CascadeMux I__715 (
            .O(N__5124),
            .I(N__5109));
    InMux I__714 (
            .O(N__5123),
            .I(N__5105));
    InMux I__713 (
            .O(N__5120),
            .I(N__5102));
    InMux I__712 (
            .O(N__5119),
            .I(N__5099));
    InMux I__711 (
            .O(N__5118),
            .I(N__5094));
    InMux I__710 (
            .O(N__5115),
            .I(N__5094));
    InMux I__709 (
            .O(N__5114),
            .I(N__5091));
    InMux I__708 (
            .O(N__5113),
            .I(N__5084));
    InMux I__707 (
            .O(N__5112),
            .I(N__5084));
    InMux I__706 (
            .O(N__5109),
            .I(N__5084));
    InMux I__705 (
            .O(N__5108),
            .I(N__5081));
    LocalMux I__704 (
            .O(N__5105),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__703 (
            .O(N__5102),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__702 (
            .O(N__5099),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__701 (
            .O(N__5094),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__700 (
            .O(N__5091),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__699 (
            .O(N__5084),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__698 (
            .O(N__5081),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    CascadeMux I__697 (
            .O(N__5066),
            .I(N__5059));
    CascadeMux I__696 (
            .O(N__5065),
            .I(N__5055));
    CascadeMux I__695 (
            .O(N__5064),
            .I(N__5050));
    CascadeMux I__694 (
            .O(N__5063),
            .I(N__5047));
    InMux I__693 (
            .O(N__5062),
            .I(N__5042));
    InMux I__692 (
            .O(N__5059),
            .I(N__5039));
    InMux I__691 (
            .O(N__5058),
            .I(N__5036));
    InMux I__690 (
            .O(N__5055),
            .I(N__5031));
    InMux I__689 (
            .O(N__5054),
            .I(N__5031));
    InMux I__688 (
            .O(N__5053),
            .I(N__5028));
    InMux I__687 (
            .O(N__5050),
            .I(N__5025));
    InMux I__686 (
            .O(N__5047),
            .I(N__5020));
    InMux I__685 (
            .O(N__5046),
            .I(N__5020));
    InMux I__684 (
            .O(N__5045),
            .I(N__5017));
    LocalMux I__683 (
            .O(N__5042),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__682 (
            .O(N__5039),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__681 (
            .O(N__5036),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__680 (
            .O(N__5031),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__679 (
            .O(N__5028),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__678 (
            .O(N__5025),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__677 (
            .O(N__5020),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__676 (
            .O(N__5017),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__675 (
            .O(N__5000),
            .I(N__4995));
    InMux I__674 (
            .O(N__4999),
            .I(N__4992));
    InMux I__673 (
            .O(N__4998),
            .I(N__4989));
    LocalMux I__672 (
            .O(N__4995),
            .I(\U712_REG_SM.N_447 ));
    LocalMux I__671 (
            .O(N__4992),
            .I(\U712_REG_SM.N_447 ));
    LocalMux I__670 (
            .O(N__4989),
            .I(\U712_REG_SM.N_447 ));
    InMux I__669 (
            .O(N__4982),
            .I(N__4976));
    InMux I__668 (
            .O(N__4981),
            .I(N__4973));
    InMux I__667 (
            .O(N__4980),
            .I(N__4968));
    InMux I__666 (
            .O(N__4979),
            .I(N__4968));
    LocalMux I__665 (
            .O(N__4976),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_6 ));
    LocalMux I__664 (
            .O(N__4973),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_6 ));
    LocalMux I__663 (
            .O(N__4968),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_6 ));
    InMux I__662 (
            .O(N__4961),
            .I(N__4958));
    LocalMux I__661 (
            .O(N__4958),
            .I(\U712_REG_SM.N_288 ));
    InMux I__660 (
            .O(N__4955),
            .I(N__4951));
    InMux I__659 (
            .O(N__4954),
            .I(N__4948));
    LocalMux I__658 (
            .O(N__4951),
            .I(LATCH_REG));
    LocalMux I__657 (
            .O(N__4948),
            .I(LATCH_REG));
    IoInMux I__656 (
            .O(N__4943),
            .I(N__4940));
    LocalMux I__655 (
            .O(N__4940),
            .I(N__4937));
    Span4Mux_s3_v I__654 (
            .O(N__4937),
            .I(N__4934));
    Span4Mux_h I__653 (
            .O(N__4934),
            .I(N__4931));
    Span4Mux_v I__652 (
            .O(N__4931),
            .I(N__4928));
    Span4Mux_v I__651 (
            .O(N__4928),
            .I(N__4925));
    Odrv4 I__650 (
            .O(N__4925),
            .I(LATCH_CLK_0_i));
    CascadeMux I__649 (
            .O(N__4922),
            .I(\U712_CHIP_RAM.N_452_cascade_ ));
    CascadeMux I__648 (
            .O(N__4919),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_ ));
    CEMux I__647 (
            .O(N__4916),
            .I(N__4913));
    LocalMux I__646 (
            .O(N__4913),
            .I(N__4910));
    Odrv12 I__645 (
            .O(N__4910),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0 ));
    IoInMux I__644 (
            .O(N__4907),
            .I(N__4904));
    LocalMux I__643 (
            .O(N__4904),
            .I(N__4901));
    IoSpan4Mux I__642 (
            .O(N__4901),
            .I(N__4898));
    IoSpan4Mux I__641 (
            .O(N__4898),
            .I(N__4895));
    Span4Mux_s1_v I__640 (
            .O(N__4895),
            .I(N__4892));
    Sp12to4 I__639 (
            .O(N__4892),
            .I(N__4889));
    Span12Mux_v I__638 (
            .O(N__4889),
            .I(N__4883));
    InMux I__637 (
            .O(N__4888),
            .I(N__4880));
    InMux I__636 (
            .O(N__4887),
            .I(N__4877));
    InMux I__635 (
            .O(N__4886),
            .I(N__4874));
    Odrv12 I__634 (
            .O(N__4883),
            .I(LDSn_c));
    LocalMux I__633 (
            .O(N__4880),
            .I(LDSn_c));
    LocalMux I__632 (
            .O(N__4877),
            .I(LDSn_c));
    LocalMux I__631 (
            .O(N__4874),
            .I(LDSn_c));
    InMux I__630 (
            .O(N__4865),
            .I(N__4856));
    InMux I__629 (
            .O(N__4864),
            .I(N__4856));
    InMux I__628 (
            .O(N__4863),
            .I(N__4853));
    InMux I__627 (
            .O(N__4862),
            .I(N__4850));
    InMux I__626 (
            .O(N__4861),
            .I(N__4847));
    LocalMux I__625 (
            .O(N__4856),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    LocalMux I__624 (
            .O(N__4853),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    LocalMux I__623 (
            .O(N__4850),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    LocalMux I__622 (
            .O(N__4847),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_0 ));
    InMux I__621 (
            .O(N__4838),
            .I(N__4835));
    LocalMux I__620 (
            .O(N__4835),
            .I(\U712_REG_SM.N_309 ));
    InMux I__619 (
            .O(N__4832),
            .I(N__4829));
    LocalMux I__618 (
            .O(N__4829),
            .I(\U712_REG_SM.STATE_COUNTER_srsts_i_i_i_a3_2_0 ));
    CascadeMux I__617 (
            .O(N__4826),
            .I(N__4822));
    InMux I__616 (
            .O(N__4825),
            .I(N__4817));
    InMux I__615 (
            .O(N__4822),
            .I(N__4817));
    LocalMux I__614 (
            .O(N__4817),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_5 ));
    SRMux I__613 (
            .O(N__4814),
            .I(N__4811));
    LocalMux I__612 (
            .O(N__4811),
            .I(N__4808));
    Odrv4 I__611 (
            .O(N__4808),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    InMux I__610 (
            .O(N__4805),
            .I(N__4802));
    LocalMux I__609 (
            .O(N__4802),
            .I(N__4799));
    Span4Mux_v I__608 (
            .O(N__4799),
            .I(N__4796));
    Span4Mux_h I__607 (
            .O(N__4796),
            .I(N__4793));
    Sp12to4 I__606 (
            .O(N__4793),
            .I(N__4790));
    Span12Mux_v I__605 (
            .O(N__4790),
            .I(N__4787));
    Odrv12 I__604 (
            .O(N__4787),
            .I(A_c_14));
    InMux I__603 (
            .O(N__4784),
            .I(N__4781));
    LocalMux I__602 (
            .O(N__4781),
            .I(N__4778));
    Span4Mux_v I__601 (
            .O(N__4778),
            .I(N__4775));
    Sp12to4 I__600 (
            .O(N__4775),
            .I(N__4772));
    Odrv12 I__599 (
            .O(N__4772),
            .I(A_c_7));
    CascadeMux I__598 (
            .O(N__4769),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5_cascade_ ));
    IoInMux I__597 (
            .O(N__4766),
            .I(N__4763));
    LocalMux I__596 (
            .O(N__4763),
            .I(N__4760));
    Span12Mux_s1_h I__595 (
            .O(N__4760),
            .I(N__4757));
    Odrv12 I__594 (
            .O(N__4757),
            .I(DBRn_c_i_0));
    InMux I__593 (
            .O(N__4754),
            .I(N__4751));
    LocalMux I__592 (
            .O(N__4751),
            .I(N__4748));
    Span4Mux_h I__591 (
            .O(N__4748),
            .I(N__4745));
    Span4Mux_v I__590 (
            .O(N__4745),
            .I(N__4742));
    Sp12to4 I__589 (
            .O(N__4742),
            .I(N__4739));
    Odrv12 I__588 (
            .O(N__4739),
            .I(A_c_20));
    CascadeMux I__587 (
            .O(N__4736),
            .I(\U712_CHIP_RAM.N_361_cascade_ ));
    IoInMux I__586 (
            .O(N__4733),
            .I(N__4730));
    LocalMux I__585 (
            .O(N__4730),
            .I(N__4727));
    Span4Mux_s3_v I__584 (
            .O(N__4727),
            .I(N__4724));
    Span4Mux_h I__583 (
            .O(N__4724),
            .I(N__4721));
    Sp12to4 I__582 (
            .O(N__4721),
            .I(N__4718));
    Span12Mux_v I__581 (
            .O(N__4718),
            .I(N__4715));
    Odrv12 I__580 (
            .O(N__4715),
            .I(BANK0_c));
    InMux I__579 (
            .O(N__4712),
            .I(N__4709));
    LocalMux I__578 (
            .O(N__4709),
            .I(\U712_CHIP_RAM.N_452 ));
    InMux I__577 (
            .O(N__4706),
            .I(N__4703));
    LocalMux I__576 (
            .O(N__4703),
            .I(N__4700));
    Odrv4 I__575 (
            .O(N__4700),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__574 (
            .O(N__4697),
            .I(N__4693));
    IoInMux I__573 (
            .O(N__4696),
            .I(N__4690));
    LocalMux I__572 (
            .O(N__4693),
            .I(N__4687));
    LocalMux I__571 (
            .O(N__4690),
            .I(N__4684));
    Span4Mux_v I__570 (
            .O(N__4687),
            .I(N__4681));
    IoSpan4Mux I__569 (
            .O(N__4684),
            .I(N__4678));
    Sp12to4 I__568 (
            .O(N__4681),
            .I(N__4675));
    IoSpan4Mux I__567 (
            .O(N__4678),
            .I(N__4672));
    Span12Mux_h I__566 (
            .O(N__4675),
            .I(N__4669));
    IoSpan4Mux I__565 (
            .O(N__4672),
            .I(N__4666));
    Odrv12 I__564 (
            .O(N__4669),
            .I(C1_c));
    Odrv4 I__563 (
            .O(N__4666),
            .I(C1_c));
    InMux I__562 (
            .O(N__4661),
            .I(N__4658));
    LocalMux I__561 (
            .O(N__4658),
            .I(N__4655));
    Odrv4 I__560 (
            .O(N__4655),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    InMux I__559 (
            .O(N__4652),
            .I(N__4649));
    LocalMux I__558 (
            .O(N__4649),
            .I(N__4646));
    Sp12to4 I__557 (
            .O(N__4646),
            .I(N__4643));
    Span12Mux_v I__556 (
            .O(N__4643),
            .I(N__4640));
    Span12Mux_h I__555 (
            .O(N__4640),
            .I(N__4637));
    Odrv12 I__554 (
            .O(N__4637),
            .I(A_c_3));
    CascadeMux I__553 (
            .O(N__4634),
            .I(\U712_CHIP_RAM.N_241_cascade_ ));
    InMux I__552 (
            .O(N__4631),
            .I(N__4628));
    LocalMux I__551 (
            .O(N__4628),
            .I(\U712_BYTE_ENABLE.N_276 ));
    CascadeMux I__550 (
            .O(N__4625),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0_cascade_ ));
    IoInMux I__549 (
            .O(N__4622),
            .I(N__4619));
    LocalMux I__548 (
            .O(N__4619),
            .I(N__4616));
    Span4Mux_s2_v I__547 (
            .O(N__4616),
            .I(N__4613));
    Span4Mux_v I__546 (
            .O(N__4613),
            .I(N__4610));
    Span4Mux_v I__545 (
            .O(N__4610),
            .I(N__4607));
    Span4Mux_v I__544 (
            .O(N__4607),
            .I(N__4604));
    Odrv4 I__543 (
            .O(N__4604),
            .I(N_47_i));
    InMux I__542 (
            .O(N__4601),
            .I(N__4597));
    InMux I__541 (
            .O(N__4600),
            .I(N__4594));
    LocalMux I__540 (
            .O(N__4597),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__539 (
            .O(N__4594),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__538 (
            .O(N__4589),
            .I(N__4585));
    InMux I__537 (
            .O(N__4588),
            .I(N__4582));
    LocalMux I__536 (
            .O(N__4585),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__535 (
            .O(N__4582),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    CascadeMux I__534 (
            .O(N__4577),
            .I(N__4573));
    InMux I__533 (
            .O(N__4576),
            .I(N__4570));
    InMux I__532 (
            .O(N__4573),
            .I(N__4567));
    LocalMux I__531 (
            .O(N__4570),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__530 (
            .O(N__4567),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__529 (
            .O(N__4562),
            .I(N__4558));
    InMux I__528 (
            .O(N__4561),
            .I(N__4555));
    LocalMux I__527 (
            .O(N__4558),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__526 (
            .O(N__4555),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__525 (
            .O(N__4550),
            .I(N__4547));
    LocalMux I__524 (
            .O(N__4547),
            .I(\U712_REG_SM.N_266 ));
    CascadeMux I__523 (
            .O(N__4544),
            .I(\U712_REG_SM.STATE_COUNTER_srsts_i_i_i_a3_3_0_cascade_ ));
    InMux I__522 (
            .O(N__4541),
            .I(N__4538));
    LocalMux I__521 (
            .O(N__4538),
            .I(N__4535));
    Span4Mux_v I__520 (
            .O(N__4535),
            .I(N__4532));
    Sp12to4 I__519 (
            .O(N__4532),
            .I(N__4529));
    Span12Mux_h I__518 (
            .O(N__4529),
            .I(N__4526));
    Span12Mux_v I__517 (
            .O(N__4526),
            .I(N__4523));
    Odrv12 I__516 (
            .O(N__4523),
            .I(REGSPACEn_c));
    InMux I__515 (
            .O(N__4520),
            .I(N__4516));
    InMux I__514 (
            .O(N__4519),
            .I(N__4513));
    LocalMux I__513 (
            .O(N__4516),
            .I(\U712_REG_SM.CYCLE_RUNZ0 ));
    LocalMux I__512 (
            .O(N__4513),
            .I(\U712_REG_SM.CYCLE_RUNZ0 ));
    InMux I__511 (
            .O(N__4508),
            .I(N__4502));
    InMux I__510 (
            .O(N__4507),
            .I(N__4497));
    InMux I__509 (
            .O(N__4506),
            .I(N__4497));
    InMux I__508 (
            .O(N__4505),
            .I(N__4494));
    LocalMux I__507 (
            .O(N__4502),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__506 (
            .O(N__4497),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__505 (
            .O(N__4494),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__504 (
            .O(N__4487),
            .I(N__4478));
    InMux I__503 (
            .O(N__4486),
            .I(N__4475));
    InMux I__502 (
            .O(N__4485),
            .I(N__4472));
    InMux I__501 (
            .O(N__4484),
            .I(N__4469));
    InMux I__500 (
            .O(N__4483),
            .I(N__4462));
    InMux I__499 (
            .O(N__4482),
            .I(N__4462));
    InMux I__498 (
            .O(N__4481),
            .I(N__4462));
    LocalMux I__497 (
            .O(N__4478),
            .I(N__4457));
    LocalMux I__496 (
            .O(N__4475),
            .I(N__4457));
    LocalMux I__495 (
            .O(N__4472),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_9 ));
    LocalMux I__494 (
            .O(N__4469),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_9 ));
    LocalMux I__493 (
            .O(N__4462),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_9 ));
    Odrv4 I__492 (
            .O(N__4457),
            .I(\U712_REG_SM.STATE_COUNTERZ0Z_9 ));
    InMux I__491 (
            .O(N__4448),
            .I(N__4443));
    InMux I__490 (
            .O(N__4447),
            .I(N__4438));
    InMux I__489 (
            .O(N__4446),
            .I(N__4438));
    LocalMux I__488 (
            .O(N__4443),
            .I(N__4433));
    LocalMux I__487 (
            .O(N__4438),
            .I(N__4433));
    Odrv4 I__486 (
            .O(N__4433),
            .I(\U712_REG_SM.N_71_i ));
    InMux I__485 (
            .O(N__4430),
            .I(N__4427));
    LocalMux I__484 (
            .O(N__4427),
            .I(N__4423));
    InMux I__483 (
            .O(N__4426),
            .I(N__4420));
    Odrv12 I__482 (
            .O(N__4423),
            .I(REG_CPU_CYCLE));
    LocalMux I__481 (
            .O(N__4420),
            .I(REG_CPU_CYCLE));
    IoInMux I__480 (
            .O(N__4415),
            .I(N__4412));
    LocalMux I__479 (
            .O(N__4412),
            .I(N__4409));
    IoSpan4Mux I__478 (
            .O(N__4409),
            .I(N__4406));
    Span4Mux_s0_h I__477 (
            .O(N__4406),
            .I(N__4403));
    Span4Mux_h I__476 (
            .O(N__4403),
            .I(N__4399));
    InMux I__475 (
            .O(N__4402),
            .I(N__4396));
    Sp12to4 I__474 (
            .O(N__4399),
            .I(N__4393));
    LocalMux I__473 (
            .O(N__4396),
            .I(N__4390));
    Span12Mux_v I__472 (
            .O(N__4393),
            .I(N__4387));
    Span4Mux_v I__471 (
            .O(N__4390),
            .I(N__4384));
    Span12Mux_h I__470 (
            .O(N__4387),
            .I(N__4381));
    Sp12to4 I__469 (
            .O(N__4384),
            .I(N__4378));
    Span12Mux_h I__468 (
            .O(N__4381),
            .I(N__4375));
    Span12Mux_h I__467 (
            .O(N__4378),
            .I(N__4372));
    Odrv12 I__466 (
            .O(N__4375),
            .I(C3_c));
    Odrv12 I__465 (
            .O(N__4372),
            .I(C3_c));
    InMux I__464 (
            .O(N__4367),
            .I(N__4364));
    LocalMux I__463 (
            .O(N__4364),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0 ));
    IoInMux I__462 (
            .O(N__4361),
            .I(N__4358));
    LocalMux I__461 (
            .O(N__4358),
            .I(N__4355));
    Span4Mux_s3_h I__460 (
            .O(N__4355),
            .I(N__4352));
    Span4Mux_h I__459 (
            .O(N__4352),
            .I(N__4349));
    Span4Mux_h I__458 (
            .O(N__4349),
            .I(N__4346));
    Sp12to4 I__457 (
            .O(N__4346),
            .I(N__4342));
    InMux I__456 (
            .O(N__4345),
            .I(N__4339));
    Odrv12 I__455 (
            .O(N__4342),
            .I(TACK_OUTn));
    LocalMux I__454 (
            .O(N__4339),
            .I(TACK_OUTn));
    CascadeMux I__453 (
            .O(N__4334),
            .I(\U712_REG_SM.N_295_cascade_ ));
    InMux I__452 (
            .O(N__4331),
            .I(N__4328));
    LocalMux I__451 (
            .O(N__4328),
            .I(\U712_REG_SM.LDSn_6_iv_i_0_0 ));
    InMux I__450 (
            .O(N__4325),
            .I(N__4318));
    InMux I__449 (
            .O(N__4324),
            .I(N__4318));
    InMux I__448 (
            .O(N__4323),
            .I(N__4315));
    LocalMux I__447 (
            .O(N__4318),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__446 (
            .O(N__4315),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__445 (
            .O(N__4310),
            .I(N__4307));
    LocalMux I__444 (
            .O(N__4307),
            .I(\U712_REG_SM.N_332 ));
    CascadeMux I__443 (
            .O(N__4304),
            .I(N__4301));
    InMux I__442 (
            .O(N__4301),
            .I(N__4298));
    LocalMux I__441 (
            .O(N__4298),
            .I(\U712_REG_SM.UDSn_6_iv_i_0_0 ));
    InMux I__440 (
            .O(N__4295),
            .I(N__4291));
    InMux I__439 (
            .O(N__4294),
            .I(N__4288));
    LocalMux I__438 (
            .O(N__4291),
            .I(\U712_REG_SM.STATE_COUNTER_RNI7KTS1Z0Z_9 ));
    LocalMux I__437 (
            .O(N__4288),
            .I(\U712_REG_SM.STATE_COUNTER_RNI7KTS1Z0Z_9 ));
    IoInMux I__436 (
            .O(N__4283),
            .I(N__4280));
    LocalMux I__435 (
            .O(N__4280),
            .I(N__4277));
    Span4Mux_s2_v I__434 (
            .O(N__4277),
            .I(N__4274));
    Span4Mux_h I__433 (
            .O(N__4274),
            .I(N__4271));
    Sp12to4 I__432 (
            .O(N__4271),
            .I(N__4268));
    Span12Mux_h I__431 (
            .O(N__4268),
            .I(N__4263));
    InMux I__430 (
            .O(N__4267),
            .I(N__4260));
    InMux I__429 (
            .O(N__4266),
            .I(N__4257));
    Odrv12 I__428 (
            .O(N__4263),
            .I(UDSn_c));
    LocalMux I__427 (
            .O(N__4260),
            .I(UDSn_c));
    LocalMux I__426 (
            .O(N__4257),
            .I(UDSn_c));
    InMux I__425 (
            .O(N__4250),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__424 (
            .O(N__4247),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__423 (
            .O(N__4244),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__422 (
            .O(N__4241),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__421 (
            .O(N__4238),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__420 (
            .O(N__4235),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__419 (
            .O(N__4232),
            .I(N__4205));
    ClkMux I__418 (
            .O(N__4231),
            .I(N__4205));
    ClkMux I__417 (
            .O(N__4230),
            .I(N__4205));
    ClkMux I__416 (
            .O(N__4229),
            .I(N__4205));
    ClkMux I__415 (
            .O(N__4228),
            .I(N__4205));
    ClkMux I__414 (
            .O(N__4227),
            .I(N__4205));
    ClkMux I__413 (
            .O(N__4226),
            .I(N__4205));
    ClkMux I__412 (
            .O(N__4225),
            .I(N__4205));
    ClkMux I__411 (
            .O(N__4224),
            .I(N__4205));
    GlobalMux I__410 (
            .O(N__4205),
            .I(N__4202));
    gio2CtrlBuf I__409 (
            .O(N__4202),
            .I(C1_c_g));
    CascadeMux I__408 (
            .O(N__4199),
            .I(\U712_REG_SM.N_330_cascade_ ));
    IoInMux I__407 (
            .O(N__4196),
            .I(N__4193));
    LocalMux I__406 (
            .O(N__4193),
            .I(N__4190));
    Span4Mux_s3_v I__405 (
            .O(N__4190),
            .I(N__4187));
    Span4Mux_h I__404 (
            .O(N__4187),
            .I(N__4184));
    Span4Mux_h I__403 (
            .O(N__4184),
            .I(N__4181));
    Sp12to4 I__402 (
            .O(N__4181),
            .I(N__4178));
    Span12Mux_s11_v I__401 (
            .O(N__4178),
            .I(N__4174));
    InMux I__400 (
            .O(N__4177),
            .I(N__4171));
    Odrv12 I__399 (
            .O(N__4174),
            .I(ASn_c));
    LocalMux I__398 (
            .O(N__4171),
            .I(ASn_c));
    IoInMux I__397 (
            .O(N__4166),
            .I(N__4163));
    LocalMux I__396 (
            .O(N__4163),
            .I(N__4160));
    IoSpan4Mux I__395 (
            .O(N__4160),
            .I(N__4157));
    Span4Mux_s2_v I__394 (
            .O(N__4157),
            .I(N__4154));
    Span4Mux_v I__393 (
            .O(N__4154),
            .I(N__4151));
    Span4Mux_v I__392 (
            .O(N__4151),
            .I(N__4147));
    InMux I__391 (
            .O(N__4150),
            .I(N__4144));
    Odrv4 I__390 (
            .O(N__4147),
            .I(REGENn_c));
    LocalMux I__389 (
            .O(N__4144),
            .I(REGENn_c));
    IoInMux I__388 (
            .O(N__4139),
            .I(N__4136));
    LocalMux I__387 (
            .O(N__4136),
            .I(N__4133));
    Span12Mux_s7_v I__386 (
            .O(N__4133),
            .I(N__4130));
    Odrv12 I__385 (
            .O(N__4130),
            .I(VBENn_c));
    InMux I__384 (
            .O(N__4127),
            .I(N__4124));
    LocalMux I__383 (
            .O(N__4124),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__382 (
            .O(N__4121),
            .I(bfn_8_10_0_));
    InMux I__381 (
            .O(N__4118),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    IoInMux I__380 (
            .O(N__4115),
            .I(N__4112));
    LocalMux I__379 (
            .O(N__4112),
            .I(N__4109));
    Span4Mux_s2_v I__378 (
            .O(N__4109),
            .I(N__4106));
    Span4Mux_v I__377 (
            .O(N__4106),
            .I(N__4103));
    Odrv4 I__376 (
            .O(N__4103),
            .I(CLK80_PLL_i_i));
    IoInMux I__375 (
            .O(N__4100),
            .I(N__4097));
    LocalMux I__374 (
            .O(N__4097),
            .I(N__4094));
    IoSpan4Mux I__373 (
            .O(N__4094),
            .I(N__4091));
    IoSpan4Mux I__372 (
            .O(N__4091),
            .I(N__4088));
    Span4Mux_s2_h I__371 (
            .O(N__4088),
            .I(N__4085));
    Span4Mux_h I__370 (
            .O(N__4085),
            .I(N__4082));
    Odrv4 I__369 (
            .O(N__4082),
            .I(N_882_i));
    CascadeMux I__368 (
            .O(N__4079),
            .I(\U712_REG_SM.N_71_i_cascade_ ));
    InMux I__367 (
            .O(N__4076),
            .I(N__4073));
    LocalMux I__366 (
            .O(N__4073),
            .I(N__4070));
    Span4Mux_v I__365 (
            .O(N__4070),
            .I(N__4067));
    Odrv4 I__364 (
            .O(N__4067),
            .I(TACK_EN_i_ess));
    CascadeMux I__363 (
            .O(N__4064),
            .I(\U712_REG_SM.N_265_cascade_ ));
    IoInMux I__362 (
            .O(N__4061),
            .I(N__4058));
    LocalMux I__361 (
            .O(N__4058),
            .I(N__4055));
    IoSpan4Mux I__360 (
            .O(N__4055),
            .I(N__4052));
    Span4Mux_s2_v I__359 (
            .O(N__4052),
            .I(N__4049));
    Sp12to4 I__358 (
            .O(N__4049),
            .I(N__4046));
    Span12Mux_v I__357 (
            .O(N__4046),
            .I(N__4043));
    Odrv12 I__356 (
            .O(N__4043),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .I(N__4229));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .I(N__4230));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__4231));
    INV \INVU712_CHIP_RAM.DMA_A20C  (
            .O(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .I(N__4225));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .I(N__4227));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .I(N__4224));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__4226));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .I(N__4228));
    INV \INVU712_REG_SM.STATE_COUNTER_2C  (
            .O(\INVU712_REG_SM.STATE_COUNTER_2C_net ),
            .I(N__8862));
    INV \INVU712_REG_SM.STATE_COUNTER_5C  (
            .O(\INVU712_REG_SM.STATE_COUNTER_5C_net ),
            .I(N__8863));
    INV \INVU712_REG_SM.C3_SYNC_0C  (
            .O(\INVU712_REG_SM.C3_SYNC_0C_net ),
            .I(N__8870));
    INV \INVU712_REG_SM.LATCH_REGC  (
            .O(\INVU712_REG_SM.LATCH_REGC_net ),
            .I(N__8865));
    INV \INVU712_REG_SM.UDSnC  (
            .O(\INVU712_REG_SM.UDSnC_net ),
            .I(N__8864));
    INV \INVU712_REG_SM.LDSnC  (
            .O(\INVU712_REG_SM.LDSnC_net ),
            .I(N__8861));
    INV \INVU712_REG_SM.REGENnC  (
            .O(\INVU712_REG_SM.REGENnC_net ),
            .I(N__8871));
    INV \INVU712_REG_SM.STATE_COUNTER_9C  (
            .O(\INVU712_REG_SM.STATE_COUNTER_9C_net ),
            .I(N__8869));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_10_0_));
    ICE_GB CLK40_PLL_derived_clock_RNIIOT (
            .USERSIGNALTOGLOBALBUFFER(N__8335),
            .GLOBALBUFFEROUTPUT(CLK40_PLL_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__8381),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__4696),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4766),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__4415),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_2_1_0.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_2_1_0.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_2_1_0.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_2_1_0 (
            .in0(N__9926),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TACKn_obuft_RNO_LC_5_15_5.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_5_15_5.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_5_15_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 TACKn_obuft_RNO_LC_5_15_5 (
            .in0(N__4076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_882_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_12_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_7_12_5  (
            .in0(N__8284),
            .in1(N__8169),
            .in2(N__8212),
            .in3(N__4323),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNIQANC1_LC_7_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIQANC1_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNIQANC1_LC_7_13_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNIQANC1_LC_7_13_4  (
            .in0(N__4505),
            .in1(N__5114),
            .in2(N__5064),
            .in3(N__4861),
            .lcout(\U712_REG_SM.N_71_i ),
            .ltout(\U712_REG_SM.N_71_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNTER_RNI7KTS1_9_LC_7_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_RNI7KTS1_9_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNTER_RNI7KTS1_9_LC_7_13_5 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_RNI7KTS1_9_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__4487),
            .in2(N__4079),
            .in3(N__6026),
            .lcout(\U712_REG_SM.STATE_COUNTER_RNI7KTS1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_14_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_14_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_14_0 .LUT_INIT=16'b0001111111111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_7_14_0  (
            .in0(N__8216),
            .in1(N__8256),
            .in2(N__8362),
            .in3(N__8498),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9922),
            .ce(N__7370),
            .sr(N__10819));
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_1_LC_7_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_1_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_1_LC_7_14_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI6FIN_1_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__5045),
            .in2(_gnd_net_),
            .in3(N__5108),
            .lcout(\U712_REG_SM.N_265 ),
            .ltout(\U712_REG_SM.N_265_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDSn_RNO_0_LC_7_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_7_14_7 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \U712_REG_SM.UDSn_RNO_0_LC_7_14_7  (
            .in0(N__9261),
            .in1(N__4266),
            .in2(N__4064),
            .in3(N__6022),
            .lcout(\U712_REG_SM.N_332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNTER_RNO_0_0_LC_7_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_RNO_0_0_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNTER_RNO_0_0_LC_7_15_0 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_RNO_0_0_LC_7_15_0  (
            .in0(N__4506),
            .in1(N__5054),
            .in2(N__5125),
            .in3(N__4481),
            .lcout(\U712_REG_SM.N_266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNTER_9_LC_7_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_9_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_9_LC_7_15_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_9_LC_7_15_1  (
            .in0(N__5119),
            .in1(N__5208),
            .in2(_gnd_net_),
            .in3(N__5062),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_9C_net ),
            .ce(),
            .sr(N__10811));
    defparam \U712_REG_SM.UDSn_RNO_1_LC_7_15_2 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_1_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_1_LC_7_15_2 .LUT_INIT=16'b1110111111001100;
    LogicCell40 \U712_REG_SM.UDSn_RNO_1_LC_7_15_2  (
            .in0(N__9260),
            .in1(N__4482),
            .in2(N__5758),
            .in3(N__4864),
            .lcout(\U712_REG_SM.UDSn_6_iv_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNTER_1_LC_7_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_1_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_1_LC_7_15_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_1_LC_7_15_3  (
            .in0(N__4865),
            .in1(N__4507),
            .in2(N__5065),
            .in3(N__5118),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_9C_net ),
            .ce(),
            .sr(N__10811));
    defparam \U712_REG_SM.ASn_LC_7_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_LC_7_15_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_LC_7_15_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \U712_REG_SM.ASn_LC_7_15_6  (
            .in0(N__4447),
            .in1(N__4177),
            .in2(_gnd_net_),
            .in3(N__4483),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_9C_net ),
            .ce(),
            .sr(N__10811));
    defparam \U712_REG_SM.CYCLE_RUN_LC_7_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.CYCLE_RUN_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.CYCLE_RUN_LC_7_15_7 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \U712_REG_SM.CYCLE_RUN_LC_7_15_7  (
            .in0(N__6049),
            .in1(N__4519),
            .in2(_gnd_net_),
            .in3(N__4446),
            .lcout(\U712_REG_SM.CYCLE_RUNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_9C_net ),
            .ce(),
            .sr(N__10811));
    defparam \U712_REG_SM.REGENn_LC_7_16_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_7_16_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_7_16_6 .LUT_INIT=16'b1111110011101110;
    LogicCell40 \U712_REG_SM.REGENn_LC_7_16_6  (
            .in0(N__4150),
            .in1(N__4485),
            .in2(N__5213),
            .in3(N__6047),
            .lcout(REGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.REGENnC_net ),
            .ce(),
            .sr(N__10807));
    defparam \U712_BUFFERS.un1_VBENn_LC_8_9_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_LC_8_9_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_LC_8_9_5  (
            .in0(N__4430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9592),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LLBE_0_i_o3_LC_8_9_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_0_i_o3_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_0_i_o3_LC_8_9_6 .LUT_INIT=16'b1111110010110011;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_0_i_o3_LC_8_9_6  (
            .in0(N__9246),
            .in1(N__9180),
            .in2(N__9094),
            .in3(N__9021),
            .lcout(\U712_BYTE_ENABLE.N_276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_8_10_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_8_10_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_8_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__4127),
            .in2(_gnd_net_),
            .in3(N__4121),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__4232),
            .ce(),
            .sr(N__4814));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_8_10_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_8_10_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_8_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__4562),
            .in2(_gnd_net_),
            .in3(N__4118),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__4232),
            .ce(),
            .sr(N__4814));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_8_10_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_8_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__4589),
            .in2(_gnd_net_),
            .in3(N__4250),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__4232),
            .ce(),
            .sr(N__4814));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_8_10_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_8_10_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_8_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__4601),
            .in2(_gnd_net_),
            .in3(N__4247),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__4232),
            .ce(),
            .sr(N__4814));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_8_10_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_8_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__4576),
            .in2(_gnd_net_),
            .in3(N__4244),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__4232),
            .ce(),
            .sr(N__4814));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_8_10_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_8_10_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_8_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__6190),
            .in2(_gnd_net_),
            .in3(N__4241),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__4232),
            .ce(),
            .sr(N__4814));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_8_10_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_8_10_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_8_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__6205),
            .in2(_gnd_net_),
            .in3(N__4238),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__4232),
            .ce(),
            .sr(N__4814));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_8_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_8_10_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_8_10_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(N__6172),
            .in2(_gnd_net_),
            .in3(N__4235),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4232),
            .ce(),
            .sr(N__4814));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_11_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_8_11_0  (
            .in0(N__7586),
            .in1(N__8582),
            .in2(N__6599),
            .in3(N__7664),
            .lcout(DMA_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9917),
            .ce(N__6524),
            .sr(N__10837));
    defparam \U712_REG_SM.LDSn_RNO_0_LC_8_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_8_12_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_REG_SM.LDSn_RNO_0_LC_8_12_6  (
            .in0(N__8997),
            .in1(N__9245),
            .in2(N__9167),
            .in3(N__4838),
            .lcout(),
            .ltout(\U712_REG_SM.N_330_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_LC_8_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_8_12_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_8_12_7 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \U712_REG_SM.LDSn_LC_8_12_7  (
            .in0(N__4331),
            .in1(N__4888),
            .in2(N__4199),
            .in3(N__4295),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.LDSnC_net ),
            .ce(),
            .sr(N__10829));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_13_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_13_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_8_13_0 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_8_13_0  (
            .in0(N__8170),
            .in1(N__4367),
            .in2(N__7394),
            .in3(N__8248),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9921),
            .ce(),
            .sr(N__10820));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_13_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_13_3 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_13_3 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_8_13_3  (
            .in0(N__4345),
            .in1(N__4324),
            .in2(N__8339),
            .in3(N__8171),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9921),
            .ce(),
            .sr(N__10820));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_13_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_8_13_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_8_13_4  (
            .in0(N__4325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9921),
            .ce(),
            .sr(N__10820));
    defparam \U712_REG_SM.LDSn_RNO_3_LC_8_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_3_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_3_LC_8_13_5 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \U712_REG_SM.LDSn_RNO_3_LC_8_13_5  (
            .in0(N__5759),
            .in1(N__4486),
            .in2(_gnd_net_),
            .in3(N__4863),
            .lcout(),
            .ltout(\U712_REG_SM.N_295_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_RNO_1_LC_8_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_1_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_1_LC_8_13_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_REG_SM.LDSn_RNO_1_LC_8_13_6  (
            .in0(N__6067),
            .in1(N__4887),
            .in2(N__4334),
            .in3(N__6025),
            .lcout(\U712_REG_SM.LDSn_6_iv_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_13_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_8_13_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_8_13_7  (
            .in0(N__8288),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9921),
            .ce(),
            .sr(N__10820));
    defparam \U712_REG_SM.UDSn_LC_8_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_8_14_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_8_14_2 .LUT_INIT=16'b1111110010101010;
    LogicCell40 \U712_REG_SM.UDSn_LC_8_14_2  (
            .in0(N__4267),
            .in1(N__4310),
            .in2(N__4304),
            .in3(N__4294),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.UDSnC_net ),
            .ce(),
            .sr(N__10812));
    defparam \U712_REG_SM.C1_SYNC_1_LC_8_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.C1_SYNC_1_LC_8_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4661),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.UDSnC_net ),
            .ce(),
            .sr(N__10812));
    defparam \U712_REG_SM.C3_SYNC_1_LC_8_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.C3_SYNC_1_LC_8_14_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__4706),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.UDSnC_net ),
            .ce(),
            .sr(N__10812));
    defparam \U712_REG_SM.STATE_COUNTER_RNO_1_0_LC_8_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_RNO_1_0_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNTER_RNO_1_0_LC_8_14_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_RNO_1_0_LC_8_14_5  (
            .in0(N__5253),
            .in1(N__4832),
            .in2(_gnd_net_),
            .in3(N__5202),
            .lcout(),
            .ltout(\U712_REG_SM.STATE_COUNTER_srsts_i_i_i_a3_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNTER_0_LC_8_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_0_LC_8_14_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNTER_0_LC_8_14_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_0_LC_8_14_6  (
            .in0(N__6048),
            .in1(N__4550),
            .in2(N__4544),
            .in3(N__6023),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.UDSnC_net ),
            .ce(),
            .sr(N__10812));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_8_14_7 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_8_14_7  (
            .in0(N__4541),
            .in1(N__4520),
            .in2(N__5653),
            .in3(N__4508),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.UDSnC_net ),
            .ce(),
            .sr(N__10812));
    defparam \U712_REG_SM.LATCH_REG_LC_8_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.LATCH_REG_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.LATCH_REG_LC_8_15_0 .LUT_INIT=16'b1010001110100000;
    LogicCell40 \U712_REG_SM.LATCH_REG_LC_8_15_0  (
            .in0(N__5892),
            .in1(N__4484),
            .in2(N__5237),
            .in3(N__4954),
            .lcout(LATCH_REG),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.LATCH_REGC_net ),
            .ce(),
            .sr(N__10808));
    defparam \U712_REG_SM.REG_WRITE_CYCLE_LC_8_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_WRITE_CYCLE_LC_8_15_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REG_WRITE_CYCLE_LC_8_15_1 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \U712_REG_SM.REG_WRITE_CYCLE_LC_8_15_1  (
            .in0(N__5756),
            .in1(N__4448),
            .in2(_gnd_net_),
            .in3(N__5893),
            .lcout(REG_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.LATCH_REGC_net ),
            .ce(),
            .sr(N__10808));
    defparam \U712_REG_SM.REG_CPU_CYCLE_LC_8_15_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CPU_CYCLE_LC_8_15_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CPU_CYCLE_LC_8_15_2 .LUT_INIT=16'b0100000011100101;
    LogicCell40 \U712_REG_SM.REG_CPU_CYCLE_LC_8_15_2  (
            .in0(N__5170),
            .in1(N__4426),
            .in2(N__5144),
            .in3(N__5206),
            .lcout(REG_CPU_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.LATCH_REGC_net ),
            .ce(),
            .sr(N__10808));
    defparam \U712_REG_SM.REG_CYCLE_LC_8_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_8_15_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_8_15_3 .LUT_INIT=16'b0011001100111010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_8_15_3  (
            .in0(N__7992),
            .in1(N__5132),
            .in2(N__5212),
            .in3(N__5000),
            .lcout(REG_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.LATCH_REGC_net ),
            .ce(),
            .sr(N__10808));
    defparam \U712_REG_SM.STATE_COUNTER_8_LC_8_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_8_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_8_LC_8_15_4 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_8_LC_8_15_4  (
            .in0(N__5255),
            .in1(N__5058),
            .in2(N__5126),
            .in3(N__5207),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.LATCH_REGC_net ),
            .ce(),
            .sr(N__10808));
    defparam \U712_REG_SM.STATE_COUNTER_7_LC_8_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_7_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_7_LC_8_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_7_LC_8_15_5  (
            .in0(N__4982),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.LATCH_REGC_net ),
            .ce(),
            .sr(N__10808));
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_16_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.C3_SYNC_0_LC_8_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4402),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.C3_SYNC_0C_net ),
            .ce(),
            .sr(N__10801));
    defparam \U712_REG_SM.C1_SYNC_0_LC_8_16_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_8_16_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.C1_SYNC_0_LC_8_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4697),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.C3_SYNC_0C_net ),
            .ce(),
            .sr(N__10801));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_8_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_8_2  (
            .in0(N__4652),
            .in1(N__9519),
            .in2(_gnd_net_),
            .in3(N__9326),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_241_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_8_3 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__10024),
            .in2(N__4634),
            .in3(N__9727),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LMBE_0_a3_i_o3_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LMBE_0_a3_i_o3_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LMBE_0_a3_i_o3_LC_9_9_1 .LUT_INIT=16'b1111010001001111;
    LogicCell40 \U712_BYTE_ENABLE.LMBE_0_a3_i_o3_LC_9_9_1  (
            .in0(N__9273),
            .in1(N__9110),
            .in2(N__9185),
            .in3(N__9022),
            .lcout(\U712_BYTE_ENABLE.N_278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_9_9_2 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_9_9_2  (
            .in0(N__7330),
            .in1(N__6949),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0 ),
            .ltout(\U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_47_i_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_47_i_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_47_i_LC_9_9_3 .LUT_INIT=16'b0010001110101111;
    LogicCell40 \U712_BYTE_ENABLE.N_47_i_LC_9_9_3  (
            .in0(N__8111),
            .in1(N__4631),
            .in2(N__4625),
            .in3(N__9591),
            .lcout(N_47_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_9_10_0 .LUT_INIT=16'b0000000001100111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_9_10_0  (
            .in0(N__10295),
            .in1(N__9665),
            .in2(N__10216),
            .in3(N__10248),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_10_3 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_10_3  (
            .in0(N__4600),
            .in1(N__4588),
            .in2(N__4577),
            .in3(N__4561),
            .lcout(\U712_CHIP_RAM.REFRESH5lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_9_10_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_9_10_6  (
            .in0(N__10294),
            .in1(N__9664),
            .in2(N__10215),
            .in3(N__10247),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_9_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_9_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_9_11_0  (
            .in0(N__4805),
            .in1(N__4784),
            .in2(_gnd_net_),
            .in3(N__9709),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_9_11_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_9_11_1  (
            .in0(N__9710),
            .in1(N__9495),
            .in2(N__4769),
            .in3(N__10658),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_11_4 .LUT_INIT=16'b1100000011010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_11_4  (
            .in0(N__5489),
            .in1(N__5535),
            .in2(N__7093),
            .in3(N__8581),
            .lcout(\U712_CHIP_RAM.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_11_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_11_5  (
            .in0(N__6147),
            .in1(N__8459),
            .in2(N__6662),
            .in3(N__7215),
            .lcout(\U712_CHIP_RAM.N_359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_9_11_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__10639),
            .in2(_gnd_net_),
            .in3(N__10873),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_9_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_9_12_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_9_12_1  (
            .in0(N__6655),
            .in1(N__4754),
            .in2(N__11192),
            .in3(N__4712),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_361_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_LC_9_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.BANK0_esr_LC_9_12_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_LC_9_12_2  (
            .in0(N__7232),
            .in1(N__6656),
            .in2(N__4736),
            .in3(N__10628),
            .lcout(BANK0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9918),
            .ce(N__5771),
            .sr(N__10821));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIH3Q74_LC_9_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIH3Q74_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIH3Q74_LC_9_12_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIH3Q74_LC_9_12_4  (
            .in0(N__5620),
            .in1(N__5583),
            .in2(N__6149),
            .in3(N__7214),
            .lcout(\U712_CHIP_RAM.N_452 ),
            .ltout(\U712_CHIP_RAM.N_452_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_12_5 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_9_12_5  (
            .in0(N__6654),
            .in1(N__7727),
            .in2(N__4922),
            .in3(N__7882),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_12_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_LC_9_12_6  (
            .in0(N__10872),
            .in1(_gnd_net_),
            .in2(N__4919),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_13_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_9_13_0  (
            .in0(N__5621),
            .in1(N__5587),
            .in2(N__7246),
            .in3(N__6148),
            .lcout(CPU_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9920),
            .ce(N__4916),
            .sr(N__10813));
    defparam \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_9_13_2 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_9_13_2  (
            .in0(N__7754),
            .in1(N__6548),
            .in2(_gnd_net_),
            .in3(N__7784),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_RNO_2_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_2_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_2_LC_9_13_3 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \U712_REG_SM.LDSn_RNO_2_LC_9_13_3  (
            .in0(N__4886),
            .in1(N__4862),
            .in2(_gnd_net_),
            .in3(N__6011),
            .lcout(\U712_REG_SM.N_309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNTER_RNO_2_0_LC_9_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_RNO_2_0_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNTER_RNO_2_0_LC_9_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_RNO_2_0_LC_9_14_0  (
            .in0(N__4979),
            .in1(N__5165),
            .in2(N__4826),
            .in3(N__5231),
            .lcout(\U712_REG_SM.STATE_COUNTER_srsts_i_i_i_a3_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNTER_5_LC_9_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_5_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_5_LC_9_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_5_LC_9_14_1  (
            .in0(N__5166),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_5C_net ),
            .ce(),
            .sr(N__10809));
    defparam \U712_REG_SM.STATE_COUNTER_4_LC_9_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_4_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_4_LC_9_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_4_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5233),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_5C_net ),
            .ce(),
            .sr(N__10809));
    defparam \U712_REG_SM.STATE_COUNTER_6_LC_9_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_6_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_6_LC_9_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_6_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4825),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_5C_net ),
            .ce(),
            .sr(N__10809));
    defparam \U712_REG_SM.STATE_COUNTER_3_LC_9_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_3_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_3_LC_9_14_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_3_LC_9_14_4  (
            .in0(N__6012),
            .in1(N__5123),
            .in2(N__5066),
            .in3(N__5960),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_5C_net ),
            .ce(),
            .sr(N__10809));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_9_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_9_14_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_9_14_6  (
            .in0(N__4980),
            .in1(N__5254),
            .in2(_gnd_net_),
            .in3(N__5232),
            .lcout(),
            .ltout(\U712_REG_SM.un18_0_i_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_LC_9_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_9_14_7 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_9_14_7  (
            .in0(N__4961),
            .in1(N__4999),
            .in2(N__5216),
            .in3(N__8249),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_5C_net ),
            .ce(),
            .sr(N__10809));
    defparam \U712_REG_SM.STATE_COUNTER_RNIFMLV_8_LC_9_15_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_RNIFMLV_8_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNTER_RNIFMLV_8_LC_9_15_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_RNIFMLV_8_LC_9_15_0  (
            .in0(N__5201),
            .in1(N__5053),
            .in2(_gnd_net_),
            .in3(N__5112),
            .lcout(),
            .ltout(\U712_REG_SM.N_442_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_15_1 .LUT_INIT=16'b0100010001000111;
    LogicCell40 \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_15_1  (
            .in0(N__5891),
            .in1(N__5171),
            .in2(N__5147),
            .in3(N__4998),
            .lcout(\U712_REG_SM.REG_CPU_CYCLE_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_15_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_15_2 .LUT_INIT=16'b0001000100011111;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_9_15_2  (
            .in0(N__5999),
            .in1(N__5889),
            .in2(N__5063),
            .in3(N__5113),
            .lcout(\U712_REG_SM.N_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_9_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_9_15_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_9_15_3  (
            .in0(N__5958),
            .in1(N__5997),
            .in2(N__5124),
            .in3(N__5046),
            .lcout(\U712_REG_SM.N_447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_9_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_9_15_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_9_15_5  (
            .in0(N__5890),
            .in1(N__4981),
            .in2(_gnd_net_),
            .in3(N__5998),
            .lcout(\U712_REG_SM.N_288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.LATCH_CLK_0_i_LC_9_15_7 .C_ON=1'b0;
    defparam \U712_BUFFERS.LATCH_CLK_0_i_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.LATCH_CLK_0_i_LC_9_15_7 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \U712_BUFFERS.LATCH_CLK_0_i_LC_9_15_7  (
            .in0(N__6086),
            .in1(N__4955),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(LATCH_CLK_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_10_7_1  (
            .in0(N__5459),
            .in1(N__5441),
            .in2(_gnd_net_),
            .in3(N__9725),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_2 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_10_7_2  (
            .in0(N__9726),
            .in1(N__9588),
            .in2(N__5420),
            .in3(N__10442),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_10_7_3  (
            .in0(N__5417),
            .in1(N__5399),
            .in2(_gnd_net_),
            .in3(N__9724),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_7_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_7_6  (
            .in0(N__9723),
            .in1(N__5384),
            .in2(_gnd_net_),
            .in3(N__5369),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_10_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_10_8_4 .LUT_INIT=16'b0101111101001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_10_8_4  (
            .in0(N__10036),
            .in1(N__10102),
            .in2(N__9741),
            .in3(N__9589),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_10_8_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(N__5495),
            .in2(N__5354),
            .in3(N__5351),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9901),
            .ce(N__9792),
            .sr(N__10844));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_10_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_10_8_7  (
            .in0(N__6266),
            .in1(N__6299),
            .in2(_gnd_net_),
            .in3(N__5321),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9901),
            .ce(N__9792),
            .sr(N__10844));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_10_9_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_10_9_0  (
            .in0(N__10874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5294),
            .lcout(\U712_CHIP_RAM.un1_CMA28_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_9_3  (
            .in0(N__5288),
            .in1(N__5270),
            .in2(_gnd_net_),
            .in3(N__9702),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_10_9_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__10301),
            .in2(_gnd_net_),
            .in3(N__10211),
            .lcout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux ),
            .ltout(\U712_CHIP_RAM.CMA_5_sn_N_5_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_9_5 .LUT_INIT=16'b0000010011110000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_9_5  (
            .in0(N__9590),
            .in1(N__10103),
            .in2(N__5498),
            .in3(N__9703),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_10_0 .LUT_INIT=16'b0101011111111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_10_0  (
            .in0(N__8497),
            .in1(N__5465),
            .in2(N__7712),
            .in3(N__7660),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_10_1 .LUT_INIT=16'b1010101010100011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_10_1  (
            .in0(N__10302),
            .in1(N__5519),
            .in2(N__6407),
            .in3(N__6369),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9910),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_10_3  (
            .in0(N__5549),
            .in1(N__6143),
            .in2(N__5540),
            .in3(N__6473),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_4 .LUT_INIT=16'b1110111100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_10_4  (
            .in0(N__6398),
            .in1(N__6371),
            .in2(N__5483),
            .in3(N__9714),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9910),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_10_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_10_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_10_5 .LUT_INIT=16'b1111000011010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_10_5  (
            .in0(N__5480),
            .in1(N__6399),
            .in2(N__10224),
            .in3(N__6368),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9910),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_10_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_3_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(N__7445),
            .in2(_gnd_net_),
            .in3(N__7505),
            .lcout(\U712_CHIP_RAM.N_392 ),
            .ltout(\U712_CHIP_RAM.N_392_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_10_7 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_10_7  (
            .in0(N__7579),
            .in1(N__7942),
            .in2(N__5468),
            .in3(N__7876),
            .lcout(\U712_CHIP_RAM.N_449 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_11_0  (
            .in0(N__5536),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5518),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_376_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_1 .LUT_INIT=16'b1110111100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_11_1  (
            .in0(N__6370),
            .in1(N__6400),
            .in2(N__5555),
            .in3(N__10260),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9913),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_0_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_0_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_0_LC_10_11_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_0_LC_10_11_2  (
            .in0(N__7578),
            .in1(N__8579),
            .in2(N__7658),
            .in3(N__6582),
            .lcout(\U712_CHIP_RAM.N_45_i ),
            .ltout(\U712_CHIP_RAM.N_45_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_10_11_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI15FJ4_LC_10_11_3  (
            .in0(N__8455),
            .in1(N__6653),
            .in2(N__5552),
            .in3(N__7867),
            .lcout(\U712_CHIP_RAM.N_324_2 ),
            .ltout(\U712_CHIP_RAM.N_324_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_10_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_10_11_4 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIFMOI5_LC_10_11_4  (
            .in0(N__6126),
            .in1(N__5624),
            .in2(N__5543),
            .in3(N__5588),
            .lcout(\U712_CHIP_RAM.N_324 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFMOI5_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFMOI5_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFMOI5_LC_10_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIFMOI5_LC_10_11_5  (
            .in0(N__8456),
            .in1(N__5507),
            .in2(N__7237),
            .in3(N__7869),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_5_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_4_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_4_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_4_LC_10_11_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNILDP34_4_LC_10_11_6  (
            .in0(N__7868),
            .in1(N__8457),
            .in2(N__7954),
            .in3(N__7119),
            .lcout(\U712_CHIP_RAM.N_450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVC_4_LC_10_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVC_4_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVC_4_LC_10_11_7 .LUT_INIT=16'b1010001010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVC_4_LC_10_11_7  (
            .in0(N__8458),
            .in1(N__7946),
            .in2(N__7236),
            .in3(N__6413),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNIVIFVCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_10_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_10_12_1 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_10_12_1  (
            .in0(N__6649),
            .in1(N__6133),
            .in2(N__5623),
            .in3(N__5582),
            .lcout(\U712_CHIP_RAM.N_252 ),
            .ltout(\U712_CHIP_RAM.N_252_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIURFN4_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIURFN4_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNIURFN4_LC_10_12_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNIURFN4_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5501),
            .in3(N__7213),
            .lcout(\U712_CHIP_RAM.N_365_1 ),
            .ltout(\U712_CHIP_RAM.N_365_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_10_12_3 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_10_12_3  (
            .in0(N__6668),
            .in1(N__7947),
            .in2(N__5777),
            .in3(N__7881),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_10_12_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_10_12_4  (
            .in0(N__10871),
            .in1(_gnd_net_),
            .in2(N__5774),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_12_5 .LUT_INIT=16'b1101111110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_10_12_5  (
            .in0(N__8488),
            .in1(N__6485),
            .in2(N__7342),
            .in3(N__6660),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9915),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_10_12_6.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_10_12_6.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_10_12_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_10_12_6 (
            .in0(N__5942),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_10_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_10_12_7 .LUT_INIT=16'b0101000001011111;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_10_12_7  (
            .in0(N__6256),
            .in1(_gnd_net_),
            .in2(N__6661),
            .in3(N__5757),
            .lcout(\U712_CHIP_RAM.N_294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_LC_10_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_10_13_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_10_13_0 .LUT_INIT=16'b0111111101000000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_10_13_0  (
            .in0(N__6494),
            .in1(N__7711),
            .in2(N__6512),
            .in3(N__5683),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9919),
            .ce(),
            .sr(N__10810));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_13_1 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_13_1  (
            .in0(N__5672),
            .in1(N__9483),
            .in2(N__5657),
            .in3(N__5622),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9919),
            .ce(),
            .sr(N__10810));
    defparam DBR_SYNC_1_LC_10_13_2.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_10_13_2.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_10_13_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_10_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5561),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9919),
            .ce(),
            .sr(N__10810));
    defparam DBR_SYNC_0_LC_10_13_3.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_10_13_3.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_10_13_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 DBR_SYNC_0_LC_10_13_3 (
            .in0(N__5938),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9919),
            .ce(),
            .sr(N__10810));
    defparam \U712_CHIP_RAM.LATCH_RAM_LC_10_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_RAM_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_RAM_LC_10_13_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.LATCH_RAM_LC_10_13_4  (
            .in0(N__6092),
            .in1(N__8578),
            .in2(N__7341),
            .in3(N__6082),
            .lcout(LATCH_RAM),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9919),
            .ce(),
            .sr(N__10810));
    defparam \U712_REG_SM.STATE_COUNTER_2_LC_10_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNTER_2_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNTER_2_LC_10_14_2 .LUT_INIT=16'b1111111110110000;
    LogicCell40 \U712_REG_SM.STATE_COUNTER_2_LC_10_14_2  (
            .in0(N__6071),
            .in1(N__5959),
            .in2(N__6024),
            .in3(N__6056),
            .lcout(\U712_REG_SM.STATE_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_2C_net ),
            .ce(),
            .sr(N__10802));
    defparam \U712_REG_SM.DBR_SYNC_1_LC_10_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_10_14_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_10_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_1_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5906),
            .lcout(\U712_REG_SM.DBR_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_2C_net ),
            .ce(),
            .sr(N__10802));
    defparam \U712_REG_SM.DBR_SYNC_0_LC_10_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_0_LC_10_14_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DBR_SYNC_0_LC_10_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_0_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5931),
            .lcout(\U712_REG_SM.DBR_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_REG_SM.STATE_COUNTER_2C_net ),
            .ce(),
            .sr(N__10802));
    defparam \U712_BUFFERS.DMA_LATCH_EN_1_i_m2_i_m2_LC_10_16_6 .C_ON=1'b0;
    defparam \U712_BUFFERS.DMA_LATCH_EN_1_i_m2_i_m2_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DMA_LATCH_EN_1_i_m2_i_m2_LC_10_16_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \U712_BUFFERS.DMA_LATCH_EN_1_i_m2_i_m2_LC_10_16_6  (
            .in0(N__7094),
            .in1(N__8005),
            .in2(_gnd_net_),
            .in3(N__5900),
            .lcout(N_289),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_7_0  (
            .in0(N__5822),
            .in1(N__5804),
            .in2(_gnd_net_),
            .in3(N__9717),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_7_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_7_1  (
            .in0(N__9718),
            .in1(N__9583),
            .in2(N__5786),
            .in3(N__8690),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_7_4 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_7_4  (
            .in0(N__9582),
            .in1(N__5783),
            .in2(N__9740),
            .in3(N__8678),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_7_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_7_7  (
            .in0(N__9719),
            .in1(N__9584),
            .in2(N__6311),
            .in3(N__10541),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_8_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_8_1  (
            .in0(N__10311),
            .in1(N__9715),
            .in2(_gnd_net_),
            .in3(N__10217),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(\U712_CHIP_RAM.CMA_5_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_8_2 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_8_2  (
            .in0(N__6286),
            .in1(N__9581),
            .in2(N__6302),
            .in3(N__10354),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_8_6 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_8_6  (
            .in0(N__9716),
            .in1(N__6293),
            .in2(N__9598),
            .in3(N__9380),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_8_7 .LUT_INIT=16'b1100101011111111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_11_8_7  (
            .in0(N__10355),
            .in1(N__6287),
            .in2(N__9597),
            .in3(N__8754),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_11_9_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_11_9_0 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_11_9_0  (
            .in0(N__6536),
            .in1(N__6941),
            .in2(N__7247),
            .in3(N__10427),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9902),
            .ce(),
            .sr(N__10830));
    defparam \U712_CHIP_RAM.DBDIR_LC_11_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_11_9_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_11_9_1 .LUT_INIT=16'b0111001011110000;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_11_9_1  (
            .in0(N__7241),
            .in1(N__6260),
            .in2(N__6223),
            .in3(N__6563),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9902),
            .ce(),
            .sr(N__10830));
    defparam \U712_CHIP_RAM.REFRESH_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_11_10_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_11_10_0  (
            .in0(N__6206),
            .in1(N__6191),
            .in2(N__6176),
            .in3(N__6158),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9907),
            .ce(),
            .sr(N__10822));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKCP34_LC_11_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKCP34_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKCP34_LC_11_10_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKCP34_LC_11_10_2  (
            .in0(N__8492),
            .in1(N__7877),
            .in2(_gnd_net_),
            .in3(N__7222),
            .lcout(\U712_CHIP_RAM.N_456 ),
            .ltout(\U712_CHIP_RAM.N_456_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_11_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_11_10_3 .LUT_INIT=16'b0000001100110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__6397),
            .in2(N__6374),
            .in3(N__7952),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8SVVB_3_LC_11_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8SVVB_3_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8SVVB_3_LC_11_10_6 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI8SVVB_3_LC_11_10_6  (
            .in0(N__8493),
            .in1(N__6902),
            .in2(N__7151),
            .in3(N__7124),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_11_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__8580),
            .in2(_gnd_net_),
            .in3(N__6347),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_11_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_11_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_11_1  (
            .in0(N__6337),
            .in1(N__7581),
            .in2(N__8634),
            .in3(N__6344),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__9911),
            .ce(N__8509),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_11_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_11_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_11_2  (
            .in0(N__6341),
            .in1(N__7462),
            .in2(N__8635),
            .in3(N__6326),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(N__9911),
            .ce(N__8509),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_11_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_11_3  (
            .in0(N__8623),
            .in1(N__7515),
            .in2(_gnd_net_),
            .in3(N__6323),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__9911),
            .ce(N__8509),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_11_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_11_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_11_4  (
            .in0(N__8629),
            .in1(N__7953),
            .in2(_gnd_net_),
            .in3(N__6320),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__9911),
            .ce(N__8509),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_11_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_11_11_5  (
            .in0(N__8624),
            .in1(N__6440),
            .in2(_gnd_net_),
            .in3(N__6317),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__9911),
            .ce(N__8509),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_11_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_11_6  (
            .in0(N__8630),
            .in1(N__6452),
            .in2(_gnd_net_),
            .in3(N__6314),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__9911),
            .ce(N__8509),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_11_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_11_7  (
            .in0(N__6464),
            .in1(N__8628),
            .in2(_gnd_net_),
            .in3(N__6476),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9911),
            .ce(N__8509),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_0_0_LC_11_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_0_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_0_0_LC_11_12_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_0_0_LC_11_12_0  (
            .in0(N__7641),
            .in1(N__7574),
            .in2(_gnd_net_),
            .in3(N__8557),
            .lcout(\U712_CHIP_RAM.N_388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_12_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_12_1  (
            .in0(N__6422),
            .in1(N__8479),
            .in2(N__7886),
            .in3(N__7948),
            .lcout(\U712_CHIP_RAM.N_363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_12_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_11_12_2  (
            .in0(N__7856),
            .in1(N__7514),
            .in2(N__7955),
            .in3(N__7123),
            .lcout(\U712_CHIP_RAM.N_351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_11_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_11_12_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_11_12_3  (
            .in0(N__6463),
            .in1(N__6451),
            .in2(_gnd_net_),
            .in3(N__6439),
            .lcout(\U712_CHIP_RAM.N_384 ),
            .ltout(\U712_CHIP_RAM.N_384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3PIP2_0_LC_11_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3PIP2_0_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3PIP2_0_LC_11_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3PIP2_0_LC_11_12_4  (
            .in0(N__7455),
            .in1(N__7575),
            .in2(N__6428),
            .in3(N__8558),
            .lcout(\U712_CHIP_RAM.N_400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_0_LC_11_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_0_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_0_LC_11_12_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_0_LC_11_12_5  (
            .in0(N__7573),
            .in1(N__8562),
            .in2(_gnd_net_),
            .in3(N__7642),
            .lcout(\U712_CHIP_RAM.N_448 ),
            .ltout(\U712_CHIP_RAM.N_448_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6B326_2_LC_11_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6B326_2_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6B326_2_LC_11_12_6 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6B326_2_LC_11_12_6  (
            .in0(N__7456),
            .in1(N__7651),
            .in2(N__6425),
            .in3(N__7400),
            .lcout(\U712_CHIP_RAM.N_255 ),
            .ltout(\U712_CHIP_RAM.N_255_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5T4O8_LC_11_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5T4O8_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5T4O8_LC_11_12_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI5T4O8_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(N__7855),
            .in2(N__6416),
            .in3(N__7271),
            .lcout(\U712_CHIP_RAM.N_269 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_11_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_11_13_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_11_13_0  (
            .in0(N__7273),
            .in1(N__7776),
            .in2(N__6611),
            .in3(N__7746),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_11_13_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_11_13_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNI892R_LC_11_13_1  (
            .in0(N__7857),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6648),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI4LVP1_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI4LVP1_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI4LVP1_LC_11_13_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI4LVP1_LC_11_13_2  (
            .in0(N__7331),
            .in1(N__7684),
            .in2(_gnd_net_),
            .in3(N__7463),
            .lcout(\U712_CHIP_RAM.N_444 ),
            .ltout(\U712_CHIP_RAM.N_444_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFGIT5_LC_11_13_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFGIT5_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFGIT5_LC_11_13_3 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNIFGIT5_LC_11_13_3  (
            .in0(N__6595),
            .in1(N__7272),
            .in2(N__6566),
            .in3(N__6559),
            .lcout(\U712_CHIP_RAM.N_334 ),
            .ltout(\U712_CHIP_RAM.N_334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI7SS3A_LC_11_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI7SS3A_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNI7SS3A_LC_11_13_4 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNI7SS3A_LC_11_13_4  (
            .in0(N__7079),
            .in1(N__7464),
            .in2(N__6539),
            .in3(N__7777),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_13_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_13_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6527),
            .in3(N__10870),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNISH5V3_LC_11_13_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNISH5V3_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNISH5V3_LC_11_13_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNISH5V3_LC_11_13_6  (
            .in0(N__9566),
            .in1(N__7747),
            .in2(N__6511),
            .in3(N__7150),
            .lcout(\U712_CHIP_RAM.N_323 ),
            .ltout(\U712_CHIP_RAM.N_323_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_13_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_13_7 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_11_13_7  (
            .in0(N__7519),
            .in1(N__9567),
            .in2(N__6488),
            .in3(N__7080),
            .lcout(\U712_CHIP_RAM.N_117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_15_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_15_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__8129),
            .in2(_gnd_net_),
            .in3(N__8122),
            .lcout(\U712_CHIP_RAM.un3_DMA_CYCLE_START ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_12_7_0 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_12_7_0  (
            .in0(N__10054),
            .in1(N__9988),
            .in2(N__10151),
            .in3(N__6863),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9896),
            .ce(N__9839),
            .sr(N__10836));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_12_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_12_7_1 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_12_7_1  (
            .in0(N__10053),
            .in1(N__8702),
            .in2(N__9996),
            .in3(N__6836),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9896),
            .ce(N__9839),
            .sr(N__10836));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_12_7_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_12_7_3  (
            .in0(N__10052),
            .in1(N__8696),
            .in2(N__9995),
            .in3(N__6809),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9896),
            .ce(N__9839),
            .sr(N__10836));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_12_7_4 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_12_7_4  (
            .in0(N__9431),
            .in1(N__9987),
            .in2(N__10058),
            .in3(N__6782),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9896),
            .ce(N__9839),
            .sr(N__10836));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_12_7_5 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_12_7_5  (
            .in0(N__6749),
            .in1(N__9593),
            .in2(N__8764),
            .in3(N__10070),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9896),
            .ce(N__9839),
            .sr(N__10836));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_12_8_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_12_8_2  (
            .in0(N__10051),
            .in1(N__8666),
            .in2(N__9997),
            .in3(N__6719),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9899),
            .ce(N__9829),
            .sr(N__10828));
    defparam \U712_BYTE_ENABLE.N_46_i_LC_12_9_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_46_i_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_46_i_LC_12_9_0 .LUT_INIT=16'b0000110111011101;
    LogicCell40 \U712_BYTE_ENABLE.N_46_i_LC_12_9_0  (
            .in0(N__6919),
            .in1(N__8107),
            .in2(N__6968),
            .in3(N__9575),
            .lcout(N_46_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UUBE_0_a2_0_a2_LC_12_9_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_0_a2_0_a2_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_0_a2_0_a2_LC_12_9_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_0_a2_0_a2_LC_12_9_1  (
            .in0(N__9272),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9093),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.UUBE_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_48_i_LC_12_9_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_48_i_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_48_i_LC_12_9_2 .LUT_INIT=16'b0000110111011101;
    LogicCell40 \U712_BYTE_ENABLE.N_48_i_LC_12_9_2  (
            .in0(N__6920),
            .in1(N__8056),
            .in2(N__7034),
            .in3(N__9576),
            .lcout(N_48_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_49_i_LC_12_9_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_49_i_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_49_i_LC_12_9_3 .LUT_INIT=16'b0100110001011111;
    LogicCell40 \U712_BYTE_ENABLE.N_49_i_LC_12_9_3  (
            .in0(N__9577),
            .in1(N__8057),
            .in2(N__7007),
            .in3(N__6995),
            .lcout(N_49_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_0_i_o3_LC_12_9_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_0_i_o3_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_0_i_o3_LC_12_9_4 .LUT_INIT=16'b1101011111010011;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_0_i_o3_LC_12_9_4  (
            .in0(N__9092),
            .in1(N__9184),
            .in2(N__9026),
            .in3(N__9271),
            .lcout(\U712_BYTE_ENABLE.N_277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_LC_12_9_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_LC_12_9_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_LC_12_9_7  (
            .in0(N__6942),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7343),
            .lcout(\U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHC4P1_2_LC_12_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHC4P1_2_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHC4P1_2_LC_12_10_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIHC4P1_2_LC_12_10_0  (
            .in0(N__8460),
            .in1(N__7941),
            .in2(N__7466),
            .in3(N__7839),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_10_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_12_10_2  (
            .in0(N__9731),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9520),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPORK3_1_LC_12_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPORK3_1_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIPORK3_1_LC_12_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIPORK3_1_LC_12_10_6  (
            .in0(N__8461),
            .in1(N__7580),
            .in2(N__7707),
            .in3(N__7659),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_325_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE6LO7_1_LC_12_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE6LO7_1_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIE6LO7_1_LC_12_10_7 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIE6LO7_1_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__6911),
            .in2(N__6905),
            .in3(N__7277),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_12_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_LC_12_11_1 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_LC_12_11_1  (
            .in0(N__7066),
            .in1(N__7854),
            .in2(N__6893),
            .in3(N__7355),
            .lcout(WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9903),
            .ce(),
            .sr(N__10806));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8ALV_LC_12_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8ALV_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8ALV_LC_12_11_2 .LUT_INIT=16'b1000100011111111;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8ALV_LC_12_11_2  (
            .in0(N__7323),
            .in1(N__7460),
            .in2(_gnd_net_),
            .in3(N__7507),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_305_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_4_LC_12_11_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_4_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_4_LC_12_11_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_4_LC_12_11_3  (
            .in0(N__7940),
            .in1(N__7852),
            .in2(N__7280),
            .in3(N__7270),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIUHSBF_LC_12_11_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIUHSBF_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIUHSBF_LC_12_11_4 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIUHSBF_LC_12_11_4  (
            .in0(N__7245),
            .in1(N__8432),
            .in2(N__7160),
            .in3(N__7157),
            .lcout(\U712_CHIP_RAM.N_202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNITVQE7_LC_12_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNITVQE7_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNITVQE7_LC_12_11_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNITVQE7_LC_12_11_5  (
            .in0(N__7143),
            .in1(N__7775),
            .in2(N__7078),
            .in3(N__7117),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_180_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_3_LC_12_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_3_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_3_LC_12_11_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_3_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__7939),
            .in2(_gnd_net_),
            .in3(N__7506),
            .lcout(\U712_CHIP_RAM.N_407 ),
            .ltout(\U712_CHIP_RAM.N_407_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_11_7 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__7853),
            .in2(N__7127),
            .in3(N__7118),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9903),
            .ce(),
            .sr(N__10806));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_12_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_12_12_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__7062),
            .in2(_gnd_net_),
            .in3(N__7454),
            .lcout(\U712_CHIP_RAM.N_257 ),
            .ltout(\U712_CHIP_RAM.N_257_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_12_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_12_12_1 .LUT_INIT=16'b0001111100010001;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_12_12_1  (
            .in0(N__8560),
            .in1(N__7461),
            .in2(N__7037),
            .in3(N__7577),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS3891_3_LC_12_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS3891_3_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS3891_3_LC_12_12_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIS3891_3_LC_12_12_3  (
            .in0(N__7938),
            .in1(N__7504),
            .in2(_gnd_net_),
            .in3(N__7828),
            .lcout(\U712_CHIP_RAM.N_396 ),
            .ltout(\U712_CHIP_RAM.N_396_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_12_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_12_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_0_LC_12_12_4  (
            .in0(N__7576),
            .in1(N__8559),
            .in2(N__7787),
            .in3(N__7643),
            .lcout(\U712_CHIP_RAM.N_436 ),
            .ltout(\U712_CHIP_RAM.N_436_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_12_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_12_12_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7757),
            .in3(N__7745),
            .lcout(\U712_CHIP_RAM.N_357 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_12_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_12_12_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_12_12_6  (
            .in0(N__7718),
            .in1(N__7703),
            .in2(_gnd_net_),
            .in3(N__7644),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_12_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_12_12_7 .LUT_INIT=16'b1111111000000010;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_12_12_7  (
            .in0(N__8204),
            .in1(N__7601),
            .in2(N__7595),
            .in3(N__7592),
            .lcout(CPU_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9909),
            .ce(),
            .sr(N__10800));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_12_13_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_12_13_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_12_13_0  (
            .in0(N__7585),
            .in1(N__8561),
            .in2(N__7523),
            .in3(N__7465),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_0_a2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_12_13_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_12_13_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_12_13_1  (
            .in0(N__8463),
            .in1(N__8358),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_274_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_13_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_13_2 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_12_13_2  (
            .in0(N__8194),
            .in1(N__7393),
            .in2(N__7376),
            .in3(N__8257),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_274_i_0_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_12_13_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_12_13_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7373),
            .in3(N__8374),
            .lcout(\U712_CYCLE_TERM.N_274_i_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_13_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_13_4 .LUT_INIT=16'b1111110010101100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_13_4  (
            .in0(N__8660),
            .in1(N__8648),
            .in2(N__8639),
            .in3(N__8594),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9912),
            .ce(N__8513),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_13_5.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_13_5.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_13_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_13_5 (
            .in0(N__8462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_13_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_13_6 .LUT_INIT=16'b0000010100001111;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_12_13_6  (
            .in0(N__8147),
            .in1(_gnd_net_),
            .in2(N__8363),
            .in3(N__8878),
            .lcout(\U712_CYCLE_TERM.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_12_14_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_12_14_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_12_14_1  (
            .in0(N__8328),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8153),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9914),
            .ce(),
            .sr(N__10799));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_14_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_12_14_5 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_12_14_5  (
            .in0(N__8264),
            .in1(N__8154),
            .in2(N__8258),
            .in3(N__8211),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9914),
            .ce(),
            .sr(N__10799));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_12_15_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_12_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8123),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9916),
            .ce(),
            .sr(N__10798));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_12_15_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_12_15_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_12_15_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__8094),
            .in2(_gnd_net_),
            .in3(N__8049),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9916),
            .ce(),
            .sr(N__10798));
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_12_16_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_12_16_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_0_a2_0_a3_LC_12_16_1  (
            .in0(N__8093),
            .in1(N__8039),
            .in2(_gnd_net_),
            .in3(N__8006),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLK40_PLL_derived_clock_RNIIOT_0_LC_12_20_2.C_ON=1'b0;
    defparam CLK40_PLL_derived_clock_RNIIOT_0_LC_12_20_2.SEQ_MODE=4'b0000;
    defparam CLK40_PLL_derived_clock_RNIIOT_0_LC_12_20_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40_PLL_derived_clock_RNIIOT_0_LC_12_20_2 (
            .in0(N__8879),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_iso_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_12_20_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_12_20_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_i_LC_12_20_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_i_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(N__9274),
            .in2(_gnd_net_),
            .in3(N__9084),
            .lcout(U712_BYTE_ENABLE_UUBE_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_6_5 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_13_6_5  (
            .in0(N__8765),
            .in1(N__8738),
            .in2(N__9602),
            .in3(N__10613),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9897),
            .ce(N__9833),
            .sr(N__10848));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_7_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_7_2  (
            .in0(N__10136),
            .in1(_gnd_net_),
            .in2(N__11188),
            .in3(N__9422),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10943),
            .ce(N__10914),
            .sr(N__10845));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_7  (
            .in0(N__9368),
            .in1(N__9421),
            .in2(_gnd_net_),
            .in3(N__11177),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10943),
            .ce(N__10914),
            .sr(N__10845));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_8_0  (
            .in0(N__11183),
            .in1(N__9414),
            .in2(_gnd_net_),
            .in3(N__10134),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__10912),
            .sr(N__10838));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_1  (
            .in0(N__10135),
            .in1(_gnd_net_),
            .in2(N__10697),
            .in3(N__11184),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net ),
            .ce(N__10912),
            .sr(N__10838));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_9_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_13_9_4  (
            .in0(N__9367),
            .in1(N__10411),
            .in2(_gnd_net_),
            .in3(N__11181),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10940),
            .ce(N__10911),
            .sr(N__10831));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_9_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_9_7  (
            .in0(N__11182),
            .in1(N__10693),
            .in2(_gnd_net_),
            .in3(N__10529),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10940),
            .ce(N__10911),
            .sr(N__10831));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_10_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_13_10_2  (
            .in0(N__11113),
            .in1(N__9360),
            .in2(_gnd_net_),
            .in3(N__9413),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__10909),
            .sr(N__10823));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_11_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_11_5  (
            .in0(N__11163),
            .in1(N__10410),
            .in2(_gnd_net_),
            .in3(N__9359),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net ),
            .ce(N__10907),
            .sr(N__10814));
    defparam \U712_BYTE_ENABLE.N_276_i_LC_13_20_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_276_i_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_276_i_LC_13_20_1 .LUT_INIT=16'b0000001101001100;
    LogicCell40 \U712_BYTE_ENABLE.N_276_i_LC_13_20_1  (
            .in0(N__9282),
            .in1(N__9177),
            .in2(N__9108),
            .in3(N__9006),
            .lcout(N_276_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_278_i_LC_13_20_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_278_i_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_278_i_LC_13_20_2 .LUT_INIT=16'b0100100001011010;
    LogicCell40 \U712_BYTE_ENABLE.N_278_i_LC_13_20_2  (
            .in0(N__9179),
            .in1(N__9284),
            .in2(N__9020),
            .in3(N__9104),
            .lcout(N_278_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_277_i_LC_13_20_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_277_i_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_277_i_LC_13_20_5 .LUT_INIT=16'b0011000011000100;
    LogicCell40 \U712_BYTE_ENABLE.N_277_i_LC_13_20_5  (
            .in0(N__9283),
            .in1(N__9178),
            .in2(N__9109),
            .in3(N__9007),
            .lcout(N_277_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CRCSn_LC_14_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_14_4_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_14_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_14_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10267),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9895),
            .ce(),
            .sr(N__10854));
    defparam \U712_CHIP_RAM.RASn_LC_14_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_14_4_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_14_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_14_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10322),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9895),
            .ce(),
            .sr(N__10854));
    defparam \U712_CHIP_RAM.CASn_LC_14_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_14_5_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_14_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_14_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9743),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9898),
            .ce(),
            .sr(N__10853));
    defparam \U712_CHIP_RAM.WEn_LC_14_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_14_5_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_14_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_14_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10231),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9898),
            .ce(),
            .sr(N__10853));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_14_7_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_14_7_1  (
            .in0(N__10321),
            .in1(N__9742),
            .in2(N__10271),
            .in3(N__10232),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9900),
            .ce(N__9837),
            .sr(N__10849));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_1  (
            .in0(N__10527),
            .in1(N__10477),
            .in2(_gnd_net_),
            .in3(N__11155),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10941),
            .ce(N__10915),
            .sr(N__10846));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_8_3  (
            .in0(N__10125),
            .in1(N__10686),
            .in2(_gnd_net_),
            .in3(N__11154),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10941),
            .ce(N__10915),
            .sr(N__10846));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_7  (
            .in0(N__10082),
            .in1(N__10600),
            .in2(_gnd_net_),
            .in3(N__11156),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10941),
            .ce(N__10915),
            .sr(N__10846));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_14_9_5 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_14_9_5  (
            .in0(N__10050),
            .in1(N__10952),
            .in2(N__9998),
            .in3(N__9437),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9908),
            .ce(N__9838),
            .sr(N__10839));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_14_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_14_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_14_10_0  (
            .in0(N__9776),
            .in1(N__9764),
            .in2(_gnd_net_),
            .in3(N__9735),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_10_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_10_1  (
            .in0(N__9736),
            .in1(N__9568),
            .in2(N__9440),
            .in3(N__10418),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_14_11_0  (
            .in0(N__10685),
            .in1(N__10528),
            .in2(_gnd_net_),
            .in3(N__11099),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net ),
            .ce(N__10908),
            .sr(N__10824));
    defparam \U712_CHIP_RAM.DMA_A20_LC_14_12_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A20_LC_14_12_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A20_LC_14_12_2 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_A20_LC_14_12_2  (
            .in0(N__11083),
            .in1(N__10646),
            .in2(N__10586),
            .in3(N__10627),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A20C_net ),
            .ce(),
            .sr(N__10815));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_15_7_3  (
            .in0(N__10601),
            .in1(N__10478),
            .in2(_gnd_net_),
            .in3(N__11112),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10942),
            .ce(N__10919),
            .sr(N__10852));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_8_7  (
            .in0(N__10599),
            .in1(N__10476),
            .in2(_gnd_net_),
            .in3(N__11153),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__10917),
            .sr(N__10850));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_9_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_9_1  (
            .in0(N__11152),
            .in1(N__10526),
            .in2(_gnd_net_),
            .in3(N__10459),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__10916),
            .sr(N__10847));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_15_9_5  (
            .in0(N__10996),
            .in1(N__11151),
            .in2(_gnd_net_),
            .in3(N__11021),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net ),
            .ce(N__10916),
            .sr(N__10847));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_10_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_15_10_1  (
            .in0(N__10412),
            .in1(N__10997),
            .in2(_gnd_net_),
            .in3(N__11150),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net ),
            .ce(N__10913),
            .sr(N__10840));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_11_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_11_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_11_1  (
            .in0(N__10991),
            .in1(N__10400),
            .in2(_gnd_net_),
            .in3(N__11087),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10939),
            .ce(N__10910),
            .sr(N__10832));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_9_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_16_9_1  (
            .in0(N__11157),
            .in1(N__11020),
            .in2(_gnd_net_),
            .in3(N__10995),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10938),
            .ce(N__10918),
            .sr(N__10851));
endmodule // U712_TOP

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Feb 4 2025 21:50:11

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U111_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U111_TOP
entity U111_TOP is
port (
    D_LL_AMIGA : inout std_logic_vector(7 downto 0);
    D_LM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UU_AMIGA : inout std_logic_vector(7 downto 0);
    D_UM_AMIGA : inout std_logic_vector(7 downto 0);
    D_LL_040 : inout std_logic_vector(7 downto 0);
    D_UU_040 : inout std_logic_vector(7 downto 0);
    D_UM_040 : inout std_logic_vector(7 downto 0);
    D_LM_040 : inout std_logic_vector(7 downto 0);
    A_AMIGA : out std_logic_vector(1 downto 0);
    A_040 : in std_logic_vector(1 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    TSn : out std_logic;
    RESETn : in std_logic;
    CLKRAMA : out std_logic;
    PORTSIZE : in std_logic;
    TEA_CPUn : out std_logic;
    CLK40B : out std_logic;
    TBI_CPUn : out std_logic;
    TAn : out std_logic;
    CPUBGn : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CLK80_CPU : out std_logic;
    BUFDIR : out std_logic;
    TCI_CPUn : out std_logic;
    TS_CPUn : in std_logic;
    CLKRAMB : out std_logic;
    CLK40A : out std_logic;
    DMAn : out std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    TACKn : in std_logic;
    BGn : in std_logic);
end U111_TOP;

-- Architecture of U111_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U111_TOP is

signal \N__8315\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7884\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6431\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5262\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5010\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4896\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4560\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4254\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4005\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3993\ : std_logic;
signal \N__3990\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3846\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3750\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3726\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3660\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3456\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3291\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3279\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3264\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3246\ : std_logic;
signal \N__3243\ : std_logic;
signal \N__3240\ : std_logic;
signal \N__3237\ : std_logic;
signal \N__3234\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3204\ : std_logic;
signal \N__3201\ : std_logic;
signal \N__3198\ : std_logic;
signal \N__3195\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3069\ : std_logic;
signal \N__3066\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3024\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3018\ : std_logic;
signal \N__3015\ : std_logic;
signal \N__3012\ : std_logic;
signal \N__3009\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2982\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2934\ : std_logic;
signal \N__2931\ : std_logic;
signal \N__2928\ : std_logic;
signal \N__2925\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2919\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2913\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2874\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2844\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2835\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2817\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2748\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2655\ : std_logic;
signal \N__2652\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2637\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2625\ : std_logic;
signal \N__2622\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2586\ : std_logic;
signal \N__2583\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2577\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2571\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2565\ : std_logic;
signal \N__2562\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2527\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2461\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2359\ : std_logic;
signal \N__2356\ : std_logic;
signal \N__2353\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2317\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2232\ : std_logic;
signal \N__2229\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \A_040_c_0\ : std_logic;
signal \A_AMIGA_c_0\ : std_logic;
signal \A_040_c_1\ : std_logic;
signal \D_LL_AMIGA_in_2\ : std_logic;
signal \un1_D_LL_AMIGA_2\ : std_logic;
signal \RnW_c_i_0\ : std_logic;
signal \D_UM_040_in_0\ : std_logic;
signal \D_LL_040_in_0\ : std_logic;
signal \un1_D_UM_040_0\ : std_logic;
signal \D_LM_AMIGA_in_1\ : std_logic;
signal \un1_D_LM_AMIGA_1\ : std_logic;
signal \D_UM_040_in_6\ : std_logic;
signal \D_LL_040_in_6\ : std_logic;
signal \un1_D_UM_040_6\ : std_logic;
signal \D_UM_040_in_4\ : std_logic;
signal \D_LL_040_in_4\ : std_logic;
signal \un1_D_UM_040_4\ : std_logic;
signal \D_UU_040_in_3\ : std_logic;
signal \D_LM_040_in_3\ : std_logic;
signal \un1_D_UU_040_3\ : std_logic;
signal \D_LM_040_in_6\ : std_logic;
signal \D_UU_040_in_6\ : std_logic;
signal \un1_D_UU_040_6\ : std_logic;
signal \D_LL_AMIGA_in_7\ : std_logic;
signal \un1_D_LL_AMIGA_7\ : std_logic;
signal \D_LL_040_in_1\ : std_logic;
signal \D_UM_040_in_1\ : std_logic;
signal \un1_D_UM_040_1\ : std_logic;
signal \D_UU_040_in_7\ : std_logic;
signal \D_LM_040_in_7\ : std_logic;
signal \un1_D_UU_040_7\ : std_logic;
signal \D_LL_AMIGA_in_4\ : std_logic;
signal \un1_D_LL_AMIGA_4\ : std_logic;
signal \D_UM_040_in_2\ : std_logic;
signal \D_LL_040_in_2\ : std_logic;
signal \un1_D_UM_040_2\ : std_logic;
signal \D_LM_AMIGA_in_3\ : std_logic;
signal \un1_D_LM_AMIGA_3\ : std_logic;
signal \D_LM_AMIGA_in_5\ : std_logic;
signal \un1_D_LM_AMIGA_5\ : std_logic;
signal \D_UU_040_in_4\ : std_logic;
signal \D_LM_040_in_4\ : std_logic;
signal \un1_D_UU_040_4\ : std_logic;
signal \D_LL_AMIGA_in_0\ : std_logic;
signal \un1_D_LL_AMIGA_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \INVU111_CYCLE_SM.TSnC_net\ : std_logic;
signal \D_LM_AMIGA_in_2\ : std_logic;
signal \un1_D_LM_AMIGA_2\ : std_logic;
signal \D_LM_AMIGA_in_6\ : std_logic;
signal \un1_D_LM_AMIGA_6\ : std_logic;
signal \D_UU_040_in_1\ : std_logic;
signal \D_LM_040_in_1\ : std_logic;
signal \un1_D_UU_040_1\ : std_logic;
signal \D_UU_040_in_2\ : std_logic;
signal \D_LM_040_in_2\ : std_logic;
signal \un1_D_UU_040_2\ : std_logic;
signal \D_LL_AMIGA_in_6\ : std_logic;
signal \un1_D_LL_AMIGA_6\ : std_logic;
signal \D_LL_040_in_3\ : std_logic;
signal \D_UM_040_in_3\ : std_logic;
signal \un1_D_UM_040_3\ : std_logic;
signal \D_LL_AMIGA_in_3\ : std_logic;
signal \un1_D_LL_AMIGA_3\ : std_logic;
signal \D_LL_AMIGA_in_1\ : std_logic;
signal \un1_D_LL_AMIGA_1\ : std_logic;
signal \D_LL_AMIGA_in_5\ : std_logic;
signal \un1_D_LL_AMIGA_5\ : std_logic;
signal \D_LM_AMIGA_in_0\ : std_logic;
signal \un1_D_LM_AMIGA_0\ : std_logic;
signal \un1_D_UM_AMIGA_0\ : std_logic;
signal \INVU111_CYCLE_SM.TA_ENC_net\ : std_logic;
signal \U111_CYCLE_SM.RESETn_c_i\ : std_logic;
signal \INVU111_CYCLE_SM.A_OUTC_net\ : std_logic;
signal \U111_CYCLE_SM.A_OUTZ0\ : std_logic;
signal \U111_CYCLE_SM.A_OUT_0\ : std_logic;
signal \D_UM_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\ : std_logic;
signal \D_LM_AMIGA_in_4\ : std_logic;
signal \un1_D_LM_AMIGA_4\ : std_logic;
signal \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \D_LM_AMIGA_in_7\ : std_logic;
signal \un1_D_LM_AMIGA_7\ : std_logic;
signal \D_UM_040_in_7\ : std_logic;
signal \D_LL_040_in_7\ : std_logic;
signal \un1_D_UM_040_7\ : std_logic;
signal \D_UU_040_in_0\ : std_logic;
signal \D_LM_040_in_0\ : std_logic;
signal \un1_D_UU_040_0\ : std_logic;
signal \D_LL_040_in_5\ : std_logic;
signal \D_UM_040_in_5\ : std_logic;
signal \un1_D_UM_040_5\ : std_logic;
signal \D_UU_040_in_5\ : std_logic;
signal \D_LM_040_in_5\ : std_logic;
signal \A_AMIGA_c_1\ : std_logic;
signal \un1_D_UU_040_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\ : std_logic;
signal \D_UU_AMIGA_in_6\ : std_logic;
signal \un1_D_UU_AMIGA_6\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\ : std_logic;
signal \D_UU_AMIGA_in_2\ : std_logic;
signal \un1_D_UU_AMIGA_2\ : std_logic;
signal \GB_BUFFER_CLK40_THRU_CO\ : std_logic;
signal \U111_CYCLE_SM.TA_ENZ0\ : std_logic;
signal \U111_CYCLE_SM_TAn_0_i\ : std_logic;
signal \U111_CYCLE_SM.un1_LW_TRANS_1_0\ : std_logic;
signal \PORTSIZE_c\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.un3_LW_CYCLE_START_cascade_\ : std_logic;
signal \INVU111_CYCLE_SM.TS_ENC_net\ : std_logic;
signal \TS_CPUn_c\ : std_logic;
signal \U111_CYCLE_SM.TS_EN_5\ : std_logic;
signal \U111_CYCLE_SM.N_69_0\ : std_logic;
signal \CLK40\ : std_logic;
signal \U111_CYCLE_SM.N_91_cascade_\ : std_logic;
signal \INVU111_CYCLE_SM.CYCLE_STATE_0C_net\ : std_logic;
signal \D_UM_AMIGA_in_6\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\ : std_logic;
signal \un1_D_UM_AMIGA_6\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLE_STARTZ0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0_cascade_\ : std_logic;
signal \INVU111_CYCLE_SM.LW_CYCLEC_net\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\ : std_logic;
signal \TACKn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLE_0\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\ : std_logic;
signal \CLK80\ : std_logic;
signal \GB_BUFFER_CLK80_THRU_CO\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\ : std_logic;
signal \D_UM_AMIGA_in_1\ : std_logic;
signal \un1_D_UM_AMIGA_1\ : std_logic;
signal \D_UM_AMIGA_in_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\ : std_logic;
signal \un1_D_UM_AMIGA_3\ : std_logic;
signal \D_UM_AMIGA_in_7\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\ : std_logic;
signal \un1_D_UM_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\ : std_logic;
signal \D_UM_AMIGA_in_4\ : std_logic;
signal \un1_D_UM_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\ : std_logic;
signal \D_UU_AMIGA_in_5\ : std_logic;
signal \un1_D_UU_AMIGA_5\ : std_logic;
signal \D_UU_AMIGA_in_3\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\ : std_logic;
signal \un1_D_UU_AMIGA_3\ : std_logic;
signal \un1_D_UM_AMIGA_2\ : std_logic;
signal \D_UM_AMIGA_in_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_2C_net\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\ : std_logic;
signal \D_UU_AMIGA_in_0\ : std_logic;
signal \un1_D_UU_AMIGA_0\ : std_logic;
signal \D_UU_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\ : std_logic;
signal \un1_D_UU_AMIGA_1\ : std_logic;
signal \D_UM_AMIGA_in_5\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\ : std_logic;
signal \un1_D_UM_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\ : std_logic;
signal \D_UU_AMIGA_in_4\ : std_logic;
signal \un1_D_UU_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLEZ0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\ : std_logic;
signal \D_UU_AMIGA_in_7\ : std_logic;
signal \un1_D_UU_AMIGA_7\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \CPUBGn_wire\ : std_logic;
signal \TEA_CPUn_wire\ : std_logic;
signal \A_040_wire\ : std_logic_vector(1 downto 0);
signal \A_AMIGA_wire\ : std_logic_vector(1 downto 0);
signal \CLK40B_wire\ : std_logic;
signal \TBI_CPUn_wire\ : std_logic;
signal \CLK40A_wire\ : std_logic;
signal \BUFDIR_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \TS_CPUn_wire\ : std_logic;
signal \CLKRAMA_wire\ : std_logic;
signal \TCI_CPUn_wire\ : std_logic;
signal \CLKRAMB_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \TAn_wire\ : std_logic;
signal \DMAn_wire\ : std_logic;
signal \CLK80_CPU_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \pll_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \TACKn_wire\ <= TACKn;
    CPUBGn <= \CPUBGn_wire\;
    TEA_CPUn <= \TEA_CPUn_wire\;
    \A_040_wire\ <= A_040;
    A_AMIGA <= \A_AMIGA_wire\;
    CLK40B <= \CLK40B_wire\;
    TBI_CPUn <= \TBI_CPUn_wire\;
    CLK40A <= \CLK40A_wire\;
    BUFDIR <= \BUFDIR_wire\;
    \SIZ_wire\ <= SIZ;
    \TS_CPUn_wire\ <= TS_CPUn;
    CLKRAMA <= \CLKRAMA_wire\;
    TCI_CPUn <= \TCI_CPUn_wire\;
    CLKRAMB <= \CLKRAMB_wire\;
    BUFENn <= \BUFENn_wire\;
    \RnW_wire\ <= RnW;
    TAn <= \TAn_wire\;
    DMAn <= \DMAn_wire\;
    CLK80_CPU <= \CLK80_CPU_wire\;
    TSn <= \TSn_wire\;
    \PORTSIZE_wire\ <= PORTSIZE;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    \pll_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_pll\ : PLL40_2F
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            SCLK => '0',
            PLLOUTGLOBALA => \CLK80\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALB => \CLK40\,
            SDI => '0',
            PLLOUTCOREA => OPEN,
            BYPASS => '0',
            RESETB => \N__4989\,
            PLLOUTCOREB => OPEN,
            LOCK => OPEN,
            SDO => OPEN,
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \pll_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__8315\
        );

    \pll_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__8315\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \D_UM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8299\,
            DIN => \N__8298\,
            DOUT => \N__8297\,
            PACKAGEPIN => D_UM_040(3)
        );

    \D_UM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8299\,
            PADOUT => \N__8298\,
            PADIN => \N__8297\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5832\,
            DIN0 => \D_UM_040_in_3\,
            DOUT0 => \N__6801\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8290\,
            DIN => \N__8289\,
            DOUT => \N__8288\,
            PACKAGEPIN => D_LL_AMIGA(1)
        );

    \D_LL_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8290\,
            PADOUT => \N__8289\,
            PADIN => \N__8288\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2460\,
            DIN0 => \D_LL_AMIGA_in_1\,
            DOUT0 => \N__2802\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8281\,
            DIN => \N__8280\,
            DOUT => \N__8279\,
            PACKAGEPIN => D_UU_AMIGA(5)
        );

    \D_UU_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8281\,
            PADOUT => \N__8280\,
            PADIN => \N__8279\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2558\,
            DIN0 => \D_UU_AMIGA_in_5\,
            DOUT0 => \N__4278\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8272\,
            DIN => \N__8271\,
            DOUT => \N__8270\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8272\,
            PADOUT => \N__8271\,
            PADIN => \N__8270\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TACKn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8263\,
            DIN => \N__8262\,
            DOUT => \N__8261\,
            PACKAGEPIN => D_UU_040(6)
        );

    \D_UU_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8263\,
            PADOUT => \N__8262\,
            PADIN => \N__8261\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5936\,
            DIN0 => \D_UU_040_in_6\,
            DOUT0 => \N__4206\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUBGn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8254\,
            DIN => \N__8253\,
            DOUT => \N__8252\,
            PACKAGEPIN => \CPUBGn_wire\
        );

    \CPUBGn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8254\,
            PADOUT => \N__8253\,
            PADIN => \N__8252\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8245\,
            DIN => \N__8244\,
            DOUT => \N__8243\,
            PACKAGEPIN => D_LL_040(7)
        );

    \D_LL_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8245\,
            PADOUT => \N__8244\,
            PADIN => \N__8243\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5948\,
            DIN0 => \D_LL_040_in_7\,
            DOUT0 => \N__2823\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8236\,
            DIN => \N__8235\,
            DOUT => \N__8234\,
            PACKAGEPIN => D_LL_AMIGA(4)
        );

    \D_LL_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8236\,
            PADOUT => \N__8235\,
            PADIN => \N__8234\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2459\,
            DIN0 => \D_LL_AMIGA_in_4\,
            DOUT0 => \N__3069\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8227\,
            DIN => \N__8226\,
            DOUT => \N__8225\,
            PACKAGEPIN => D_UM_AMIGA(3)
        );

    \D_UM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8227\,
            PADOUT => \N__8226\,
            PADIN => \N__8225\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2543\,
            DIN0 => \D_UM_AMIGA_in_3\,
            DOUT0 => \N__3732\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8218\,
            DIN => \N__8217\,
            DOUT => \N__8216\,
            PACKAGEPIN => D_UU_040(3)
        );

    \D_UU_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8218\,
            PADOUT => \N__8217\,
            PADIN => \N__8216\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5885\,
            DIN0 => \D_UU_040_in_3\,
            DOUT0 => \N__6486\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEA_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8209\,
            DIN => \N__8208\,
            DOUT => \N__8207\,
            PACKAGEPIN => \TEA_CPUn_wire\
        );

    \TEA_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8209\,
            PADOUT => \N__8208\,
            PADIN => \N__8207\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4990\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8200\,
            DIN => \N__8199\,
            DOUT => \N__8198\,
            PACKAGEPIN => \A_040_wire\(1)
        );

    \A_040_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8200\,
            PADOUT => \N__8199\,
            PADIN => \N__8198\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8191\,
            DIN => \N__8190\,
            DOUT => \N__8189\,
            PACKAGEPIN => D_LM_AMIGA(3)
        );

    \D_LM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8191\,
            PADOUT => \N__8190\,
            PADIN => \N__8189\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2427\,
            DIN0 => \D_LM_AMIGA_in_3\,
            DOUT0 => \N__2985\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8182\,
            DIN => \N__8181\,
            DOUT => \N__8180\,
            PACKAGEPIN => D_LM_040(0)
        );

    \D_LM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8182\,
            PADOUT => \N__8181\,
            PADIN => \N__8180\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5949\,
            DIN0 => \D_LM_040_in_0\,
            DOUT0 => \N__4176\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8173\,
            DIN => \N__8172\,
            DOUT => \N__8171\,
            PACKAGEPIN => D_UM_AMIGA(6)
        );

    \D_UM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8173\,
            PADOUT => \N__8172\,
            PADIN => \N__8171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2557\,
            DIN0 => \D_UM_AMIGA_in_6\,
            DOUT0 => \N__3108\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8164\,
            DIN => \N__8163\,
            DOUT => \N__8162\,
            PACKAGEPIN => D_LM_AMIGA(4)
        );

    \D_LM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8164\,
            PADOUT => \N__8163\,
            PADIN => \N__8162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2472\,
            DIN0 => \D_LM_AMIGA_in_4\,
            DOUT0 => \N__3381\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8155\,
            DIN => \N__8154\,
            DOUT => \N__8153\,
            PACKAGEPIN => \A_AMIGA_wire\(1)
        );

    \A_AMIGA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8155\,
            PADOUT => \N__8154\,
            PADIN => \N__8153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4400\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8146\,
            DIN => \N__8145\,
            DOUT => \N__8144\,
            PACKAGEPIN => D_LM_040(7)
        );

    \D_LM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8146\,
            PADOUT => \N__8145\,
            PADIN => \N__8144\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5749\,
            DIN0 => \D_LM_040_in_7\,
            DOUT0 => \N__4920\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8137\,
            DIN => \N__8136\,
            DOUT => \N__8135\,
            PACKAGEPIN => D_UM_040(4)
        );

    \D_UM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8137\,
            PADOUT => \N__8136\,
            PADIN => \N__8135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5886\,
            DIN0 => \D_UM_040_in_4\,
            DOUT0 => \N__6639\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8128\,
            DIN => \N__8127\,
            DOUT => \N__8126\,
            PACKAGEPIN => \CLK40B_wire\
        );

    \CLK40B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8128\,
            PADOUT => \N__8127\,
            PADIN => \N__8126\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5478\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8119\,
            DIN => \N__8118\,
            DOUT => \N__8117\,
            PACKAGEPIN => D_UU_AMIGA(0)
        );

    \D_UU_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8119\,
            PADOUT => \N__8118\,
            PADIN => \N__8117\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2407\,
            DIN0 => \D_UU_AMIGA_in_0\,
            DOUT0 => \N__4743\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8110\,
            DIN => \N__8109\,
            DOUT => \N__8108\,
            PACKAGEPIN => \A_040_wire\(0)
        );

    \A_040_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8110\,
            PADOUT => \N__8109\,
            PADIN => \N__8108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8101\,
            DIN => \N__8100\,
            DOUT => \N__8099\,
            PACKAGEPIN => D_LM_AMIGA(0)
        );

    \D_LM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8101\,
            PADOUT => \N__8100\,
            PADIN => \N__8099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2409\,
            DIN0 => \D_LM_AMIGA_in_0\,
            DOUT0 => \N__4797\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8092\,
            DIN => \N__8091\,
            DOUT => \N__8090\,
            PACKAGEPIN => D_UM_040(1)
        );

    \D_UM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8092\,
            PADOUT => \N__8091\,
            PADIN => \N__8090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5830\,
            DIN0 => \D_UM_040_in_1\,
            DOUT0 => \N__6882\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8083\,
            DIN => \N__8082\,
            DOUT => \N__8081\,
            PACKAGEPIN => \TBI_CPUn_wire\
        );

    \TBI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8083\,
            PADOUT => \N__8082\,
            PADIN => \N__8081\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5430\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8074\,
            DIN => \N__8073\,
            DOUT => \N__8072\,
            PACKAGEPIN => \CLK40A_wire\
        );

    \CLK40A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8074\,
            PADOUT => \N__8073\,
            PADIN => \N__8072\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5477\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8065\,
            DIN => \N__8064\,
            DOUT => \N__8063\,
            PACKAGEPIN => D_LM_040(3)
        );

    \D_LM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8065\,
            PADOUT => \N__8064\,
            PADIN => \N__8063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5911\,
            DIN0 => \D_LM_040_in_3\,
            DOUT0 => \N__3459\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8056\,
            DIN => \N__8055\,
            DOUT => \N__8054\,
            PACKAGEPIN => D_LL_040(4)
        );

    \D_LL_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8056\,
            PADOUT => \N__8055\,
            PADIN => \N__8054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5983\,
            DIN0 => \D_LL_040_in_4\,
            DOUT0 => \N__3573\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8047\,
            DIN => \N__8046\,
            DOUT => \N__8045\,
            PACKAGEPIN => D_LL_AMIGA(7)
        );

    \D_LL_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8047\,
            PADOUT => \N__8046\,
            PADIN => \N__8045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2408\,
            DIN0 => \D_LL_AMIGA_in_7\,
            DOUT0 => \N__4875\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8038\,
            DIN => \N__8037\,
            DOUT => \N__8036\,
            PACKAGEPIN => D_UU_AMIGA(7)
        );

    \D_UU_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8038\,
            PADOUT => \N__8037\,
            PADIN => \N__8036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2555\,
            DIN0 => \D_UU_AMIGA_in_7\,
            DOUT0 => \N__2655\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8029\,
            DIN => \N__8028\,
            DOUT => \N__8027\,
            PACKAGEPIN => \BUFDIR_wire\
        );

    \BUFDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8029\,
            PADOUT => \N__8028\,
            PADIN => \N__8027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5967\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8020\,
            DIN => \N__8019\,
            DOUT => \N__8018\,
            PACKAGEPIN => D_LM_AMIGA(5)
        );

    \D_LM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8020\,
            PADOUT => \N__8019\,
            PADIN => \N__8018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2511\,
            DIN0 => \D_LM_AMIGA_in_5\,
            DOUT0 => \N__4617\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8011\,
            DIN => \N__8010\,
            DOUT => \N__8009\,
            PACKAGEPIN => D_UU_040(4)
        );

    \D_UU_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8011\,
            PADOUT => \N__8010\,
            PADIN => \N__8009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5939\,
            DIN0 => \D_UU_040_in_4\,
            DOUT0 => \N__6900\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8002\,
            DIN => \N__8001\,
            DOUT => \N__8000\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8002\,
            PADOUT => \N__8001\,
            PADIN => \N__8000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7993\,
            DIN => \N__7992\,
            DOUT => \N__7991\,
            PACKAGEPIN => D_LM_040(6)
        );

    \D_LM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7993\,
            PADOUT => \N__7992\,
            PADIN => \N__7991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5744\,
            DIN0 => \D_LM_040_in_6\,
            DOUT0 => \N__3228\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7984\,
            DIN => \N__7983\,
            DOUT => \N__7982\,
            PACKAGEPIN => D_UM_040(5)
        );

    \D_UM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7984\,
            PADOUT => \N__7983\,
            PADIN => \N__7982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5887\,
            DIN0 => \D_UM_040_in_5\,
            DOUT0 => \N__6981\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TS_CPUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7975\,
            DIN => \N__7974\,
            DOUT => \N__7973\,
            PACKAGEPIN => \TS_CPUn_wire\
        );

    \TS_CPUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7975\,
            PADOUT => \N__7974\,
            PADIN => \N__7973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TS_CPUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7966\,
            DIN => \N__7965\,
            DOUT => \N__7964\,
            PACKAGEPIN => D_LL_040(1)
        );

    \D_LL_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7966\,
            PADOUT => \N__7965\,
            PADIN => \N__7964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5982\,
            DIN0 => \D_LL_040_in_1\,
            DOUT0 => \N__3654\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7957\,
            DIN => \N__7956\,
            DOUT => \N__7955\,
            PACKAGEPIN => D_LL_AMIGA(3)
        );

    \D_LL_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7957\,
            PADOUT => \N__7956\,
            PADIN => \N__7955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2508\,
            DIN0 => \D_LL_AMIGA_in_3\,
            DOUT0 => \N__3800\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7948\,
            DIN => \N__7947\,
            DOUT => \N__7946\,
            PACKAGEPIN => D_UM_AMIGA(5)
        );

    \D_UM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7948\,
            PADOUT => \N__7947\,
            PADIN => \N__7946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2535\,
            DIN0 => \D_UM_AMIGA_in_5\,
            DOUT0 => \N__4659\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7939\,
            DIN => \N__7938\,
            DOUT => \N__7937\,
            PACKAGEPIN => D_UU_040(1)
        );

    \D_UU_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7939\,
            PADOUT => \N__7938\,
            PADIN => \N__7937\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5833\,
            DIN0 => \D_UU_040_in_1\,
            DOUT0 => \N__7059\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7930\,
            DIN => \N__7929\,
            DOUT => \N__7928\,
            PACKAGEPIN => D_UU_AMIGA(3)
        );

    \D_UU_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7930\,
            PADOUT => \N__7929\,
            PADIN => \N__7928\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2559\,
            DIN0 => \D_UU_AMIGA_in_3\,
            DOUT0 => \N__2940\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7921\,
            DIN => \N__7920\,
            DOUT => \N__7919\,
            PACKAGEPIN => D_LM_AMIGA(1)
        );

    \D_LM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7921\,
            PADOUT => \N__7920\,
            PADIN => \N__7919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2426\,
            DIN0 => \D_LM_AMIGA_in_1\,
            DOUT0 => \N__3987\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7912\,
            DIN => \N__7911\,
            DOUT => \N__7910\,
            PACKAGEPIN => D_LM_040(2)
        );

    \D_LM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7912\,
            PADOUT => \N__7911\,
            PADIN => \N__7910\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5947\,
            DIN0 => \D_LM_040_in_2\,
            DOUT0 => \N__3264\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7903\,
            DIN => \N__7902\,
            DOUT => \N__7901\,
            PACKAGEPIN => D_LL_040(5)
        );

    \D_LL_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7903\,
            PADOUT => \N__7902\,
            PADIN => \N__7901\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5950\,
            DIN0 => \D_LL_040_in_5\,
            DOUT0 => \N__3612\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7894\,
            DIN => \N__7893\,
            DOUT => \N__7892\,
            PACKAGEPIN => D_LL_AMIGA(6)
        );

    \D_LL_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7894\,
            PADOUT => \N__7893\,
            PADIN => \N__7892\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2410\,
            DIN0 => \D_LL_AMIGA_in_6\,
            DOUT0 => \N__3156\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7885\,
            DIN => \N__7884\,
            DOUT => \N__7883\,
            PACKAGEPIN => D_UU_AMIGA(6)
        );

    \D_UU_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7885\,
            PADOUT => \N__7884\,
            PADIN => \N__7883\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2556\,
            DIN0 => \D_UU_AMIGA_in_6\,
            DOUT0 => \N__2856\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7876\,
            DIN => \N__7875\,
            DOUT => \N__7874\,
            PACKAGEPIN => D_UM_AMIGA(1)
        );

    \D_UM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7876\,
            PADOUT => \N__7875\,
            PADIN => \N__7874\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2512\,
            DIN0 => \D_UM_AMIGA_in_1\,
            DOUT0 => \N__2736\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7867\,
            DIN => \N__7866\,
            DOUT => \N__7865\,
            PACKAGEPIN => D_UU_040(5)
        );

    \D_UU_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7867\,
            PADOUT => \N__7866\,
            PADIN => \N__7865\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5888\,
            DIN0 => \D_UU_040_in_5\,
            DOUT0 => \N__6561\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7858\,
            DIN => \N__7857\,
            DOUT => \N__7856\,
            PACKAGEPIN => \CLKRAMA_wire\
        );

    \CLKRAMA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7858\,
            PADOUT => \N__7857\,
            PADIN => \N__7856\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6195\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7849\,
            DIN => \N__7848\,
            DOUT => \N__7847\,
            PACKAGEPIN => D_UM_040(2)
        );

    \D_UM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7849\,
            PADOUT => \N__7848\,
            PADIN => \N__7847\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5777\,
            DIN0 => \D_UM_040_in_2\,
            DOUT0 => \N__6465\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7840\,
            DIN => \N__7839\,
            DOUT => \N__7838\,
            PACKAGEPIN => D_LL_040(2)
        );

    \D_LL_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7840\,
            PADOUT => \N__7839\,
            PADIN => \N__7838\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5968\,
            DIN0 => \D_LL_040_in_2\,
            DOUT0 => \N__2583\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7831\,
            DIN => \N__7830\,
            DOUT => \N__7829\,
            PACKAGEPIN => \TCI_CPUn_wire\
        );

    \TCI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7831\,
            PADOUT => \N__7830\,
            PADIN => \N__7829\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4994\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7822\,
            DIN => \N__7821\,
            DOUT => \N__7820\,
            PACKAGEPIN => \CLKRAMB_wire\
        );

    \CLKRAMB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7822\,
            PADOUT => \N__7821\,
            PADIN => \N__7820\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6188\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7813\,
            DIN => \N__7812\,
            DOUT => \N__7811\,
            PACKAGEPIN => D_LL_AMIGA(2)
        );

    \D_LL_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7813\,
            PADOUT => \N__7812\,
            PADIN => \N__7811\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2509\,
            DIN0 => \D_LL_AMIGA_in_2\,
            DOUT0 => \N__3534\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7804\,
            DIN => \N__7803\,
            DOUT => \N__7802\,
            PACKAGEPIN => D_UM_AMIGA(4)
        );

    \D_UM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7804\,
            PADOUT => \N__7803\,
            PADIN => \N__7802\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2545\,
            DIN0 => \D_UM_AMIGA_in_4\,
            DOUT0 => \N__3027\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7795\,
            DIN => \N__7794\,
            DOUT => \N__7793\,
            PACKAGEPIN => D_UU_AMIGA(2)
        );

    \D_UU_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7795\,
            PADOUT => \N__7794\,
            PADIN => \N__7793\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2406\,
            DIN0 => \D_UU_AMIGA_in_2\,
            DOUT0 => \N__3867\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7786\,
            DIN => \N__7785\,
            DOUT => \N__7784\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7786\,
            PADOUT => \N__7785\,
            PADIN => \N__7784\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7777\,
            DIN => \N__7776\,
            DOUT => \N__7775\,
            PACKAGEPIN => D_LM_AMIGA(6)
        );

    \D_LM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7777\,
            PADOUT => \N__7776\,
            PADIN => \N__7775\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2514\,
            DIN0 => \D_LM_AMIGA_in_6\,
            DOUT0 => \N__2919\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7768\,
            DIN => \N__7767\,
            DOUT => \N__7766\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7768\,
            PADOUT => \N__7767\,
            PADIN => \N__7766\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7759\,
            DIN => \N__7758\,
            DOUT => \N__7757\,
            PACKAGEPIN => D_LM_040(5)
        );

    \D_LM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7759\,
            PADOUT => \N__7758\,
            PADIN => \N__7757\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5821\,
            DIN0 => \D_LM_040_in_5\,
            DOUT0 => \N__3426\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7750\,
            DIN => \N__7749\,
            DOUT => \N__7748\,
            PACKAGEPIN => D_UM_040(6)
        );

    \D_UM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7750\,
            PADOUT => \N__7749\,
            PADIN => \N__7748\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5748\,
            DIN0 => \D_UM_040_in_6\,
            DOUT0 => \N__6009\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7741\,
            DIN => \N__7740\,
            DOUT => \N__7739\,
            PACKAGEPIN => \TAn_wire\
        );

    \TAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7741\,
            PADOUT => \N__7740\,
            PADIN => \N__7739\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5429\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMAn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7732\,
            DIN => \N__7731\,
            DOUT => \N__7730\,
            PACKAGEPIN => \DMAn_wire\
        );

    \DMAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7732\,
            PADOUT => \N__7731\,
            PADIN => \N__7730\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4998\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7723\,
            DIN => \N__7722\,
            DOUT => \N__7721\,
            PACKAGEPIN => D_LL_040(6)
        );

    \D_LL_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7723\,
            PADOUT => \N__7722\,
            PADIN => \N__7721\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5951\,
            DIN0 => \D_LL_040_in_6\,
            DOUT0 => \N__3825\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7714\,
            DIN => \N__7713\,
            DOUT => \N__7712\,
            PACKAGEPIN => D_LL_AMIGA(5)
        );

    \D_LL_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7714\,
            PADOUT => \N__7713\,
            PADIN => \N__7712\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2411\,
            DIN0 => \D_LL_AMIGA_in_5\,
            DOUT0 => \N__4725\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7705\,
            DIN => \N__7704\,
            DOUT => \N__7703\,
            PACKAGEPIN => D_UM_AMIGA(0)
        );

    \D_UM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7705\,
            PADOUT => \N__7704\,
            PADIN => \N__7703\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2471\,
            DIN0 => \D_UM_AMIGA_in_0\,
            DOUT0 => \N__2238\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7696\,
            DIN => \N__7695\,
            DOUT => \N__7694\,
            PACKAGEPIN => D_UU_040(2)
        );

    \D_UU_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7696\,
            PADOUT => \N__7695\,
            PADIN => \N__7694\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5938\,
            DIN0 => \D_UU_040_in_2\,
            DOUT0 => \N__5493\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7687\,
            DIN => \N__7686\,
            DOUT => \N__7685\,
            PACKAGEPIN => D_LM_AMIGA(2)
        );

    \D_LM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7687\,
            PADOUT => \N__7686\,
            PADIN => \N__7685\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2470\,
            DIN0 => \D_LM_AMIGA_in_2\,
            DOUT0 => \N__3905\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK80_CPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7678\,
            DIN => \N__7677\,
            DOUT => \N__7676\,
            PACKAGEPIN => \CLK80_CPU_wire\
        );

    \CLK80_CPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7678\,
            PADOUT => \N__7677\,
            PADIN => \N__7676\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6187\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7669\,
            DIN => \N__7668\,
            DOUT => \N__7667\,
            PACKAGEPIN => D_LL_040(3)
        );

    \D_LL_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7669\,
            PADOUT => \N__7668\,
            PADIN => \N__7667\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5984\,
            DIN0 => \D_LL_040_in_3\,
            DOUT0 => \N__3693\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7660\,
            DIN => \N__7659\,
            DOUT => \N__7658\,
            PACKAGEPIN => D_LM_040(1)
        );

    \D_LM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7660\,
            PADOUT => \N__7659\,
            PADIN => \N__7658\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5946\,
            DIN0 => \D_LM_040_in_1\,
            DOUT0 => \N__3195\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7651\,
            DIN => \N__7650\,
            DOUT => \N__7649\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7651\,
            PADOUT => \N__7650\,
            PADIN => \N__7649\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3291\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7642\,
            DIN => \N__7641\,
            DOUT => \N__7640\,
            PACKAGEPIN => D_UM_AMIGA(7)
        );

    \D_UM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7642\,
            PADOUT => \N__7641\,
            PADIN => \N__7640\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2544\,
            DIN0 => \D_UM_AMIGA_in_7\,
            DOUT0 => \N__4830\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7633\,
            DIN => \N__7632\,
            DOUT => \N__7631\,
            PACKAGEPIN => D_LM_AMIGA(7)
        );

    \D_LM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7633\,
            PADOUT => \N__7632\,
            PADIN => \N__7631\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2513\,
            DIN0 => \D_LM_AMIGA_in_7\,
            DOUT0 => \N__2700\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7624\,
            DIN => \N__7623\,
            DOUT => \N__7622\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7624\,
            PADOUT => \N__7623\,
            PADIN => \N__7622\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PORTSIZE_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7615\,
            DIN => \N__7614\,
            DOUT => \N__7613\,
            PACKAGEPIN => \A_AMIGA_wire\(0)
        );

    \A_AMIGA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7615\,
            PADOUT => \N__7614\,
            PADIN => \N__7613\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2622\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7606\,
            DIN => \N__7605\,
            DOUT => \N__7604\,
            PACKAGEPIN => D_LM_040(4)
        );

    \D_LM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7606\,
            PADOUT => \N__7605\,
            PADIN => \N__7604\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5866\,
            DIN0 => \D_LM_040_in_4\,
            DOUT0 => \N__4032\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7597\,
            DIN => \N__7596\,
            DOUT => \N__7595\,
            PACKAGEPIN => D_UM_040(7)
        );

    \D_UM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7597\,
            PADOUT => \N__7596\,
            PADIN => \N__7595\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5831\,
            DIN0 => \D_UM_040_in_7\,
            DOUT0 => \N__6717\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7588\,
            DIN => \N__7587\,
            DOUT => \N__7586\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7588\,
            PADOUT => \N__7587\,
            PADIN => \N__7586\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7579\,
            DIN => \N__7578\,
            DOUT => \N__7577\,
            PACKAGEPIN => D_UU_AMIGA(1)
        );

    \D_UU_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7579\,
            PADOUT => \N__7578\,
            PADIN => \N__7577\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2542\,
            DIN0 => \D_UU_AMIGA_in_1\,
            DOUT0 => \N__3945\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7570\,
            DIN => \N__7569\,
            DOUT => \N__7568\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7570\,
            PADOUT => \N__7569\,
            PADIN => \N__7568\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5476\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7561\,
            DIN => \N__7560\,
            DOUT => \N__7559\,
            PACKAGEPIN => D_UM_040(0)
        );

    \D_UM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7561\,
            PADOUT => \N__7560\,
            PADIN => \N__7559\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5820\,
            DIN0 => \D_UM_040_in_0\,
            DOUT0 => \N__4155\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7552\,
            DIN => \N__7551\,
            DOUT => \N__7550\,
            PACKAGEPIN => D_LL_AMIGA(0)
        );

    \D_LL_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7552\,
            PADOUT => \N__7551\,
            PADIN => \N__7550\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2510\,
            DIN0 => \D_LL_AMIGA_in_0\,
            DOUT0 => \N__2283\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7543\,
            DIN => \N__7542\,
            DOUT => \N__7541\,
            PACKAGEPIN => D_UU_AMIGA(4)
        );

    \D_UU_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7543\,
            PADOUT => \N__7542\,
            PADIN => \N__7541\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2534\,
            DIN0 => \D_UU_AMIGA_in_4\,
            DOUT0 => \N__3342\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7534\,
            DIN => \N__7533\,
            DOUT => \N__7532\,
            PACKAGEPIN => D_UU_040(7)
        );

    \D_UU_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7534\,
            PADOUT => \N__7533\,
            PADIN => \N__7532\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5935\,
            DIN0 => \D_UU_040_in_7\,
            DOUT0 => \N__7290\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7525\,
            DIN => \N__7524\,
            DOUT => \N__7523\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7525\,
            PADOUT => \N__7524\,
            PADIN => \N__7523\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7516\,
            DIN => \N__7515\,
            DOUT => \N__7514\,
            PACKAGEPIN => D_LL_040(0)
        );

    \D_LL_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7516\,
            PADOUT => \N__7515\,
            PADIN => \N__7514\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5985\,
            DIN0 => \D_LL_040_in_0\,
            DOUT0 => \N__3312\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7507\,
            DIN => \N__7506\,
            DOUT => \N__7505\,
            PACKAGEPIN => D_UM_AMIGA(2)
        );

    \D_UM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7507\,
            PADOUT => \N__7506\,
            PADIN => \N__7505\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2473\,
            DIN0 => \D_UM_AMIGA_in_2\,
            DOUT0 => \N__3492\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7498\,
            DIN => \N__7497\,
            DOUT => \N__7496\,
            PACKAGEPIN => D_UU_040(0)
        );

    \D_UU_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7498\,
            PADOUT => \N__7497\,
            PADIN => \N__7496\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5937\,
            DIN0 => \D_UU_040_in_0\,
            DOUT0 => \N__7134\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1948\ : InMux
    port map (
            O => \N__7479\,
            I => \N__7473\
        );

    \I__1947\ : InMux
    port map (
            O => \N__7478\,
            I => \N__7473\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__7473\,
            I => \N__7457\
        );

    \I__1945\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7450\
        );

    \I__1944\ : InMux
    port map (
            O => \N__7471\,
            I => \N__7450\
        );

    \I__1943\ : InMux
    port map (
            O => \N__7470\,
            I => \N__7450\
        );

    \I__1942\ : InMux
    port map (
            O => \N__7469\,
            I => \N__7445\
        );

    \I__1941\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7445\
        );

    \I__1940\ : InMux
    port map (
            O => \N__7467\,
            I => \N__7440\
        );

    \I__1939\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7440\
        );

    \I__1938\ : InMux
    port map (
            O => \N__7465\,
            I => \N__7435\
        );

    \I__1937\ : InMux
    port map (
            O => \N__7464\,
            I => \N__7435\
        );

    \I__1936\ : InMux
    port map (
            O => \N__7463\,
            I => \N__7430\
        );

    \I__1935\ : InMux
    port map (
            O => \N__7462\,
            I => \N__7430\
        );

    \I__1934\ : InMux
    port map (
            O => \N__7461\,
            I => \N__7427\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__7460\,
            I => \N__7420\
        );

    \I__1932\ : Sp12to4
    port map (
            O => \N__7457\,
            I => \N__7416\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__7450\,
            I => \N__7411\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__7445\,
            I => \N__7411\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__7440\,
            I => \N__7404\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__7435\,
            I => \N__7404\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__7430\,
            I => \N__7404\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__7427\,
            I => \N__7401\
        );

    \I__1925\ : InMux
    port map (
            O => \N__7426\,
            I => \N__7398\
        );

    \I__1924\ : InMux
    port map (
            O => \N__7425\,
            I => \N__7395\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__7424\,
            I => \N__7392\
        );

    \I__1922\ : InMux
    port map (
            O => \N__7423\,
            I => \N__7389\
        );

    \I__1921\ : InMux
    port map (
            O => \N__7420\,
            I => \N__7384\
        );

    \I__1920\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7384\
        );

    \I__1919\ : Span12Mux_v
    port map (
            O => \N__7416\,
            I => \N__7380\
        );

    \I__1918\ : Span4Mux_v
    port map (
            O => \N__7411\,
            I => \N__7377\
        );

    \I__1917\ : Span4Mux_v
    port map (
            O => \N__7404\,
            I => \N__7368\
        );

    \I__1916\ : Span4Mux_v
    port map (
            O => \N__7401\,
            I => \N__7368\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__7398\,
            I => \N__7368\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__7395\,
            I => \N__7368\
        );

    \I__1913\ : InMux
    port map (
            O => \N__7392\,
            I => \N__7365\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__7389\,
            I => \N__7360\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__7384\,
            I => \N__7360\
        );

    \I__1910\ : InMux
    port map (
            O => \N__7383\,
            I => \N__7357\
        );

    \I__1909\ : Odrv12
    port map (
            O => \N__7380\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__7377\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__7368\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__7365\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__7360\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__7357\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1903\ : InMux
    port map (
            O => \N__7344\,
            I => \N__7341\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__7341\,
            I => \N__7338\
        );

    \I__1901\ : Odrv12
    port map (
            O => \N__7338\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__1900\ : InMux
    port map (
            O => \N__7335\,
            I => \N__7331\
        );

    \I__1899\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7328\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__7331\,
            I => \N__7324\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__7328\,
            I => \N__7321\
        );

    \I__1896\ : InMux
    port map (
            O => \N__7327\,
            I => \N__7318\
        );

    \I__1895\ : Span4Mux_v
    port map (
            O => \N__7324\,
            I => \N__7315\
        );

    \I__1894\ : Span4Mux_v
    port map (
            O => \N__7321\,
            I => \N__7312\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__7318\,
            I => \N__7309\
        );

    \I__1892\ : Span4Mux_h
    port map (
            O => \N__7315\,
            I => \N__7306\
        );

    \I__1891\ : Span4Mux_v
    port map (
            O => \N__7312\,
            I => \N__7301\
        );

    \I__1890\ : Span4Mux_v
    port map (
            O => \N__7309\,
            I => \N__7301\
        );

    \I__1889\ : Sp12to4
    port map (
            O => \N__7306\,
            I => \N__7296\
        );

    \I__1888\ : Sp12to4
    port map (
            O => \N__7301\,
            I => \N__7296\
        );

    \I__1887\ : Span12Mux_h
    port map (
            O => \N__7296\,
            I => \N__7293\
        );

    \I__1886\ : Odrv12
    port map (
            O => \N__7293\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__1885\ : IoInMux
    port map (
            O => \N__7290\,
            I => \N__7287\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__7287\,
            I => \N__7284\
        );

    \I__1883\ : Span12Mux_s11_v
    port map (
            O => \N__7284\,
            I => \N__7281\
        );

    \I__1882\ : Span12Mux_h
    port map (
            O => \N__7281\,
            I => \N__7278\
        );

    \I__1881\ : Odrv12
    port map (
            O => \N__7278\,
            I => \un1_D_UU_AMIGA_7\
        );

    \I__1880\ : CEMux
    port map (
            O => \N__7275\,
            I => \N__7268\
        );

    \I__1879\ : CEMux
    port map (
            O => \N__7274\,
            I => \N__7265\
        );

    \I__1878\ : CEMux
    port map (
            O => \N__7273\,
            I => \N__7262\
        );

    \I__1877\ : CEMux
    port map (
            O => \N__7272\,
            I => \N__7259\
        );

    \I__1876\ : CEMux
    port map (
            O => \N__7271\,
            I => \N__7256\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__7268\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__7265\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__7262\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__7259\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__7256\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1870\ : SRMux
    port map (
            O => \N__7245\,
            I => \N__7240\
        );

    \I__1869\ : SRMux
    port map (
            O => \N__7244\,
            I => \N__7237\
        );

    \I__1868\ : SRMux
    port map (
            O => \N__7243\,
            I => \N__7233\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__7240\,
            I => \N__7229\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__7237\,
            I => \N__7226\
        );

    \I__1865\ : SRMux
    port map (
            O => \N__7236\,
            I => \N__7223\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__7233\,
            I => \N__7220\
        );

    \I__1863\ : SRMux
    port map (
            O => \N__7232\,
            I => \N__7217\
        );

    \I__1862\ : Span4Mux_v
    port map (
            O => \N__7229\,
            I => \N__7212\
        );

    \I__1861\ : Span4Mux_v
    port map (
            O => \N__7226\,
            I => \N__7212\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__7223\,
            I => \N__7205\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__7220\,
            I => \N__7205\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__7217\,
            I => \N__7205\
        );

    \I__1857\ : Span4Mux_h
    port map (
            O => \N__7212\,
            I => \N__7202\
        );

    \I__1856\ : Span4Mux_v
    port map (
            O => \N__7205\,
            I => \N__7199\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__7202\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__7199\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\
        );

    \I__1853\ : InMux
    port map (
            O => \N__7194\,
            I => \N__7191\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__7191\,
            I => \N__7188\
        );

    \I__1851\ : Odrv12
    port map (
            O => \N__7188\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__7185\,
            I => \N__7182\
        );

    \I__1849\ : InMux
    port map (
            O => \N__7182\,
            I => \N__7179\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__7179\,
            I => \N__7175\
        );

    \I__1847\ : InMux
    port map (
            O => \N__7178\,
            I => \N__7172\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__7175\,
            I => \N__7168\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__7172\,
            I => \N__7165\
        );

    \I__1844\ : InMux
    port map (
            O => \N__7171\,
            I => \N__7162\
        );

    \I__1843\ : Span4Mux_v
    port map (
            O => \N__7168\,
            I => \N__7159\
        );

    \I__1842\ : Span4Mux_v
    port map (
            O => \N__7165\,
            I => \N__7154\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__7162\,
            I => \N__7154\
        );

    \I__1840\ : Sp12to4
    port map (
            O => \N__7159\,
            I => \N__7151\
        );

    \I__1839\ : Sp12to4
    port map (
            O => \N__7154\,
            I => \N__7148\
        );

    \I__1838\ : Span12Mux_h
    port map (
            O => \N__7151\,
            I => \N__7145\
        );

    \I__1837\ : Span12Mux_v
    port map (
            O => \N__7148\,
            I => \N__7142\
        );

    \I__1836\ : Span12Mux_v
    port map (
            O => \N__7145\,
            I => \N__7137\
        );

    \I__1835\ : Span12Mux_h
    port map (
            O => \N__7142\,
            I => \N__7137\
        );

    \I__1834\ : Odrv12
    port map (
            O => \N__7137\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1833\ : IoInMux
    port map (
            O => \N__7134\,
            I => \N__7131\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__7131\,
            I => \N__7128\
        );

    \I__1831\ : Span4Mux_s3_v
    port map (
            O => \N__7128\,
            I => \N__7125\
        );

    \I__1830\ : Span4Mux_h
    port map (
            O => \N__7125\,
            I => \N__7122\
        );

    \I__1829\ : Sp12to4
    port map (
            O => \N__7122\,
            I => \N__7119\
        );

    \I__1828\ : Span12Mux_s8_v
    port map (
            O => \N__7119\,
            I => \N__7116\
        );

    \I__1827\ : Odrv12
    port map (
            O => \N__7116\,
            I => \un1_D_UU_AMIGA_0\
        );

    \I__1826\ : InMux
    port map (
            O => \N__7113\,
            I => \N__7110\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__7110\,
            I => \N__7106\
        );

    \I__1824\ : InMux
    port map (
            O => \N__7109\,
            I => \N__7103\
        );

    \I__1823\ : Span4Mux_v
    port map (
            O => \N__7106\,
            I => \N__7099\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__7103\,
            I => \N__7096\
        );

    \I__1821\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7093\
        );

    \I__1820\ : Span4Mux_v
    port map (
            O => \N__7099\,
            I => \N__7090\
        );

    \I__1819\ : Span4Mux_v
    port map (
            O => \N__7096\,
            I => \N__7085\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__7093\,
            I => \N__7085\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__7090\,
            I => \N__7082\
        );

    \I__1816\ : Span4Mux_v
    port map (
            O => \N__7085\,
            I => \N__7079\
        );

    \I__1815\ : Sp12to4
    port map (
            O => \N__7082\,
            I => \N__7074\
        );

    \I__1814\ : Sp12to4
    port map (
            O => \N__7079\,
            I => \N__7074\
        );

    \I__1813\ : Span12Mux_h
    port map (
            O => \N__7074\,
            I => \N__7071\
        );

    \I__1812\ : Odrv12
    port map (
            O => \N__7071\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__1811\ : InMux
    port map (
            O => \N__7068\,
            I => \N__7065\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__7065\,
            I => \N__7062\
        );

    \I__1809\ : Odrv12
    port map (
            O => \N__7062\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__1808\ : IoInMux
    port map (
            O => \N__7059\,
            I => \N__7056\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__7056\,
            I => \N__7053\
        );

    \I__1806\ : IoSpan4Mux
    port map (
            O => \N__7053\,
            I => \N__7050\
        );

    \I__1805\ : IoSpan4Mux
    port map (
            O => \N__7050\,
            I => \N__7047\
        );

    \I__1804\ : Span4Mux_s2_h
    port map (
            O => \N__7047\,
            I => \N__7044\
        );

    \I__1803\ : Sp12to4
    port map (
            O => \N__7044\,
            I => \N__7041\
        );

    \I__1802\ : Odrv12
    port map (
            O => \N__7041\,
            I => \un1_D_UU_AMIGA_1\
        );

    \I__1801\ : InMux
    port map (
            O => \N__7038\,
            I => \N__7035\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__7035\,
            I => \N__7031\
        );

    \I__1799\ : InMux
    port map (
            O => \N__7034\,
            I => \N__7027\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__7031\,
            I => \N__7024\
        );

    \I__1797\ : InMux
    port map (
            O => \N__7030\,
            I => \N__7021\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__7027\,
            I => \N__7018\
        );

    \I__1795\ : Sp12to4
    port map (
            O => \N__7024\,
            I => \N__7015\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__7021\,
            I => \N__7012\
        );

    \I__1793\ : Span12Mux_v
    port map (
            O => \N__7018\,
            I => \N__7009\
        );

    \I__1792\ : Span12Mux_h
    port map (
            O => \N__7015\,
            I => \N__7006\
        );

    \I__1791\ : Span12Mux_s7_v
    port map (
            O => \N__7012\,
            I => \N__7003\
        );

    \I__1790\ : Span12Mux_h
    port map (
            O => \N__7009\,
            I => \N__7000\
        );

    \I__1789\ : Span12Mux_v
    port map (
            O => \N__7006\,
            I => \N__6995\
        );

    \I__1788\ : Span12Mux_h
    port map (
            O => \N__7003\,
            I => \N__6995\
        );

    \I__1787\ : Odrv12
    port map (
            O => \N__7000\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1786\ : Odrv12
    port map (
            O => \N__6995\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1785\ : InMux
    port map (
            O => \N__6990\,
            I => \N__6987\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__6987\,
            I => \N__6984\
        );

    \I__1783\ : Odrv12
    port map (
            O => \N__6984\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__1782\ : IoInMux
    port map (
            O => \N__6981\,
            I => \N__6978\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__6978\,
            I => \N__6975\
        );

    \I__1780\ : Span4Mux_s2_v
    port map (
            O => \N__6975\,
            I => \N__6972\
        );

    \I__1779\ : Span4Mux_h
    port map (
            O => \N__6972\,
            I => \N__6969\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__6969\,
            I => \N__6966\
        );

    \I__1777\ : Sp12to4
    port map (
            O => \N__6966\,
            I => \N__6963\
        );

    \I__1776\ : Odrv12
    port map (
            O => \N__6963\,
            I => \un1_D_UM_AMIGA_5\
        );

    \I__1775\ : InMux
    port map (
            O => \N__6960\,
            I => \N__6957\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__6957\,
            I => \N__6954\
        );

    \I__1773\ : Odrv12
    port map (
            O => \N__6954\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__1772\ : CascadeMux
    port map (
            O => \N__6951\,
            I => \N__6947\
        );

    \I__1771\ : InMux
    port map (
            O => \N__6950\,
            I => \N__6943\
        );

    \I__1770\ : InMux
    port map (
            O => \N__6947\,
            I => \N__6940\
        );

    \I__1769\ : InMux
    port map (
            O => \N__6946\,
            I => \N__6937\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__6943\,
            I => \N__6934\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__6940\,
            I => \N__6931\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__6937\,
            I => \N__6928\
        );

    \I__1765\ : Span4Mux_v
    port map (
            O => \N__6934\,
            I => \N__6925\
        );

    \I__1764\ : Span4Mux_v
    port map (
            O => \N__6931\,
            I => \N__6922\
        );

    \I__1763\ : Span4Mux_v
    port map (
            O => \N__6928\,
            I => \N__6919\
        );

    \I__1762\ : Sp12to4
    port map (
            O => \N__6925\,
            I => \N__6914\
        );

    \I__1761\ : Sp12to4
    port map (
            O => \N__6922\,
            I => \N__6914\
        );

    \I__1760\ : Sp12to4
    port map (
            O => \N__6919\,
            I => \N__6911\
        );

    \I__1759\ : Span12Mux_h
    port map (
            O => \N__6914\,
            I => \N__6908\
        );

    \I__1758\ : Span12Mux_h
    port map (
            O => \N__6911\,
            I => \N__6905\
        );

    \I__1757\ : Odrv12
    port map (
            O => \N__6908\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1756\ : Odrv12
    port map (
            O => \N__6905\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1755\ : IoInMux
    port map (
            O => \N__6900\,
            I => \N__6897\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__6897\,
            I => \N__6894\
        );

    \I__1753\ : Span4Mux_s3_v
    port map (
            O => \N__6894\,
            I => \N__6891\
        );

    \I__1752\ : Span4Mux_h
    port map (
            O => \N__6891\,
            I => \N__6888\
        );

    \I__1751\ : Span4Mux_h
    port map (
            O => \N__6888\,
            I => \N__6885\
        );

    \I__1750\ : Odrv4
    port map (
            O => \N__6885\,
            I => \un1_D_UU_AMIGA_4\
        );

    \I__1749\ : IoInMux
    port map (
            O => \N__6882\,
            I => \N__6879\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__6879\,
            I => \N__6876\
        );

    \I__1747\ : IoSpan4Mux
    port map (
            O => \N__6876\,
            I => \N__6873\
        );

    \I__1746\ : Span4Mux_s2_h
    port map (
            O => \N__6873\,
            I => \N__6870\
        );

    \I__1745\ : Sp12to4
    port map (
            O => \N__6870\,
            I => \N__6867\
        );

    \I__1744\ : Span12Mux_h
    port map (
            O => \N__6867\,
            I => \N__6864\
        );

    \I__1743\ : Odrv12
    port map (
            O => \N__6864\,
            I => \un1_D_UM_AMIGA_1\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__6861\,
            I => \N__6858\
        );

    \I__1741\ : InMux
    port map (
            O => \N__6858\,
            I => \N__6855\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__6855\,
            I => \N__6850\
        );

    \I__1739\ : InMux
    port map (
            O => \N__6854\,
            I => \N__6847\
        );

    \I__1738\ : InMux
    port map (
            O => \N__6853\,
            I => \N__6844\
        );

    \I__1737\ : Span4Mux_v
    port map (
            O => \N__6850\,
            I => \N__6841\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__6847\,
            I => \N__6836\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__6844\,
            I => \N__6836\
        );

    \I__1734\ : Span4Mux_v
    port map (
            O => \N__6841\,
            I => \N__6833\
        );

    \I__1733\ : Span4Mux_v
    port map (
            O => \N__6836\,
            I => \N__6830\
        );

    \I__1732\ : Sp12to4
    port map (
            O => \N__6833\,
            I => \N__6827\
        );

    \I__1731\ : Span4Mux_v
    port map (
            O => \N__6830\,
            I => \N__6824\
        );

    \I__1730\ : Span12Mux_h
    port map (
            O => \N__6827\,
            I => \N__6821\
        );

    \I__1729\ : Sp12to4
    port map (
            O => \N__6824\,
            I => \N__6818\
        );

    \I__1728\ : Span12Mux_v
    port map (
            O => \N__6821\,
            I => \N__6813\
        );

    \I__1727\ : Span12Mux_h
    port map (
            O => \N__6818\,
            I => \N__6813\
        );

    \I__1726\ : Odrv12
    port map (
            O => \N__6813\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1725\ : InMux
    port map (
            O => \N__6810\,
            I => \N__6807\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__6807\,
            I => \N__6804\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__6804\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__1722\ : IoInMux
    port map (
            O => \N__6801\,
            I => \N__6798\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__6798\,
            I => \N__6795\
        );

    \I__1720\ : Span4Mux_s0_h
    port map (
            O => \N__6795\,
            I => \N__6792\
        );

    \I__1719\ : Span4Mux_h
    port map (
            O => \N__6792\,
            I => \N__6789\
        );

    \I__1718\ : Sp12to4
    port map (
            O => \N__6789\,
            I => \N__6786\
        );

    \I__1717\ : Span12Mux_s11_v
    port map (
            O => \N__6786\,
            I => \N__6783\
        );

    \I__1716\ : Span12Mux_h
    port map (
            O => \N__6783\,
            I => \N__6780\
        );

    \I__1715\ : Odrv12
    port map (
            O => \N__6780\,
            I => \un1_D_UM_AMIGA_3\
        );

    \I__1714\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6773\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__6776\,
            I => \N__6770\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__6773\,
            I => \N__6767\
        );

    \I__1711\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6763\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__6767\,
            I => \N__6760\
        );

    \I__1709\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6757\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__6763\,
            I => \N__6754\
        );

    \I__1707\ : Span4Mux_v
    port map (
            O => \N__6760\,
            I => \N__6749\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__6757\,
            I => \N__6749\
        );

    \I__1705\ : Span4Mux_v
    port map (
            O => \N__6754\,
            I => \N__6746\
        );

    \I__1704\ : Span4Mux_v
    port map (
            O => \N__6749\,
            I => \N__6743\
        );

    \I__1703\ : Sp12to4
    port map (
            O => \N__6746\,
            I => \N__6740\
        );

    \I__1702\ : Sp12to4
    port map (
            O => \N__6743\,
            I => \N__6737\
        );

    \I__1701\ : Span12Mux_v
    port map (
            O => \N__6740\,
            I => \N__6734\
        );

    \I__1700\ : Span12Mux_h
    port map (
            O => \N__6737\,
            I => \N__6731\
        );

    \I__1699\ : Odrv12
    port map (
            O => \N__6734\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1698\ : Odrv12
    port map (
            O => \N__6731\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1697\ : InMux
    port map (
            O => \N__6726\,
            I => \N__6723\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__6723\,
            I => \N__6720\
        );

    \I__1695\ : Odrv12
    port map (
            O => \N__6720\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__1694\ : IoInMux
    port map (
            O => \N__6717\,
            I => \N__6714\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__6714\,
            I => \N__6711\
        );

    \I__1692\ : IoSpan4Mux
    port map (
            O => \N__6711\,
            I => \N__6708\
        );

    \I__1691\ : Span4Mux_s3_h
    port map (
            O => \N__6708\,
            I => \N__6705\
        );

    \I__1690\ : Span4Mux_h
    port map (
            O => \N__6705\,
            I => \N__6702\
        );

    \I__1689\ : Span4Mux_h
    port map (
            O => \N__6702\,
            I => \N__6699\
        );

    \I__1688\ : Span4Mux_h
    port map (
            O => \N__6699\,
            I => \N__6696\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__6696\,
            I => \un1_D_UM_AMIGA_7\
        );

    \I__1686\ : InMux
    port map (
            O => \N__6693\,
            I => \N__6690\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__6690\,
            I => \N__6687\
        );

    \I__1684\ : Odrv12
    port map (
            O => \N__6687\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__1683\ : InMux
    port map (
            O => \N__6684\,
            I => \N__6681\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__6681\,
            I => \N__6678\
        );

    \I__1681\ : Span4Mux_v
    port map (
            O => \N__6678\,
            I => \N__6675\
        );

    \I__1680\ : Span4Mux_v
    port map (
            O => \N__6675\,
            I => \N__6671\
        );

    \I__1679\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6668\
        );

    \I__1678\ : Span4Mux_v
    port map (
            O => \N__6671\,
            I => \N__6663\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__6668\,
            I => \N__6663\
        );

    \I__1676\ : Span4Mux_h
    port map (
            O => \N__6663\,
            I => \N__6659\
        );

    \I__1675\ : InMux
    port map (
            O => \N__6662\,
            I => \N__6656\
        );

    \I__1674\ : Span4Mux_v
    port map (
            O => \N__6659\,
            I => \N__6651\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__6656\,
            I => \N__6651\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__6651\,
            I => \N__6648\
        );

    \I__1671\ : Sp12to4
    port map (
            O => \N__6648\,
            I => \N__6645\
        );

    \I__1670\ : Span12Mux_h
    port map (
            O => \N__6645\,
            I => \N__6642\
        );

    \I__1669\ : Odrv12
    port map (
            O => \N__6642\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1668\ : IoInMux
    port map (
            O => \N__6639\,
            I => \N__6636\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__6636\,
            I => \N__6633\
        );

    \I__1666\ : Span4Mux_s3_v
    port map (
            O => \N__6633\,
            I => \N__6630\
        );

    \I__1665\ : Span4Mux_v
    port map (
            O => \N__6630\,
            I => \N__6627\
        );

    \I__1664\ : Sp12to4
    port map (
            O => \N__6627\,
            I => \N__6624\
        );

    \I__1663\ : Span12Mux_h
    port map (
            O => \N__6624\,
            I => \N__6621\
        );

    \I__1662\ : Odrv12
    port map (
            O => \N__6621\,
            I => \un1_D_UM_AMIGA_4\
        );

    \I__1661\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6615\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__6615\,
            I => \N__6612\
        );

    \I__1659\ : Odrv12
    port map (
            O => \N__6612\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__6609\,
            I => \N__6605\
        );

    \I__1657\ : InMux
    port map (
            O => \N__6608\,
            I => \N__6602\
        );

    \I__1656\ : InMux
    port map (
            O => \N__6605\,
            I => \N__6599\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__6602\,
            I => \N__6596\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__6599\,
            I => \N__6592\
        );

    \I__1653\ : Span4Mux_v
    port map (
            O => \N__6596\,
            I => \N__6589\
        );

    \I__1652\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6586\
        );

    \I__1651\ : Span4Mux_v
    port map (
            O => \N__6592\,
            I => \N__6583\
        );

    \I__1650\ : Span4Mux_v
    port map (
            O => \N__6589\,
            I => \N__6578\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__6586\,
            I => \N__6578\
        );

    \I__1648\ : Span4Mux_v
    port map (
            O => \N__6583\,
            I => \N__6573\
        );

    \I__1647\ : Span4Mux_h
    port map (
            O => \N__6578\,
            I => \N__6573\
        );

    \I__1646\ : Span4Mux_v
    port map (
            O => \N__6573\,
            I => \N__6570\
        );

    \I__1645\ : Span4Mux_h
    port map (
            O => \N__6570\,
            I => \N__6567\
        );

    \I__1644\ : Sp12to4
    port map (
            O => \N__6567\,
            I => \N__6564\
        );

    \I__1643\ : Odrv12
    port map (
            O => \N__6564\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1642\ : IoInMux
    port map (
            O => \N__6561\,
            I => \N__6558\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__6558\,
            I => \N__6555\
        );

    \I__1640\ : IoSpan4Mux
    port map (
            O => \N__6555\,
            I => \N__6552\
        );

    \I__1639\ : IoSpan4Mux
    port map (
            O => \N__6552\,
            I => \N__6549\
        );

    \I__1638\ : Sp12to4
    port map (
            O => \N__6549\,
            I => \N__6546\
        );

    \I__1637\ : Span12Mux_s6_v
    port map (
            O => \N__6546\,
            I => \N__6543\
        );

    \I__1636\ : Odrv12
    port map (
            O => \N__6543\,
            I => \un1_D_UU_AMIGA_5\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__6540\,
            I => \N__6537\
        );

    \I__1634\ : InMux
    port map (
            O => \N__6537\,
            I => \N__6534\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__6534\,
            I => \N__6530\
        );

    \I__1632\ : InMux
    port map (
            O => \N__6533\,
            I => \N__6527\
        );

    \I__1631\ : Span4Mux_v
    port map (
            O => \N__6530\,
            I => \N__6523\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__6527\,
            I => \N__6520\
        );

    \I__1629\ : InMux
    port map (
            O => \N__6526\,
            I => \N__6517\
        );

    \I__1628\ : Span4Mux_v
    port map (
            O => \N__6523\,
            I => \N__6514\
        );

    \I__1627\ : Span4Mux_v
    port map (
            O => \N__6520\,
            I => \N__6509\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__6517\,
            I => \N__6509\
        );

    \I__1625\ : Span4Mux_v
    port map (
            O => \N__6514\,
            I => \N__6504\
        );

    \I__1624\ : Span4Mux_v
    port map (
            O => \N__6509\,
            I => \N__6504\
        );

    \I__1623\ : Sp12to4
    port map (
            O => \N__6504\,
            I => \N__6501\
        );

    \I__1622\ : Span12Mux_h
    port map (
            O => \N__6501\,
            I => \N__6498\
        );

    \I__1621\ : Odrv12
    port map (
            O => \N__6498\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__1620\ : InMux
    port map (
            O => \N__6495\,
            I => \N__6492\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__6492\,
            I => \N__6489\
        );

    \I__1618\ : Odrv12
    port map (
            O => \N__6489\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__1617\ : IoInMux
    port map (
            O => \N__6486\,
            I => \N__6483\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__6483\,
            I => \N__6480\
        );

    \I__1615\ : Span4Mux_s2_v
    port map (
            O => \N__6480\,
            I => \N__6477\
        );

    \I__1614\ : Span4Mux_h
    port map (
            O => \N__6477\,
            I => \N__6474\
        );

    \I__1613\ : Span4Mux_v
    port map (
            O => \N__6474\,
            I => \N__6471\
        );

    \I__1612\ : Sp12to4
    port map (
            O => \N__6471\,
            I => \N__6468\
        );

    \I__1611\ : Odrv12
    port map (
            O => \N__6468\,
            I => \un1_D_UU_AMIGA_3\
        );

    \I__1610\ : IoInMux
    port map (
            O => \N__6465\,
            I => \N__6462\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__6462\,
            I => \N__6459\
        );

    \I__1608\ : IoSpan4Mux
    port map (
            O => \N__6459\,
            I => \N__6456\
        );

    \I__1607\ : Span4Mux_s2_h
    port map (
            O => \N__6456\,
            I => \N__6453\
        );

    \I__1606\ : Sp12to4
    port map (
            O => \N__6453\,
            I => \N__6450\
        );

    \I__1605\ : Odrv12
    port map (
            O => \N__6450\,
            I => \un1_D_UM_AMIGA_2\
        );

    \I__1604\ : InMux
    port map (
            O => \N__6447\,
            I => \N__6442\
        );

    \I__1603\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6439\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__6445\,
            I => \N__6436\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__6442\,
            I => \N__6431\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__6439\,
            I => \N__6431\
        );

    \I__1599\ : InMux
    port map (
            O => \N__6436\,
            I => \N__6428\
        );

    \I__1598\ : Span4Mux_v
    port map (
            O => \N__6431\,
            I => \N__6425\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__6428\,
            I => \N__6422\
        );

    \I__1596\ : Sp12to4
    port map (
            O => \N__6425\,
            I => \N__6419\
        );

    \I__1595\ : Span12Mux_v
    port map (
            O => \N__6422\,
            I => \N__6416\
        );

    \I__1594\ : Span12Mux_h
    port map (
            O => \N__6419\,
            I => \N__6413\
        );

    \I__1593\ : Odrv12
    port map (
            O => \N__6416\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1592\ : Odrv12
    port map (
            O => \N__6413\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1591\ : InMux
    port map (
            O => \N__6408\,
            I => \N__6405\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__6405\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__6402\,
            I => \U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0_cascade_\
        );

    \I__1588\ : InMux
    port map (
            O => \N__6399\,
            I => \N__6395\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__6398\,
            I => \N__6389\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__6395\,
            I => \N__6382\
        );

    \I__1585\ : InMux
    port map (
            O => \N__6394\,
            I => \N__6377\
        );

    \I__1584\ : InMux
    port map (
            O => \N__6393\,
            I => \N__6377\
        );

    \I__1583\ : InMux
    port map (
            O => \N__6392\,
            I => \N__6374\
        );

    \I__1582\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6369\
        );

    \I__1581\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6369\
        );

    \I__1580\ : InMux
    port map (
            O => \N__6387\,
            I => \N__6362\
        );

    \I__1579\ : InMux
    port map (
            O => \N__6386\,
            I => \N__6362\
        );

    \I__1578\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6362\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__6382\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__6377\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__6374\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__6369\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__6362\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__6351\,
            I => \N__6347\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__6350\,
            I => \N__6343\
        );

    \I__1570\ : InMux
    port map (
            O => \N__6347\,
            I => \N__6336\
        );

    \I__1569\ : InMux
    port map (
            O => \N__6346\,
            I => \N__6336\
        );

    \I__1568\ : InMux
    port map (
            O => \N__6343\,
            I => \N__6331\
        );

    \I__1567\ : InMux
    port map (
            O => \N__6342\,
            I => \N__6331\
        );

    \I__1566\ : InMux
    port map (
            O => \N__6341\,
            I => \N__6328\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__6336\,
            I => \N__6323\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__6331\,
            I => \N__6323\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__6328\,
            I => \N__6320\
        );

    \I__1562\ : Span4Mux_v
    port map (
            O => \N__6323\,
            I => \N__6317\
        );

    \I__1561\ : Span4Mux_h
    port map (
            O => \N__6320\,
            I => \N__6314\
        );

    \I__1560\ : Sp12to4
    port map (
            O => \N__6317\,
            I => \N__6311\
        );

    \I__1559\ : Span4Mux_v
    port map (
            O => \N__6314\,
            I => \N__6308\
        );

    \I__1558\ : Span12Mux_h
    port map (
            O => \N__6311\,
            I => \N__6305\
        );

    \I__1557\ : Span4Mux_v
    port map (
            O => \N__6308\,
            I => \N__6302\
        );

    \I__1556\ : Span12Mux_v
    port map (
            O => \N__6305\,
            I => \N__6299\
        );

    \I__1555\ : Span4Mux_v
    port map (
            O => \N__6302\,
            I => \N__6296\
        );

    \I__1554\ : Odrv12
    port map (
            O => \N__6299\,
            I => \TACKn_c\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__6296\,
            I => \TACKn_c\
        );

    \I__1552\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6285\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__6290\,
            I => \N__6277\
        );

    \I__1550\ : InMux
    port map (
            O => \N__6289\,
            I => \N__6272\
        );

    \I__1549\ : InMux
    port map (
            O => \N__6288\,
            I => \N__6272\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__6285\,
            I => \N__6269\
        );

    \I__1547\ : InMux
    port map (
            O => \N__6284\,
            I => \N__6266\
        );

    \I__1546\ : InMux
    port map (
            O => \N__6283\,
            I => \N__6261\
        );

    \I__1545\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6261\
        );

    \I__1544\ : InMux
    port map (
            O => \N__6281\,
            I => \N__6254\
        );

    \I__1543\ : InMux
    port map (
            O => \N__6280\,
            I => \N__6254\
        );

    \I__1542\ : InMux
    port map (
            O => \N__6277\,
            I => \N__6254\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__6272\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__6269\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__6266\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__6261\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__6254\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1536\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6240\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__6240\,
            I => \U111_CYCLE_SM.LW_CYCLE_0\
        );

    \I__1534\ : InMux
    port map (
            O => \N__6237\,
            I => \N__6234\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__6234\,
            I => \N__6221\
        );

    \I__1532\ : ClkMux
    port map (
            O => \N__6233\,
            I => \N__6198\
        );

    \I__1531\ : ClkMux
    port map (
            O => \N__6232\,
            I => \N__6198\
        );

    \I__1530\ : ClkMux
    port map (
            O => \N__6231\,
            I => \N__6198\
        );

    \I__1529\ : ClkMux
    port map (
            O => \N__6230\,
            I => \N__6198\
        );

    \I__1528\ : ClkMux
    port map (
            O => \N__6229\,
            I => \N__6198\
        );

    \I__1527\ : ClkMux
    port map (
            O => \N__6228\,
            I => \N__6198\
        );

    \I__1526\ : ClkMux
    port map (
            O => \N__6227\,
            I => \N__6198\
        );

    \I__1525\ : ClkMux
    port map (
            O => \N__6226\,
            I => \N__6198\
        );

    \I__1524\ : ClkMux
    port map (
            O => \N__6225\,
            I => \N__6198\
        );

    \I__1523\ : ClkMux
    port map (
            O => \N__6224\,
            I => \N__6198\
        );

    \I__1522\ : Glb2LocalMux
    port map (
            O => \N__6221\,
            I => \N__6198\
        );

    \I__1521\ : GlobalMux
    port map (
            O => \N__6198\,
            I => \CLK80\
        );

    \I__1520\ : IoInMux
    port map (
            O => \N__6195\,
            I => \N__6192\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__6192\,
            I => \N__6189\
        );

    \I__1518\ : IoSpan4Mux
    port map (
            O => \N__6189\,
            I => \N__6184\
        );

    \I__1517\ : IoInMux
    port map (
            O => \N__6188\,
            I => \N__6181\
        );

    \I__1516\ : IoInMux
    port map (
            O => \N__6187\,
            I => \N__6178\
        );

    \I__1515\ : IoSpan4Mux
    port map (
            O => \N__6184\,
            I => \N__6173\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__6181\,
            I => \N__6173\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__6178\,
            I => \N__6170\
        );

    \I__1512\ : IoSpan4Mux
    port map (
            O => \N__6173\,
            I => \N__6167\
        );

    \I__1511\ : IoSpan4Mux
    port map (
            O => \N__6170\,
            I => \N__6164\
        );

    \I__1510\ : Span4Mux_s2_v
    port map (
            O => \N__6167\,
            I => \N__6161\
        );

    \I__1509\ : Span4Mux_s2_h
    port map (
            O => \N__6164\,
            I => \N__6158\
        );

    \I__1508\ : Sp12to4
    port map (
            O => \N__6161\,
            I => \N__6155\
        );

    \I__1507\ : Sp12to4
    port map (
            O => \N__6158\,
            I => \N__6152\
        );

    \I__1506\ : Span12Mux_s9_v
    port map (
            O => \N__6155\,
            I => \N__6149\
        );

    \I__1505\ : Span12Mux_h
    port map (
            O => \N__6152\,
            I => \N__6146\
        );

    \I__1504\ : Odrv12
    port map (
            O => \N__6149\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1503\ : Odrv12
    port map (
            O => \N__6146\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__1502\ : InMux
    port map (
            O => \N__6141\,
            I => \N__6138\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__6138\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__6135\,
            I => \N__6132\
        );

    \I__1499\ : InMux
    port map (
            O => \N__6132\,
            I => \N__6129\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__6129\,
            I => \N__6124\
        );

    \I__1497\ : InMux
    port map (
            O => \N__6128\,
            I => \N__6121\
        );

    \I__1496\ : InMux
    port map (
            O => \N__6127\,
            I => \N__6118\
        );

    \I__1495\ : Span4Mux_v
    port map (
            O => \N__6124\,
            I => \N__6115\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__6121\,
            I => \N__6110\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__6118\,
            I => \N__6110\
        );

    \I__1492\ : Sp12to4
    port map (
            O => \N__6115\,
            I => \N__6107\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__6110\,
            I => \N__6104\
        );

    \I__1490\ : Span12Mux_h
    port map (
            O => \N__6107\,
            I => \N__6101\
        );

    \I__1489\ : Sp12to4
    port map (
            O => \N__6104\,
            I => \N__6098\
        );

    \I__1488\ : Span12Mux_v
    port map (
            O => \N__6101\,
            I => \N__6093\
        );

    \I__1487\ : Span12Mux_h
    port map (
            O => \N__6098\,
            I => \N__6093\
        );

    \I__1486\ : Odrv12
    port map (
            O => \N__6093\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1485\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6084\
        );

    \I__1484\ : InMux
    port map (
            O => \N__6089\,
            I => \N__6081\
        );

    \I__1483\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6076\
        );

    \I__1482\ : InMux
    port map (
            O => \N__6087\,
            I => \N__6076\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__6084\,
            I => \N__6072\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__6081\,
            I => \N__6069\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__6076\,
            I => \N__6066\
        );

    \I__1478\ : ClkMux
    port map (
            O => \N__6075\,
            I => \N__6057\
        );

    \I__1477\ : Glb2LocalMux
    port map (
            O => \N__6072\,
            I => \N__6057\
        );

    \I__1476\ : Glb2LocalMux
    port map (
            O => \N__6069\,
            I => \N__6057\
        );

    \I__1475\ : Glb2LocalMux
    port map (
            O => \N__6066\,
            I => \N__6057\
        );

    \I__1474\ : GlobalMux
    port map (
            O => \N__6057\,
            I => \CLK40\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__6054\,
            I => \U111_CYCLE_SM.N_91_cascade_\
        );

    \I__1472\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6048\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__6048\,
            I => \N__6045\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__6045\,
            I => \N__6042\
        );

    \I__1469\ : Span4Mux_v
    port map (
            O => \N__6042\,
            I => \N__6037\
        );

    \I__1468\ : InMux
    port map (
            O => \N__6041\,
            I => \N__6034\
        );

    \I__1467\ : InMux
    port map (
            O => \N__6040\,
            I => \N__6031\
        );

    \I__1466\ : Sp12to4
    port map (
            O => \N__6037\,
            I => \N__6024\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__6034\,
            I => \N__6024\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__6031\,
            I => \N__6024\
        );

    \I__1463\ : Span12Mux_h
    port map (
            O => \N__6024\,
            I => \N__6021\
        );

    \I__1462\ : Span12Mux_v
    port map (
            O => \N__6021\,
            I => \N__6018\
        );

    \I__1461\ : Odrv12
    port map (
            O => \N__6018\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__1460\ : InMux
    port map (
            O => \N__6015\,
            I => \N__6012\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__6012\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__1458\ : IoInMux
    port map (
            O => \N__6009\,
            I => \N__6006\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__6006\,
            I => \N__6003\
        );

    \I__1456\ : Span4Mux_s3_h
    port map (
            O => \N__6003\,
            I => \N__6000\
        );

    \I__1455\ : Span4Mux_h
    port map (
            O => \N__6000\,
            I => \N__5997\
        );

    \I__1454\ : Span4Mux_h
    port map (
            O => \N__5997\,
            I => \N__5994\
        );

    \I__1453\ : Span4Mux_h
    port map (
            O => \N__5994\,
            I => \N__5991\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__5991\,
            I => \un1_D_UM_AMIGA_6\
        );

    \I__1451\ : CascadeMux
    port map (
            O => \N__5988\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\
        );

    \I__1450\ : IoInMux
    port map (
            O => \N__5985\,
            I => \N__5978\
        );

    \I__1449\ : IoInMux
    port map (
            O => \N__5984\,
            I => \N__5975\
        );

    \I__1448\ : IoInMux
    port map (
            O => \N__5983\,
            I => \N__5972\
        );

    \I__1447\ : IoInMux
    port map (
            O => \N__5982\,
            I => \N__5969\
        );

    \I__1446\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5964\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__5978\,
            I => \N__5955\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__5975\,
            I => \N__5955\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__5972\,
            I => \N__5955\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__5969\,
            I => \N__5955\
        );

    \I__1441\ : IoInMux
    port map (
            O => \N__5968\,
            I => \N__5952\
        );

    \I__1440\ : IoInMux
    port map (
            O => \N__5967\,
            I => \N__5943\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__5964\,
            I => \N__5940\
        );

    \I__1438\ : IoSpan4Mux
    port map (
            O => \N__5955\,
            I => \N__5930\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__5952\,
            I => \N__5930\
        );

    \I__1436\ : IoInMux
    port map (
            O => \N__5951\,
            I => \N__5927\
        );

    \I__1435\ : IoInMux
    port map (
            O => \N__5950\,
            I => \N__5924\
        );

    \I__1434\ : IoInMux
    port map (
            O => \N__5949\,
            I => \N__5921\
        );

    \I__1433\ : IoInMux
    port map (
            O => \N__5948\,
            I => \N__5918\
        );

    \I__1432\ : IoInMux
    port map (
            O => \N__5947\,
            I => \N__5915\
        );

    \I__1431\ : IoInMux
    port map (
            O => \N__5946\,
            I => \N__5912\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__5943\,
            I => \N__5908\
        );

    \I__1429\ : Span4Mux_h
    port map (
            O => \N__5940\,
            I => \N__5905\
        );

    \I__1428\ : IoInMux
    port map (
            O => \N__5939\,
            I => \N__5901\
        );

    \I__1427\ : IoInMux
    port map (
            O => \N__5938\,
            I => \N__5898\
        );

    \I__1426\ : IoInMux
    port map (
            O => \N__5937\,
            I => \N__5895\
        );

    \I__1425\ : IoInMux
    port map (
            O => \N__5936\,
            I => \N__5892\
        );

    \I__1424\ : IoInMux
    port map (
            O => \N__5935\,
            I => \N__5889\
        );

    \I__1423\ : IoSpan4Mux
    port map (
            O => \N__5930\,
            I => \N__5870\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__5927\,
            I => \N__5870\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__5924\,
            I => \N__5870\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__5921\,
            I => \N__5870\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__5918\,
            I => \N__5870\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__5915\,
            I => \N__5870\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__5912\,
            I => \N__5870\
        );

    \I__1416\ : IoInMux
    port map (
            O => \N__5911\,
            I => \N__5867\
        );

    \I__1415\ : Span4Mux_s3_v
    port map (
            O => \N__5908\,
            I => \N__5863\
        );

    \I__1414\ : Span4Mux_v
    port map (
            O => \N__5905\,
            I => \N__5860\
        );

    \I__1413\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5857\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__5901\,
            I => \N__5846\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__5898\,
            I => \N__5846\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__5895\,
            I => \N__5846\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__5892\,
            I => \N__5846\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__5889\,
            I => \N__5846\
        );

    \I__1407\ : IoInMux
    port map (
            O => \N__5888\,
            I => \N__5843\
        );

    \I__1406\ : IoInMux
    port map (
            O => \N__5887\,
            I => \N__5840\
        );

    \I__1405\ : IoInMux
    port map (
            O => \N__5886\,
            I => \N__5837\
        );

    \I__1404\ : IoInMux
    port map (
            O => \N__5885\,
            I => \N__5834\
        );

    \I__1403\ : IoSpan4Mux
    port map (
            O => \N__5870\,
            I => \N__5825\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__5867\,
            I => \N__5825\
        );

    \I__1401\ : IoInMux
    port map (
            O => \N__5866\,
            I => \N__5822\
        );

    \I__1400\ : Span4Mux_v
    port map (
            O => \N__5863\,
            I => \N__5817\
        );

    \I__1399\ : Span4Mux_h
    port map (
            O => \N__5860\,
            I => \N__5812\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__5857\,
            I => \N__5812\
        );

    \I__1397\ : IoSpan4Mux
    port map (
            O => \N__5846\,
            I => \N__5801\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__5843\,
            I => \N__5801\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__5840\,
            I => \N__5801\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__5837\,
            I => \N__5801\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__5834\,
            I => \N__5801\
        );

    \I__1392\ : IoInMux
    port map (
            O => \N__5833\,
            I => \N__5798\
        );

    \I__1391\ : IoInMux
    port map (
            O => \N__5832\,
            I => \N__5795\
        );

    \I__1390\ : IoInMux
    port map (
            O => \N__5831\,
            I => \N__5792\
        );

    \I__1389\ : IoInMux
    port map (
            O => \N__5830\,
            I => \N__5789\
        );

    \I__1388\ : IoSpan4Mux
    port map (
            O => \N__5825\,
            I => \N__5784\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__5822\,
            I => \N__5784\
        );

    \I__1386\ : IoInMux
    port map (
            O => \N__5821\,
            I => \N__5781\
        );

    \I__1385\ : IoInMux
    port map (
            O => \N__5820\,
            I => \N__5778\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__5817\,
            I => \N__5774\
        );

    \I__1383\ : Span4Mux_v
    port map (
            O => \N__5812\,
            I => \N__5771\
        );

    \I__1382\ : IoSpan4Mux
    port map (
            O => \N__5801\,
            I => \N__5760\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__5798\,
            I => \N__5760\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__5795\,
            I => \N__5760\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__5792\,
            I => \N__5760\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__5789\,
            I => \N__5760\
        );

    \I__1377\ : IoSpan4Mux
    port map (
            O => \N__5784\,
            I => \N__5753\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__5781\,
            I => \N__5753\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__5778\,
            I => \N__5753\
        );

    \I__1374\ : IoInMux
    port map (
            O => \N__5777\,
            I => \N__5750\
        );

    \I__1373\ : Sp12to4
    port map (
            O => \N__5774\,
            I => \N__5745\
        );

    \I__1372\ : Sp12to4
    port map (
            O => \N__5771\,
            I => \N__5741\
        );

    \I__1371\ : IoSpan4Mux
    port map (
            O => \N__5760\,
            I => \N__5738\
        );

    \I__1370\ : IoSpan4Mux
    port map (
            O => \N__5753\,
            I => \N__5733\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__5750\,
            I => \N__5733\
        );

    \I__1368\ : IoInMux
    port map (
            O => \N__5749\,
            I => \N__5730\
        );

    \I__1367\ : IoInMux
    port map (
            O => \N__5748\,
            I => \N__5727\
        );

    \I__1366\ : Span12Mux_h
    port map (
            O => \N__5745\,
            I => \N__5724\
        );

    \I__1365\ : IoInMux
    port map (
            O => \N__5744\,
            I => \N__5721\
        );

    \I__1364\ : Span12Mux_h
    port map (
            O => \N__5741\,
            I => \N__5718\
        );

    \I__1363\ : IoSpan4Mux
    port map (
            O => \N__5738\,
            I => \N__5713\
        );

    \I__1362\ : IoSpan4Mux
    port map (
            O => \N__5733\,
            I => \N__5713\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__5730\,
            I => \N__5710\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__5727\,
            I => \N__5707\
        );

    \I__1359\ : Span12Mux_h
    port map (
            O => \N__5724\,
            I => \N__5702\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__5721\,
            I => \N__5702\
        );

    \I__1357\ : Odrv12
    port map (
            O => \N__5718\,
            I => \RnW_c\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__5713\,
            I => \RnW_c\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__5710\,
            I => \RnW_c\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__5707\,
            I => \RnW_c\
        );

    \I__1353\ : Odrv12
    port map (
            O => \N__5702\,
            I => \RnW_c\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__5691\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_\
        );

    \I__1351\ : InMux
    port map (
            O => \N__5688\,
            I => \N__5685\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__5685\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\
        );

    \I__1349\ : CascadeMux
    port map (
            O => \N__5682\,
            I => \N__5675\
        );

    \I__1348\ : InMux
    port map (
            O => \N__5681\,
            I => \N__5672\
        );

    \I__1347\ : InMux
    port map (
            O => \N__5680\,
            I => \N__5669\
        );

    \I__1346\ : InMux
    port map (
            O => \N__5679\,
            I => \N__5666\
        );

    \I__1345\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5663\
        );

    \I__1344\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5660\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__5672\,
            I => \N__5657\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__5669\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__5666\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__5663\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__5660\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__5657\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__1337\ : InMux
    port map (
            O => \N__5646\,
            I => \N__5640\
        );

    \I__1336\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5637\
        );

    \I__1335\ : CascadeMux
    port map (
            O => \N__5644\,
            I => \N__5632\
        );

    \I__1334\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5628\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__5640\,
            I => \N__5623\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__5637\,
            I => \N__5623\
        );

    \I__1331\ : InMux
    port map (
            O => \N__5636\,
            I => \N__5618\
        );

    \I__1330\ : InMux
    port map (
            O => \N__5635\,
            I => \N__5618\
        );

    \I__1329\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5613\
        );

    \I__1328\ : InMux
    port map (
            O => \N__5631\,
            I => \N__5613\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__5628\,
            I => \N__5610\
        );

    \I__1326\ : Span4Mux_v
    port map (
            O => \N__5623\,
            I => \N__5602\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__5618\,
            I => \N__5602\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__5613\,
            I => \N__5602\
        );

    \I__1323\ : Span4Mux_v
    port map (
            O => \N__5610\,
            I => \N__5598\
        );

    \I__1322\ : InMux
    port map (
            O => \N__5609\,
            I => \N__5595\
        );

    \I__1321\ : Span4Mux_v
    port map (
            O => \N__5602\,
            I => \N__5592\
        );

    \I__1320\ : InMux
    port map (
            O => \N__5601\,
            I => \N__5589\
        );

    \I__1319\ : Sp12to4
    port map (
            O => \N__5598\,
            I => \N__5584\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__5595\,
            I => \N__5584\
        );

    \I__1317\ : Span4Mux_h
    port map (
            O => \N__5592\,
            I => \N__5581\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__5589\,
            I => \N__5578\
        );

    \I__1315\ : Span12Mux_h
    port map (
            O => \N__5584\,
            I => \N__5575\
        );

    \I__1314\ : Sp12to4
    port map (
            O => \N__5581\,
            I => \N__5572\
        );

    \I__1313\ : Span4Mux_v
    port map (
            O => \N__5578\,
            I => \N__5569\
        );

    \I__1312\ : Span12Mux_v
    port map (
            O => \N__5575\,
            I => \N__5566\
        );

    \I__1311\ : Span12Mux_v
    port map (
            O => \N__5572\,
            I => \N__5561\
        );

    \I__1310\ : Sp12to4
    port map (
            O => \N__5569\,
            I => \N__5561\
        );

    \I__1309\ : Odrv12
    port map (
            O => \N__5566\,
            I => \RESETn_c\
        );

    \I__1308\ : Odrv12
    port map (
            O => \N__5561\,
            I => \RESETn_c\
        );

    \I__1307\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5553\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__5553\,
            I => \N__5550\
        );

    \I__1305\ : Span4Mux_v
    port map (
            O => \N__5550\,
            I => \N__5547\
        );

    \I__1304\ : Odrv4
    port map (
            O => \N__5547\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__5544\,
            I => \N__5541\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5537\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5534\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__5537\,
            I => \N__5531\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__5534\,
            I => \N__5528\
        );

    \I__1298\ : Span4Mux_v
    port map (
            O => \N__5531\,
            I => \N__5524\
        );

    \I__1297\ : Span4Mux_v
    port map (
            O => \N__5528\,
            I => \N__5521\
        );

    \I__1296\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5518\
        );

    \I__1295\ : Span4Mux_v
    port map (
            O => \N__5524\,
            I => \N__5515\
        );

    \I__1294\ : Span4Mux_v
    port map (
            O => \N__5521\,
            I => \N__5510\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__5518\,
            I => \N__5510\
        );

    \I__1292\ : Span4Mux_v
    port map (
            O => \N__5515\,
            I => \N__5507\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__5510\,
            I => \N__5504\
        );

    \I__1290\ : Sp12to4
    port map (
            O => \N__5507\,
            I => \N__5499\
        );

    \I__1289\ : Sp12to4
    port map (
            O => \N__5504\,
            I => \N__5499\
        );

    \I__1288\ : Span12Mux_h
    port map (
            O => \N__5499\,
            I => \N__5496\
        );

    \I__1287\ : Odrv12
    port map (
            O => \N__5496\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__1286\ : IoInMux
    port map (
            O => \N__5493\,
            I => \N__5490\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__5490\,
            I => \N__5487\
        );

    \I__1284\ : Span12Mux_s11_v
    port map (
            O => \N__5487\,
            I => \N__5484\
        );

    \I__1283\ : Span12Mux_h
    port map (
            O => \N__5484\,
            I => \N__5481\
        );

    \I__1282\ : Odrv12
    port map (
            O => \N__5481\,
            I => \un1_D_UU_AMIGA_2\
        );

    \I__1281\ : IoInMux
    port map (
            O => \N__5478\,
            I => \N__5473\
        );

    \I__1280\ : IoInMux
    port map (
            O => \N__5477\,
            I => \N__5470\
        );

    \I__1279\ : IoInMux
    port map (
            O => \N__5476\,
            I => \N__5467\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5473\,
            I => \N__5464\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5470\,
            I => \N__5461\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__5467\,
            I => \N__5458\
        );

    \I__1275\ : Span12Mux_s4_v
    port map (
            O => \N__5464\,
            I => \N__5455\
        );

    \I__1274\ : Span12Mux_s9_h
    port map (
            O => \N__5461\,
            I => \N__5450\
        );

    \I__1273\ : Span12Mux_s10_h
    port map (
            O => \N__5458\,
            I => \N__5450\
        );

    \I__1272\ : Odrv12
    port map (
            O => \N__5455\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__1271\ : Odrv12
    port map (
            O => \N__5450\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__5445\,
            I => \N__5441\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5438\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5435\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__5438\,
            I => \U111_CYCLE_SM.TA_ENZ0\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__5435\,
            I => \U111_CYCLE_SM.TA_ENZ0\
        );

    \I__1265\ : IoInMux
    port map (
            O => \N__5430\,
            I => \N__5426\
        );

    \I__1264\ : IoInMux
    port map (
            O => \N__5429\,
            I => \N__5423\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5426\,
            I => \N__5420\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__5423\,
            I => \N__5417\
        );

    \I__1261\ : Span4Mux_s3_v
    port map (
            O => \N__5420\,
            I => \N__5414\
        );

    \I__1260\ : Span4Mux_s2_v
    port map (
            O => \N__5417\,
            I => \N__5411\
        );

    \I__1259\ : Sp12to4
    port map (
            O => \N__5414\,
            I => \N__5408\
        );

    \I__1258\ : Span4Mux_h
    port map (
            O => \N__5411\,
            I => \N__5405\
        );

    \I__1257\ : Span12Mux_s11_h
    port map (
            O => \N__5408\,
            I => \N__5402\
        );

    \I__1256\ : Span4Mux_v
    port map (
            O => \N__5405\,
            I => \N__5399\
        );

    \I__1255\ : Span12Mux_v
    port map (
            O => \N__5402\,
            I => \N__5396\
        );

    \I__1254\ : Sp12to4
    port map (
            O => \N__5399\,
            I => \N__5393\
        );

    \I__1253\ : Odrv12
    port map (
            O => \N__5396\,
            I => \U111_CYCLE_SM_TAn_0_i\
        );

    \I__1252\ : Odrv12
    port map (
            O => \N__5393\,
            I => \U111_CYCLE_SM_TAn_0_i\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5388\,
            I => \N__5381\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5387\,
            I => \N__5381\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5375\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5381\,
            I => \N__5369\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5363\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5379\,
            I => \N__5360\
        );

    \I__1245\ : InMux
    port map (
            O => \N__5378\,
            I => \N__5357\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5375\,
            I => \N__5353\
        );

    \I__1243\ : InMux
    port map (
            O => \N__5374\,
            I => \N__5349\
        );

    \I__1242\ : InMux
    port map (
            O => \N__5373\,
            I => \N__5345\
        );

    \I__1241\ : InMux
    port map (
            O => \N__5372\,
            I => \N__5334\
        );

    \I__1240\ : Span4Mux_h
    port map (
            O => \N__5369\,
            I => \N__5331\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5368\,
            I => \N__5328\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5367\,
            I => \N__5323\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5323\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__5363\,
            I => \N__5318\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__5360\,
            I => \N__5313\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5357\,
            I => \N__5313\
        );

    \I__1233\ : InMux
    port map (
            O => \N__5356\,
            I => \N__5310\
        );

    \I__1232\ : Span4Mux_h
    port map (
            O => \N__5353\,
            I => \N__5304\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5352\,
            I => \N__5301\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5349\,
            I => \N__5298\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5295\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5345\,
            I => \N__5292\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5344\,
            I => \N__5289\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5343\,
            I => \N__5286\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5281\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5281\
        );

    \I__1223\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5276\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5276\
        );

    \I__1221\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5272\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5337\,
            I => \N__5269\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5334\,
            I => \N__5265\
        );

    \I__1218\ : Span4Mux_v
    port map (
            O => \N__5331\,
            I => \N__5262\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__5328\,
            I => \N__5259\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__5323\,
            I => \N__5256\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5322\,
            I => \N__5251\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5251\
        );

    \I__1213\ : Span4Mux_h
    port map (
            O => \N__5318\,
            I => \N__5246\
        );

    \I__1212\ : Span4Mux_v
    port map (
            O => \N__5313\,
            I => \N__5246\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5310\,
            I => \N__5243\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5240\
        );

    \I__1209\ : InMux
    port map (
            O => \N__5308\,
            I => \N__5237\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5307\,
            I => \N__5234\
        );

    \I__1207\ : Span4Mux_v
    port map (
            O => \N__5304\,
            I => \N__5229\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__5301\,
            I => \N__5229\
        );

    \I__1205\ : Span4Mux_v
    port map (
            O => \N__5298\,
            I => \N__5223\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5295\,
            I => \N__5223\
        );

    \I__1203\ : Span4Mux_v
    port map (
            O => \N__5292\,
            I => \N__5216\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5289\,
            I => \N__5216\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__5286\,
            I => \N__5216\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5281\,
            I => \N__5211\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5276\,
            I => \N__5211\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5208\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5272\,
            I => \N__5205\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5269\,
            I => \N__5202\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5199\
        );

    \I__1194\ : Span4Mux_h
    port map (
            O => \N__5265\,
            I => \N__5195\
        );

    \I__1193\ : Span4Mux_v
    port map (
            O => \N__5262\,
            I => \N__5190\
        );

    \I__1192\ : Span4Mux_h
    port map (
            O => \N__5259\,
            I => \N__5190\
        );

    \I__1191\ : Span4Mux_v
    port map (
            O => \N__5256\,
            I => \N__5185\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__5251\,
            I => \N__5185\
        );

    \I__1189\ : Span4Mux_v
    port map (
            O => \N__5246\,
            I => \N__5174\
        );

    \I__1188\ : Span4Mux_h
    port map (
            O => \N__5243\,
            I => \N__5174\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5240\,
            I => \N__5174\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5237\,
            I => \N__5174\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__5234\,
            I => \N__5174\
        );

    \I__1184\ : Span4Mux_v
    port map (
            O => \N__5229\,
            I => \N__5171\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5228\,
            I => \N__5168\
        );

    \I__1182\ : Span4Mux_h
    port map (
            O => \N__5223\,
            I => \N__5165\
        );

    \I__1181\ : Span4Mux_h
    port map (
            O => \N__5216\,
            I => \N__5158\
        );

    \I__1180\ : Span4Mux_v
    port map (
            O => \N__5211\,
            I => \N__5158\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5208\,
            I => \N__5158\
        );

    \I__1178\ : Span4Mux_v
    port map (
            O => \N__5205\,
            I => \N__5151\
        );

    \I__1177\ : Span4Mux_h
    port map (
            O => \N__5202\,
            I => \N__5151\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__5199\,
            I => \N__5151\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5198\,
            I => \N__5148\
        );

    \I__1174\ : Sp12to4
    port map (
            O => \N__5195\,
            I => \N__5145\
        );

    \I__1173\ : Span4Mux_h
    port map (
            O => \N__5190\,
            I => \N__5140\
        );

    \I__1172\ : Span4Mux_v
    port map (
            O => \N__5185\,
            I => \N__5140\
        );

    \I__1171\ : Span4Mux_v
    port map (
            O => \N__5174\,
            I => \N__5137\
        );

    \I__1170\ : Sp12to4
    port map (
            O => \N__5171\,
            I => \N__5132\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__5168\,
            I => \N__5132\
        );

    \I__1168\ : Span4Mux_v
    port map (
            O => \N__5165\,
            I => \N__5123\
        );

    \I__1167\ : Span4Mux_v
    port map (
            O => \N__5158\,
            I => \N__5123\
        );

    \I__1166\ : Span4Mux_h
    port map (
            O => \N__5151\,
            I => \N__5123\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5148\,
            I => \N__5123\
        );

    \I__1164\ : Odrv12
    port map (
            O => \N__5145\,
            I => \U111_CYCLE_SM.un1_LW_TRANS_1_0\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__5140\,
            I => \U111_CYCLE_SM.un1_LW_TRANS_1_0\
        );

    \I__1162\ : Odrv4
    port map (
            O => \N__5137\,
            I => \U111_CYCLE_SM.un1_LW_TRANS_1_0\
        );

    \I__1161\ : Odrv12
    port map (
            O => \N__5132\,
            I => \U111_CYCLE_SM.un1_LW_TRANS_1_0\
        );

    \I__1160\ : Odrv4
    port map (
            O => \N__5123\,
            I => \U111_CYCLE_SM.un1_LW_TRANS_1_0\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5112\,
            I => \N__5106\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5111\,
            I => \N__5106\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5106\,
            I => \N__5103\
        );

    \I__1156\ : Span12Mux_h
    port map (
            O => \N__5103\,
            I => \N__5100\
        );

    \I__1155\ : Span12Mux_v
    port map (
            O => \N__5100\,
            I => \N__5097\
        );

    \I__1154\ : Odrv12
    port map (
            O => \N__5097\,
            I => \PORTSIZE_c\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5094\,
            I => \N__5088\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5093\,
            I => \N__5088\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5088\,
            I => \N__5085\
        );

    \I__1150\ : Span12Mux_h
    port map (
            O => \N__5085\,
            I => \N__5082\
        );

    \I__1149\ : Span12Mux_v
    port map (
            O => \N__5082\,
            I => \N__5079\
        );

    \I__1148\ : Odrv12
    port map (
            O => \N__5079\,
            I => \SIZ_c_1\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__5076\,
            I => \N__5073\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5073\,
            I => \N__5067\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5072\,
            I => \N__5067\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__5067\,
            I => \N__5064\
        );

    \I__1143\ : Span12Mux_h
    port map (
            O => \N__5064\,
            I => \N__5061\
        );

    \I__1142\ : Span12Mux_v
    port map (
            O => \N__5061\,
            I => \N__5058\
        );

    \I__1141\ : Odrv12
    port map (
            O => \N__5058\,
            I => \SIZ_c_0\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5052\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5052\,
            I => \N__5049\
        );

    \I__1138\ : Span4Mux_h
    port map (
            O => \N__5049\,
            I => \N__5044\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5048\,
            I => \N__5039\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5039\
        );

    \I__1135\ : Sp12to4
    port map (
            O => \N__5044\,
            I => \N__5036\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__5039\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__1133\ : Odrv12
    port map (
            O => \N__5036\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__5031\,
            I => \U111_CYCLE_SM.un3_LW_CYCLE_START_cascade_\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5028\,
            I => \N__5025\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__5025\,
            I => \N__5022\
        );

    \I__1129\ : Span4Mux_h
    port map (
            O => \N__5022\,
            I => \N__5019\
        );

    \I__1128\ : Sp12to4
    port map (
            O => \N__5019\,
            I => \N__5016\
        );

    \I__1127\ : Span12Mux_v
    port map (
            O => \N__5016\,
            I => \N__5013\
        );

    \I__1126\ : Odrv12
    port map (
            O => \N__5013\,
            I => \TS_CPUn_c\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5010\,
            I => \N__5007\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5007\,
            I => \U111_CYCLE_SM.TS_EN_5\
        );

    \I__1123\ : InMux
    port map (
            O => \N__5004\,
            I => \N__5001\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__5001\,
            I => \U111_CYCLE_SM.N_69_0\
        );

    \I__1121\ : IoInMux
    port map (
            O => \N__4998\,
            I => \N__4995\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__4995\,
            I => \N__4991\
        );

    \I__1119\ : IoInMux
    port map (
            O => \N__4994\,
            I => \N__4986\
        );

    \I__1118\ : IoSpan4Mux
    port map (
            O => \N__4991\,
            I => \N__4983\
        );

    \I__1117\ : IoInMux
    port map (
            O => \N__4990\,
            I => \N__4978\
        );

    \I__1116\ : IoInMux
    port map (
            O => \N__4989\,
            I => \N__4978\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__4986\,
            I => \N__4975\
        );

    \I__1114\ : IoSpan4Mux
    port map (
            O => \N__4983\,
            I => \N__4972\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__4978\,
            I => \N__4969\
        );

    \I__1112\ : Span4Mux_s3_h
    port map (
            O => \N__4975\,
            I => \N__4966\
        );

    \I__1111\ : IoSpan4Mux
    port map (
            O => \N__4972\,
            I => \N__4961\
        );

    \I__1110\ : IoSpan4Mux
    port map (
            O => \N__4969\,
            I => \N__4961\
        );

    \I__1109\ : Span4Mux_v
    port map (
            O => \N__4966\,
            I => \N__4958\
        );

    \I__1108\ : Span4Mux_s2_v
    port map (
            O => \N__4961\,
            I => \N__4955\
        );

    \I__1107\ : Sp12to4
    port map (
            O => \N__4958\,
            I => \N__4952\
        );

    \I__1106\ : Span4Mux_v
    port map (
            O => \N__4955\,
            I => \N__4949\
        );

    \I__1105\ : Span12Mux_h
    port map (
            O => \N__4952\,
            I => \N__4946\
        );

    \I__1104\ : Span4Mux_v
    port map (
            O => \N__4949\,
            I => \N__4943\
        );

    \I__1103\ : Odrv12
    port map (
            O => \N__4946\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__4943\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1101\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4935\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__4935\,
            I => \N__4932\
        );

    \I__1099\ : Span4Mux_v
    port map (
            O => \N__4932\,
            I => \N__4929\
        );

    \I__1098\ : Span4Mux_h
    port map (
            O => \N__4929\,
            I => \N__4926\
        );

    \I__1097\ : Sp12to4
    port map (
            O => \N__4926\,
            I => \N__4923\
        );

    \I__1096\ : Odrv12
    port map (
            O => \N__4923\,
            I => \D_LM_AMIGA_in_7\
        );

    \I__1095\ : IoInMux
    port map (
            O => \N__4920\,
            I => \N__4917\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__4917\,
            I => \N__4914\
        );

    \I__1093\ : IoSpan4Mux
    port map (
            O => \N__4914\,
            I => \N__4911\
        );

    \I__1092\ : Span4Mux_s2_h
    port map (
            O => \N__4911\,
            I => \N__4908\
        );

    \I__1091\ : Span4Mux_h
    port map (
            O => \N__4908\,
            I => \N__4905\
        );

    \I__1090\ : Sp12to4
    port map (
            O => \N__4905\,
            I => \N__4902\
        );

    \I__1089\ : Odrv12
    port map (
            O => \N__4902\,
            I => \un1_D_LM_AMIGA_7\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__4899\,
            I => \N__4896\
        );

    \I__1087\ : InMux
    port map (
            O => \N__4896\,
            I => \N__4893\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__4893\,
            I => \N__4890\
        );

    \I__1085\ : Span4Mux_v
    port map (
            O => \N__4890\,
            I => \N__4887\
        );

    \I__1084\ : Span4Mux_v
    port map (
            O => \N__4887\,
            I => \N__4884\
        );

    \I__1083\ : Sp12to4
    port map (
            O => \N__4884\,
            I => \N__4881\
        );

    \I__1082\ : Span12Mux_h
    port map (
            O => \N__4881\,
            I => \N__4878\
        );

    \I__1081\ : Odrv12
    port map (
            O => \N__4878\,
            I => \D_UM_040_in_7\
        );

    \I__1080\ : IoInMux
    port map (
            O => \N__4875\,
            I => \N__4872\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__4872\,
            I => \N__4869\
        );

    \I__1078\ : IoSpan4Mux
    port map (
            O => \N__4869\,
            I => \N__4865\
        );

    \I__1077\ : InMux
    port map (
            O => \N__4868\,
            I => \N__4862\
        );

    \I__1076\ : Span4Mux_s3_h
    port map (
            O => \N__4865\,
            I => \N__4859\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__4862\,
            I => \N__4856\
        );

    \I__1074\ : Sp12to4
    port map (
            O => \N__4859\,
            I => \N__4853\
        );

    \I__1073\ : Sp12to4
    port map (
            O => \N__4856\,
            I => \N__4850\
        );

    \I__1072\ : Span12Mux_v
    port map (
            O => \N__4853\,
            I => \N__4847\
        );

    \I__1071\ : Span12Mux_v
    port map (
            O => \N__4850\,
            I => \N__4844\
        );

    \I__1070\ : Span12Mux_h
    port map (
            O => \N__4847\,
            I => \N__4841\
        );

    \I__1069\ : Span12Mux_h
    port map (
            O => \N__4844\,
            I => \N__4838\
        );

    \I__1068\ : Span12Mux_h
    port map (
            O => \N__4841\,
            I => \N__4833\
        );

    \I__1067\ : Span12Mux_v
    port map (
            O => \N__4838\,
            I => \N__4833\
        );

    \I__1066\ : Odrv12
    port map (
            O => \N__4833\,
            I => \D_LL_040_in_7\
        );

    \I__1065\ : IoInMux
    port map (
            O => \N__4830\,
            I => \N__4827\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__4827\,
            I => \N__4824\
        );

    \I__1063\ : Span12Mux_s2_h
    port map (
            O => \N__4824\,
            I => \N__4821\
        );

    \I__1062\ : Span12Mux_h
    port map (
            O => \N__4821\,
            I => \N__4818\
        );

    \I__1061\ : Odrv12
    port map (
            O => \N__4818\,
            I => \un1_D_UM_040_7\
        );

    \I__1060\ : InMux
    port map (
            O => \N__4815\,
            I => \N__4812\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__4812\,
            I => \N__4809\
        );

    \I__1058\ : Sp12to4
    port map (
            O => \N__4809\,
            I => \N__4806\
        );

    \I__1057\ : Span12Mux_v
    port map (
            O => \N__4806\,
            I => \N__4803\
        );

    \I__1056\ : Span12Mux_h
    port map (
            O => \N__4803\,
            I => \N__4800\
        );

    \I__1055\ : Odrv12
    port map (
            O => \N__4800\,
            I => \D_UU_040_in_0\
        );

    \I__1054\ : IoInMux
    port map (
            O => \N__4797\,
            I => \N__4793\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__4796\,
            I => \N__4790\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__4793\,
            I => \N__4787\
        );

    \I__1051\ : InMux
    port map (
            O => \N__4790\,
            I => \N__4784\
        );

    \I__1050\ : IoSpan4Mux
    port map (
            O => \N__4787\,
            I => \N__4781\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__4784\,
            I => \N__4778\
        );

    \I__1048\ : IoSpan4Mux
    port map (
            O => \N__4781\,
            I => \N__4775\
        );

    \I__1047\ : Span4Mux_h
    port map (
            O => \N__4778\,
            I => \N__4772\
        );

    \I__1046\ : Span4Mux_s2_h
    port map (
            O => \N__4775\,
            I => \N__4769\
        );

    \I__1045\ : Sp12to4
    port map (
            O => \N__4772\,
            I => \N__4766\
        );

    \I__1044\ : Sp12to4
    port map (
            O => \N__4769\,
            I => \N__4763\
        );

    \I__1043\ : Span12Mux_v
    port map (
            O => \N__4766\,
            I => \N__4760\
        );

    \I__1042\ : Span12Mux_h
    port map (
            O => \N__4763\,
            I => \N__4757\
        );

    \I__1041\ : Span12Mux_v
    port map (
            O => \N__4760\,
            I => \N__4754\
        );

    \I__1040\ : Span12Mux_h
    port map (
            O => \N__4757\,
            I => \N__4751\
        );

    \I__1039\ : Span12Mux_h
    port map (
            O => \N__4754\,
            I => \N__4748\
        );

    \I__1038\ : Odrv12
    port map (
            O => \N__4751\,
            I => \D_LM_040_in_0\
        );

    \I__1037\ : Odrv12
    port map (
            O => \N__4748\,
            I => \D_LM_040_in_0\
        );

    \I__1036\ : IoInMux
    port map (
            O => \N__4743\,
            I => \N__4740\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__4740\,
            I => \N__4737\
        );

    \I__1034\ : Span4Mux_s3_v
    port map (
            O => \N__4737\,
            I => \N__4734\
        );

    \I__1033\ : Sp12to4
    port map (
            O => \N__4734\,
            I => \N__4731\
        );

    \I__1032\ : Span12Mux_h
    port map (
            O => \N__4731\,
            I => \N__4728\
        );

    \I__1031\ : Odrv12
    port map (
            O => \N__4728\,
            I => \un1_D_UU_040_0\
        );

    \I__1030\ : IoInMux
    port map (
            O => \N__4725\,
            I => \N__4721\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__4724\,
            I => \N__4718\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4721\,
            I => \N__4715\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4712\
        );

    \I__1026\ : IoSpan4Mux
    port map (
            O => \N__4715\,
            I => \N__4709\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__4712\,
            I => \N__4706\
        );

    \I__1024\ : Span4Mux_s3_h
    port map (
            O => \N__4709\,
            I => \N__4703\
        );

    \I__1023\ : Sp12to4
    port map (
            O => \N__4706\,
            I => \N__4700\
        );

    \I__1022\ : Sp12to4
    port map (
            O => \N__4703\,
            I => \N__4697\
        );

    \I__1021\ : Span12Mux_v
    port map (
            O => \N__4700\,
            I => \N__4694\
        );

    \I__1020\ : Span12Mux_v
    port map (
            O => \N__4697\,
            I => \N__4691\
        );

    \I__1019\ : Span12Mux_v
    port map (
            O => \N__4694\,
            I => \N__4686\
        );

    \I__1018\ : Span12Mux_h
    port map (
            O => \N__4691\,
            I => \N__4686\
        );

    \I__1017\ : Span12Mux_h
    port map (
            O => \N__4686\,
            I => \N__4683\
        );

    \I__1016\ : Odrv12
    port map (
            O => \N__4683\,
            I => \D_LL_040_in_5\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4680\,
            I => \N__4677\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__4677\,
            I => \N__4674\
        );

    \I__1013\ : Span4Mux_v
    port map (
            O => \N__4674\,
            I => \N__4671\
        );

    \I__1012\ : Span4Mux_h
    port map (
            O => \N__4671\,
            I => \N__4668\
        );

    \I__1011\ : Sp12to4
    port map (
            O => \N__4668\,
            I => \N__4665\
        );

    \I__1010\ : Span12Mux_h
    port map (
            O => \N__4665\,
            I => \N__4662\
        );

    \I__1009\ : Odrv12
    port map (
            O => \N__4662\,
            I => \D_UM_040_in_5\
        );

    \I__1008\ : IoInMux
    port map (
            O => \N__4659\,
            I => \N__4656\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4656\,
            I => \N__4653\
        );

    \I__1006\ : IoSpan4Mux
    port map (
            O => \N__4653\,
            I => \N__4650\
        );

    \I__1005\ : IoSpan4Mux
    port map (
            O => \N__4650\,
            I => \N__4647\
        );

    \I__1004\ : Span4Mux_s2_v
    port map (
            O => \N__4647\,
            I => \N__4644\
        );

    \I__1003\ : Span4Mux_v
    port map (
            O => \N__4644\,
            I => \N__4641\
        );

    \I__1002\ : Odrv4
    port map (
            O => \N__4641\,
            I => \un1_D_UM_040_5\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4638\,
            I => \N__4635\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4635\,
            I => \N__4632\
        );

    \I__999\ : Span4Mux_v
    port map (
            O => \N__4632\,
            I => \N__4629\
        );

    \I__998\ : Span4Mux_h
    port map (
            O => \N__4629\,
            I => \N__4626\
        );

    \I__997\ : Sp12to4
    port map (
            O => \N__4626\,
            I => \N__4623\
        );

    \I__996\ : Span12Mux_h
    port map (
            O => \N__4623\,
            I => \N__4620\
        );

    \I__995\ : Odrv12
    port map (
            O => \N__4620\,
            I => \D_UU_040_in_5\
        );

    \I__994\ : IoInMux
    port map (
            O => \N__4617\,
            I => \N__4614\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4614\,
            I => \N__4610\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__4613\,
            I => \N__4607\
        );

    \I__991\ : IoSpan4Mux
    port map (
            O => \N__4610\,
            I => \N__4604\
        );

    \I__990\ : InMux
    port map (
            O => \N__4607\,
            I => \N__4601\
        );

    \I__989\ : Span4Mux_s2_h
    port map (
            O => \N__4604\,
            I => \N__4598\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4601\,
            I => \N__4595\
        );

    \I__987\ : Span4Mux_v
    port map (
            O => \N__4598\,
            I => \N__4592\
        );

    \I__986\ : Span4Mux_v
    port map (
            O => \N__4595\,
            I => \N__4589\
        );

    \I__985\ : Sp12to4
    port map (
            O => \N__4592\,
            I => \N__4586\
        );

    \I__984\ : Sp12to4
    port map (
            O => \N__4589\,
            I => \N__4583\
        );

    \I__983\ : Span12Mux_s9_h
    port map (
            O => \N__4586\,
            I => \N__4580\
        );

    \I__982\ : Span12Mux_h
    port map (
            O => \N__4583\,
            I => \N__4577\
        );

    \I__981\ : Span12Mux_h
    port map (
            O => \N__4580\,
            I => \N__4574\
        );

    \I__980\ : Span12Mux_v
    port map (
            O => \N__4577\,
            I => \N__4571\
        );

    \I__979\ : Odrv12
    port map (
            O => \N__4574\,
            I => \D_LM_040_in_5\
        );

    \I__978\ : Odrv12
    port map (
            O => \N__4571\,
            I => \D_LM_040_in_5\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__4566\,
            I => \N__4555\
        );

    \I__976\ : InMux
    port map (
            O => \N__4565\,
            I => \N__4549\
        );

    \I__975\ : InMux
    port map (
            O => \N__4564\,
            I => \N__4549\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__4563\,
            I => \N__4546\
        );

    \I__973\ : InMux
    port map (
            O => \N__4562\,
            I => \N__4543\
        );

    \I__972\ : InMux
    port map (
            O => \N__4561\,
            I => \N__4540\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__4560\,
            I => \N__4536\
        );

    \I__970\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4533\
        );

    \I__969\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4530\
        );

    \I__968\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4527\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__4554\,
            I => \N__4522\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4549\,
            I => \N__4519\
        );

    \I__965\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4516\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__4543\,
            I => \N__4511\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__4540\,
            I => \N__4511\
        );

    \I__962\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4508\
        );

    \I__961\ : InMux
    port map (
            O => \N__4536\,
            I => \N__4505\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4533\,
            I => \N__4496\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4530\,
            I => \N__4496\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4527\,
            I => \N__4496\
        );

    \I__957\ : InMux
    port map (
            O => \N__4526\,
            I => \N__4493\
        );

    \I__956\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4487\
        );

    \I__955\ : InMux
    port map (
            O => \N__4522\,
            I => \N__4487\
        );

    \I__954\ : Span4Mux_v
    port map (
            O => \N__4519\,
            I => \N__4482\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4516\,
            I => \N__4482\
        );

    \I__952\ : Span4Mux_v
    port map (
            O => \N__4511\,
            I => \N__4473\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4508\,
            I => \N__4473\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__4505\,
            I => \N__4473\
        );

    \I__949\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4470\
        );

    \I__948\ : InMux
    port map (
            O => \N__4503\,
            I => \N__4467\
        );

    \I__947\ : Span4Mux_v
    port map (
            O => \N__4496\,
            I => \N__4461\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4493\,
            I => \N__4461\
        );

    \I__945\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4458\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4487\,
            I => \N__4454\
        );

    \I__943\ : Span4Mux_v
    port map (
            O => \N__4482\,
            I => \N__4445\
        );

    \I__942\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4440\
        );

    \I__941\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4440\
        );

    \I__940\ : Span4Mux_v
    port map (
            O => \N__4473\,
            I => \N__4431\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4470\,
            I => \N__4431\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4467\,
            I => \N__4431\
        );

    \I__937\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4428\
        );

    \I__936\ : Span4Mux_v
    port map (
            O => \N__4461\,
            I => \N__4422\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4458\,
            I => \N__4422\
        );

    \I__934\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4419\
        );

    \I__933\ : Span4Mux_v
    port map (
            O => \N__4454\,
            I => \N__4416\
        );

    \I__932\ : InMux
    port map (
            O => \N__4453\,
            I => \N__4413\
        );

    \I__931\ : InMux
    port map (
            O => \N__4452\,
            I => \N__4410\
        );

    \I__930\ : InMux
    port map (
            O => \N__4451\,
            I => \N__4404\
        );

    \I__929\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4404\
        );

    \I__928\ : InMux
    port map (
            O => \N__4449\,
            I => \N__4401\
        );

    \I__927\ : InMux
    port map (
            O => \N__4448\,
            I => \N__4397\
        );

    \I__926\ : Span4Mux_v
    port map (
            O => \N__4445\,
            I => \N__4392\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4440\,
            I => \N__4392\
        );

    \I__924\ : InMux
    port map (
            O => \N__4439\,
            I => \N__4387\
        );

    \I__923\ : InMux
    port map (
            O => \N__4438\,
            I => \N__4387\
        );

    \I__922\ : Span4Mux_v
    port map (
            O => \N__4431\,
            I => \N__4382\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4428\,
            I => \N__4382\
        );

    \I__920\ : InMux
    port map (
            O => \N__4427\,
            I => \N__4379\
        );

    \I__919\ : Span4Mux_v
    port map (
            O => \N__4422\,
            I => \N__4374\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4419\,
            I => \N__4374\
        );

    \I__917\ : Span4Mux_v
    port map (
            O => \N__4416\,
            I => \N__4367\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4413\,
            I => \N__4367\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__4410\,
            I => \N__4367\
        );

    \I__914\ : InMux
    port map (
            O => \N__4409\,
            I => \N__4364\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4404\,
            I => \N__4358\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__4401\,
            I => \N__4358\
        );

    \I__911\ : IoInMux
    port map (
            O => \N__4400\,
            I => \N__4355\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4397\,
            I => \N__4352\
        );

    \I__909\ : Span4Mux_v
    port map (
            O => \N__4392\,
            I => \N__4347\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4387\,
            I => \N__4347\
        );

    \I__907\ : Span4Mux_v
    port map (
            O => \N__4382\,
            I => \N__4342\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4379\,
            I => \N__4342\
        );

    \I__905\ : Span4Mux_v
    port map (
            O => \N__4374\,
            I => \N__4338\
        );

    \I__904\ : Span4Mux_v
    port map (
            O => \N__4367\,
            I => \N__4333\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4364\,
            I => \N__4333\
        );

    \I__902\ : InMux
    port map (
            O => \N__4363\,
            I => \N__4330\
        );

    \I__901\ : Span12Mux_h
    port map (
            O => \N__4358\,
            I => \N__4327\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4355\,
            I => \N__4324\
        );

    \I__899\ : Span12Mux_h
    port map (
            O => \N__4352\,
            I => \N__4321\
        );

    \I__898\ : Span4Mux_v
    port map (
            O => \N__4347\,
            I => \N__4318\
        );

    \I__897\ : Span4Mux_v
    port map (
            O => \N__4342\,
            I => \N__4315\
        );

    \I__896\ : InMux
    port map (
            O => \N__4341\,
            I => \N__4312\
        );

    \I__895\ : Span4Mux_h
    port map (
            O => \N__4338\,
            I => \N__4305\
        );

    \I__894\ : Span4Mux_v
    port map (
            O => \N__4333\,
            I => \N__4305\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4330\,
            I => \N__4305\
        );

    \I__892\ : Span12Mux_v
    port map (
            O => \N__4327\,
            I => \N__4302\
        );

    \I__891\ : Span4Mux_s3_v
    port map (
            O => \N__4324\,
            I => \N__4299\
        );

    \I__890\ : Span12Mux_v
    port map (
            O => \N__4321\,
            I => \N__4290\
        );

    \I__889\ : Sp12to4
    port map (
            O => \N__4318\,
            I => \N__4290\
        );

    \I__888\ : Sp12to4
    port map (
            O => \N__4315\,
            I => \N__4290\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__4312\,
            I => \N__4290\
        );

    \I__886\ : Span4Mux_v
    port map (
            O => \N__4305\,
            I => \N__4287\
        );

    \I__885\ : Odrv12
    port map (
            O => \N__4302\,
            I => \A_AMIGA_c_1\
        );

    \I__884\ : Odrv4
    port map (
            O => \N__4299\,
            I => \A_AMIGA_c_1\
        );

    \I__883\ : Odrv12
    port map (
            O => \N__4290\,
            I => \A_AMIGA_c_1\
        );

    \I__882\ : Odrv4
    port map (
            O => \N__4287\,
            I => \A_AMIGA_c_1\
        );

    \I__881\ : IoInMux
    port map (
            O => \N__4278\,
            I => \N__4275\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4275\,
            I => \N__4272\
        );

    \I__879\ : Span12Mux_s2_h
    port map (
            O => \N__4272\,
            I => \N__4269\
        );

    \I__878\ : Span12Mux_h
    port map (
            O => \N__4269\,
            I => \N__4266\
        );

    \I__877\ : Odrv12
    port map (
            O => \N__4266\,
            I => \un1_D_UU_040_5\
        );

    \I__876\ : InMux
    port map (
            O => \N__4263\,
            I => \N__4260\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4260\,
            I => \N__4257\
        );

    \I__874\ : Span4Mux_v
    port map (
            O => \N__4257\,
            I => \N__4254\
        );

    \I__873\ : Odrv4
    port map (
            O => \N__4254\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__4251\,
            I => \N__4248\
        );

    \I__871\ : InMux
    port map (
            O => \N__4248\,
            I => \N__4244\
        );

    \I__870\ : InMux
    port map (
            O => \N__4247\,
            I => \N__4241\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4244\,
            I => \N__4237\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4241\,
            I => \N__4234\
        );

    \I__867\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4231\
        );

    \I__866\ : Span4Mux_v
    port map (
            O => \N__4237\,
            I => \N__4228\
        );

    \I__865\ : Span4Mux_v
    port map (
            O => \N__4234\,
            I => \N__4223\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4231\,
            I => \N__4223\
        );

    \I__863\ : Span4Mux_v
    port map (
            O => \N__4228\,
            I => \N__4220\
        );

    \I__862\ : Span4Mux_v
    port map (
            O => \N__4223\,
            I => \N__4217\
        );

    \I__861\ : Sp12to4
    port map (
            O => \N__4220\,
            I => \N__4212\
        );

    \I__860\ : Sp12to4
    port map (
            O => \N__4217\,
            I => \N__4212\
        );

    \I__859\ : Span12Mux_h
    port map (
            O => \N__4212\,
            I => \N__4209\
        );

    \I__858\ : Odrv12
    port map (
            O => \N__4209\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__857\ : IoInMux
    port map (
            O => \N__4206\,
            I => \N__4203\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4203\,
            I => \N__4200\
        );

    \I__855\ : IoSpan4Mux
    port map (
            O => \N__4200\,
            I => \N__4197\
        );

    \I__854\ : Sp12to4
    port map (
            O => \N__4197\,
            I => \N__4194\
        );

    \I__853\ : Span12Mux_s6_v
    port map (
            O => \N__4194\,
            I => \N__4191\
        );

    \I__852\ : Odrv12
    port map (
            O => \N__4191\,
            I => \un1_D_UU_AMIGA_6\
        );

    \I__851\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4185\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4185\,
            I => \N__4182\
        );

    \I__849\ : Span12Mux_h
    port map (
            O => \N__4182\,
            I => \N__4179\
        );

    \I__848\ : Odrv12
    port map (
            O => \N__4179\,
            I => \D_LM_AMIGA_in_0\
        );

    \I__847\ : IoInMux
    port map (
            O => \N__4176\,
            I => \N__4173\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4173\,
            I => \N__4170\
        );

    \I__845\ : IoSpan4Mux
    port map (
            O => \N__4170\,
            I => \N__4167\
        );

    \I__844\ : IoSpan4Mux
    port map (
            O => \N__4167\,
            I => \N__4164\
        );

    \I__843\ : Sp12to4
    port map (
            O => \N__4164\,
            I => \N__4161\
        );

    \I__842\ : Span12Mux_s7_h
    port map (
            O => \N__4161\,
            I => \N__4158\
        );

    \I__841\ : Odrv12
    port map (
            O => \N__4158\,
            I => \un1_D_LM_AMIGA_0\
        );

    \I__840\ : IoInMux
    port map (
            O => \N__4155\,
            I => \N__4152\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4152\,
            I => \N__4149\
        );

    \I__838\ : Span12Mux_s9_h
    port map (
            O => \N__4149\,
            I => \N__4146\
        );

    \I__837\ : Odrv12
    port map (
            O => \N__4146\,
            I => \un1_D_UM_AMIGA_0\
        );

    \I__836\ : SRMux
    port map (
            O => \N__4143\,
            I => \N__4140\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4140\,
            I => \N__4137\
        );

    \I__834\ : Odrv4
    port map (
            O => \N__4137\,
            I => \U111_CYCLE_SM.RESETn_c_i\
        );

    \I__833\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4131\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4131\,
            I => \N__4128\
        );

    \I__831\ : Span4Mux_h
    port map (
            O => \N__4128\,
            I => \N__4125\
        );

    \I__830\ : Sp12to4
    port map (
            O => \N__4125\,
            I => \N__4122\
        );

    \I__829\ : Span12Mux_v
    port map (
            O => \N__4122\,
            I => \N__4118\
        );

    \I__828\ : InMux
    port map (
            O => \N__4121\,
            I => \N__4115\
        );

    \I__827\ : Odrv12
    port map (
            O => \N__4118\,
            I => \U111_CYCLE_SM.A_OUTZ0\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4115\,
            I => \U111_CYCLE_SM.A_OUTZ0\
        );

    \I__825\ : InMux
    port map (
            O => \N__4110\,
            I => \N__4107\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4107\,
            I => \U111_CYCLE_SM.A_OUT_0\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__4104\,
            I => \N__4101\
        );

    \I__822\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4098\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4098\,
            I => \N__4095\
        );

    \I__820\ : Span4Mux_v
    port map (
            O => \N__4095\,
            I => \N__4091\
        );

    \I__819\ : InMux
    port map (
            O => \N__4094\,
            I => \N__4088\
        );

    \I__818\ : Span4Mux_v
    port map (
            O => \N__4091\,
            I => \N__4085\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4088\,
            I => \N__4082\
        );

    \I__816\ : Span4Mux_v
    port map (
            O => \N__4085\,
            I => \N__4078\
        );

    \I__815\ : Span4Mux_v
    port map (
            O => \N__4082\,
            I => \N__4075\
        );

    \I__814\ : InMux
    port map (
            O => \N__4081\,
            I => \N__4072\
        );

    \I__813\ : Sp12to4
    port map (
            O => \N__4078\,
            I => \N__4065\
        );

    \I__812\ : Sp12to4
    port map (
            O => \N__4075\,
            I => \N__4065\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4072\,
            I => \N__4065\
        );

    \I__810\ : Span12Mux_h
    port map (
            O => \N__4065\,
            I => \N__4062\
        );

    \I__809\ : Odrv12
    port map (
            O => \N__4062\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__808\ : InMux
    port map (
            O => \N__4059\,
            I => \N__4056\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4056\,
            I => \N__4053\
        );

    \I__806\ : Odrv12
    port map (
            O => \N__4053\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__805\ : InMux
    port map (
            O => \N__4050\,
            I => \N__4047\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__4047\,
            I => \N__4044\
        );

    \I__803\ : Span4Mux_v
    port map (
            O => \N__4044\,
            I => \N__4041\
        );

    \I__802\ : Sp12to4
    port map (
            O => \N__4041\,
            I => \N__4038\
        );

    \I__801\ : Span12Mux_h
    port map (
            O => \N__4038\,
            I => \N__4035\
        );

    \I__800\ : Odrv12
    port map (
            O => \N__4035\,
            I => \D_LM_AMIGA_in_4\
        );

    \I__799\ : IoInMux
    port map (
            O => \N__4032\,
            I => \N__4029\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4029\,
            I => \N__4026\
        );

    \I__797\ : IoSpan4Mux
    port map (
            O => \N__4026\,
            I => \N__4023\
        );

    \I__796\ : IoSpan4Mux
    port map (
            O => \N__4023\,
            I => \N__4020\
        );

    \I__795\ : Span4Mux_s2_h
    port map (
            O => \N__4020\,
            I => \N__4017\
        );

    \I__794\ : Sp12to4
    port map (
            O => \N__4017\,
            I => \N__4014\
        );

    \I__793\ : Span12Mux_s10_h
    port map (
            O => \N__4014\,
            I => \N__4011\
        );

    \I__792\ : Odrv12
    port map (
            O => \N__4011\,
            I => \un1_D_LM_AMIGA_4\
        );

    \I__791\ : InMux
    port map (
            O => \N__4008\,
            I => \N__4005\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4005\,
            I => \N__4002\
        );

    \I__789\ : Span4Mux_v
    port map (
            O => \N__4002\,
            I => \N__3999\
        );

    \I__788\ : Span4Mux_v
    port map (
            O => \N__3999\,
            I => \N__3996\
        );

    \I__787\ : Sp12to4
    port map (
            O => \N__3996\,
            I => \N__3993\
        );

    \I__786\ : Span12Mux_h
    port map (
            O => \N__3993\,
            I => \N__3990\
        );

    \I__785\ : Odrv12
    port map (
            O => \N__3990\,
            I => \D_UU_040_in_1\
        );

    \I__784\ : IoInMux
    port map (
            O => \N__3987\,
            I => \N__3983\
        );

    \I__783\ : InMux
    port map (
            O => \N__3986\,
            I => \N__3980\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__3983\,
            I => \N__3977\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__3980\,
            I => \N__3974\
        );

    \I__780\ : Span4Mux_s3_h
    port map (
            O => \N__3977\,
            I => \N__3971\
        );

    \I__779\ : Span4Mux_h
    port map (
            O => \N__3974\,
            I => \N__3968\
        );

    \I__778\ : Sp12to4
    port map (
            O => \N__3971\,
            I => \N__3965\
        );

    \I__777\ : Sp12to4
    port map (
            O => \N__3968\,
            I => \N__3962\
        );

    \I__776\ : Span12Mux_v
    port map (
            O => \N__3965\,
            I => \N__3959\
        );

    \I__775\ : Span12Mux_v
    port map (
            O => \N__3962\,
            I => \N__3956\
        );

    \I__774\ : Span12Mux_h
    port map (
            O => \N__3959\,
            I => \N__3951\
        );

    \I__773\ : Span12Mux_v
    port map (
            O => \N__3956\,
            I => \N__3951\
        );

    \I__772\ : Span12Mux_h
    port map (
            O => \N__3951\,
            I => \N__3948\
        );

    \I__771\ : Odrv12
    port map (
            O => \N__3948\,
            I => \D_LM_040_in_1\
        );

    \I__770\ : IoInMux
    port map (
            O => \N__3945\,
            I => \N__3942\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__3942\,
            I => \N__3939\
        );

    \I__768\ : IoSpan4Mux
    port map (
            O => \N__3939\,
            I => \N__3936\
        );

    \I__767\ : Sp12to4
    port map (
            O => \N__3936\,
            I => \N__3933\
        );

    \I__766\ : Span12Mux_s6_h
    port map (
            O => \N__3933\,
            I => \N__3930\
        );

    \I__765\ : Odrv12
    port map (
            O => \N__3930\,
            I => \un1_D_UU_040_1\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__3927\,
            I => \N__3924\
        );

    \I__763\ : InMux
    port map (
            O => \N__3924\,
            I => \N__3921\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__3921\,
            I => \N__3918\
        );

    \I__761\ : Span4Mux_v
    port map (
            O => \N__3918\,
            I => \N__3915\
        );

    \I__760\ : Sp12to4
    port map (
            O => \N__3915\,
            I => \N__3912\
        );

    \I__759\ : Span12Mux_h
    port map (
            O => \N__3912\,
            I => \N__3909\
        );

    \I__758\ : Odrv12
    port map (
            O => \N__3909\,
            I => \D_UU_040_in_2\
        );

    \I__757\ : InMux
    port map (
            O => \N__3906\,
            I => \N__3902\
        );

    \I__756\ : IoInMux
    port map (
            O => \N__3905\,
            I => \N__3899\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__3902\,
            I => \N__3896\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__3899\,
            I => \N__3893\
        );

    \I__753\ : Sp12to4
    port map (
            O => \N__3896\,
            I => \N__3890\
        );

    \I__752\ : Span12Mux_s9_h
    port map (
            O => \N__3893\,
            I => \N__3887\
        );

    \I__751\ : Span12Mux_v
    port map (
            O => \N__3890\,
            I => \N__3884\
        );

    \I__750\ : Span12Mux_v
    port map (
            O => \N__3887\,
            I => \N__3881\
        );

    \I__749\ : Span12Mux_v
    port map (
            O => \N__3884\,
            I => \N__3878\
        );

    \I__748\ : Span12Mux_h
    port map (
            O => \N__3881\,
            I => \N__3875\
        );

    \I__747\ : Span12Mux_h
    port map (
            O => \N__3878\,
            I => \N__3872\
        );

    \I__746\ : Odrv12
    port map (
            O => \N__3875\,
            I => \D_LM_040_in_2\
        );

    \I__745\ : Odrv12
    port map (
            O => \N__3872\,
            I => \D_LM_040_in_2\
        );

    \I__744\ : IoInMux
    port map (
            O => \N__3867\,
            I => \N__3864\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3864\,
            I => \N__3861\
        );

    \I__742\ : IoSpan4Mux
    port map (
            O => \N__3861\,
            I => \N__3858\
        );

    \I__741\ : IoSpan4Mux
    port map (
            O => \N__3858\,
            I => \N__3855\
        );

    \I__740\ : Span4Mux_s2_v
    port map (
            O => \N__3855\,
            I => \N__3852\
        );

    \I__739\ : Span4Mux_v
    port map (
            O => \N__3852\,
            I => \N__3849\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__3849\,
            I => \un1_D_UU_040_2\
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__3846\,
            I => \N__3843\
        );

    \I__736\ : InMux
    port map (
            O => \N__3843\,
            I => \N__3840\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__3840\,
            I => \N__3837\
        );

    \I__734\ : Span4Mux_v
    port map (
            O => \N__3837\,
            I => \N__3834\
        );

    \I__733\ : Span4Mux_h
    port map (
            O => \N__3834\,
            I => \N__3831\
        );

    \I__732\ : Sp12to4
    port map (
            O => \N__3831\,
            I => \N__3828\
        );

    \I__731\ : Odrv12
    port map (
            O => \N__3828\,
            I => \D_LL_AMIGA_in_6\
        );

    \I__730\ : IoInMux
    port map (
            O => \N__3825\,
            I => \N__3822\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3822\,
            I => \N__3819\
        );

    \I__728\ : Span4Mux_s3_h
    port map (
            O => \N__3819\,
            I => \N__3816\
        );

    \I__727\ : Span4Mux_v
    port map (
            O => \N__3816\,
            I => \N__3813\
        );

    \I__726\ : Span4Mux_v
    port map (
            O => \N__3813\,
            I => \N__3810\
        );

    \I__725\ : Span4Mux_h
    port map (
            O => \N__3810\,
            I => \N__3807\
        );

    \I__724\ : Sp12to4
    port map (
            O => \N__3807\,
            I => \N__3804\
        );

    \I__723\ : Odrv12
    port map (
            O => \N__3804\,
            I => \un1_D_LL_AMIGA_6\
        );

    \I__722\ : InMux
    port map (
            O => \N__3801\,
            I => \N__3797\
        );

    \I__721\ : IoInMux
    port map (
            O => \N__3800\,
            I => \N__3794\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__3797\,
            I => \N__3791\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3794\,
            I => \N__3788\
        );

    \I__718\ : Span4Mux_v
    port map (
            O => \N__3791\,
            I => \N__3785\
        );

    \I__717\ : Span4Mux_s3_h
    port map (
            O => \N__3788\,
            I => \N__3782\
        );

    \I__716\ : Sp12to4
    port map (
            O => \N__3785\,
            I => \N__3779\
        );

    \I__715\ : Sp12to4
    port map (
            O => \N__3782\,
            I => \N__3776\
        );

    \I__714\ : Span12Mux_h
    port map (
            O => \N__3779\,
            I => \N__3773\
        );

    \I__713\ : Span12Mux_v
    port map (
            O => \N__3776\,
            I => \N__3770\
        );

    \I__712\ : Span12Mux_v
    port map (
            O => \N__3773\,
            I => \N__3767\
        );

    \I__711\ : Span12Mux_h
    port map (
            O => \N__3770\,
            I => \N__3764\
        );

    \I__710\ : Span12Mux_v
    port map (
            O => \N__3767\,
            I => \N__3759\
        );

    \I__709\ : Span12Mux_h
    port map (
            O => \N__3764\,
            I => \N__3759\
        );

    \I__708\ : Odrv12
    port map (
            O => \N__3759\,
            I => \D_LL_040_in_3\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__3756\,
            I => \N__3753\
        );

    \I__706\ : InMux
    port map (
            O => \N__3753\,
            I => \N__3750\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__3750\,
            I => \N__3747\
        );

    \I__704\ : Span4Mux_h
    port map (
            O => \N__3747\,
            I => \N__3744\
        );

    \I__703\ : Sp12to4
    port map (
            O => \N__3744\,
            I => \N__3741\
        );

    \I__702\ : Span12Mux_v
    port map (
            O => \N__3741\,
            I => \N__3738\
        );

    \I__701\ : Span12Mux_h
    port map (
            O => \N__3738\,
            I => \N__3735\
        );

    \I__700\ : Odrv12
    port map (
            O => \N__3735\,
            I => \D_UM_040_in_3\
        );

    \I__699\ : IoInMux
    port map (
            O => \N__3732\,
            I => \N__3729\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3729\,
            I => \N__3726\
        );

    \I__697\ : IoSpan4Mux
    port map (
            O => \N__3726\,
            I => \N__3723\
        );

    \I__696\ : Span4Mux_s3_h
    port map (
            O => \N__3723\,
            I => \N__3720\
        );

    \I__695\ : Span4Mux_h
    port map (
            O => \N__3720\,
            I => \N__3717\
        );

    \I__694\ : Span4Mux_h
    port map (
            O => \N__3717\,
            I => \N__3714\
        );

    \I__693\ : Odrv4
    port map (
            O => \N__3714\,
            I => \un1_D_UM_040_3\
        );

    \I__692\ : InMux
    port map (
            O => \N__3711\,
            I => \N__3708\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__3708\,
            I => \N__3705\
        );

    \I__690\ : Span4Mux_v
    port map (
            O => \N__3705\,
            I => \N__3702\
        );

    \I__689\ : Span4Mux_h
    port map (
            O => \N__3702\,
            I => \N__3699\
        );

    \I__688\ : Sp12to4
    port map (
            O => \N__3699\,
            I => \N__3696\
        );

    \I__687\ : Odrv12
    port map (
            O => \N__3696\,
            I => \D_LL_AMIGA_in_3\
        );

    \I__686\ : IoInMux
    port map (
            O => \N__3693\,
            I => \N__3690\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3690\,
            I => \N__3687\
        );

    \I__684\ : IoSpan4Mux
    port map (
            O => \N__3687\,
            I => \N__3684\
        );

    \I__683\ : Sp12to4
    port map (
            O => \N__3684\,
            I => \N__3681\
        );

    \I__682\ : Span12Mux_s7_v
    port map (
            O => \N__3681\,
            I => \N__3678\
        );

    \I__681\ : Span12Mux_h
    port map (
            O => \N__3678\,
            I => \N__3675\
        );

    \I__680\ : Odrv12
    port map (
            O => \N__3675\,
            I => \un1_D_LL_AMIGA_3\
        );

    \I__679\ : InMux
    port map (
            O => \N__3672\,
            I => \N__3669\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3669\,
            I => \N__3666\
        );

    \I__677\ : Span4Mux_v
    port map (
            O => \N__3666\,
            I => \N__3663\
        );

    \I__676\ : Sp12to4
    port map (
            O => \N__3663\,
            I => \N__3660\
        );

    \I__675\ : Span12Mux_h
    port map (
            O => \N__3660\,
            I => \N__3657\
        );

    \I__674\ : Odrv12
    port map (
            O => \N__3657\,
            I => \D_LL_AMIGA_in_1\
        );

    \I__673\ : IoInMux
    port map (
            O => \N__3654\,
            I => \N__3651\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3651\,
            I => \N__3648\
        );

    \I__671\ : IoSpan4Mux
    port map (
            O => \N__3648\,
            I => \N__3645\
        );

    \I__670\ : Span4Mux_s3_h
    port map (
            O => \N__3645\,
            I => \N__3642\
        );

    \I__669\ : Sp12to4
    port map (
            O => \N__3642\,
            I => \N__3639\
        );

    \I__668\ : Span12Mux_h
    port map (
            O => \N__3639\,
            I => \N__3636\
        );

    \I__667\ : Odrv12
    port map (
            O => \N__3636\,
            I => \un1_D_LL_AMIGA_1\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__3633\,
            I => \N__3630\
        );

    \I__665\ : InMux
    port map (
            O => \N__3630\,
            I => \N__3627\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3627\,
            I => \N__3624\
        );

    \I__663\ : Span4Mux_v
    port map (
            O => \N__3624\,
            I => \N__3621\
        );

    \I__662\ : Sp12to4
    port map (
            O => \N__3621\,
            I => \N__3618\
        );

    \I__661\ : Span12Mux_h
    port map (
            O => \N__3618\,
            I => \N__3615\
        );

    \I__660\ : Odrv12
    port map (
            O => \N__3615\,
            I => \D_LL_AMIGA_in_5\
        );

    \I__659\ : IoInMux
    port map (
            O => \N__3612\,
            I => \N__3609\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3609\,
            I => \N__3606\
        );

    \I__657\ : Span4Mux_s1_h
    port map (
            O => \N__3606\,
            I => \N__3603\
        );

    \I__656\ : Span4Mux_h
    port map (
            O => \N__3603\,
            I => \N__3600\
        );

    \I__655\ : Sp12to4
    port map (
            O => \N__3600\,
            I => \N__3597\
        );

    \I__654\ : Span12Mux_s9_v
    port map (
            O => \N__3597\,
            I => \N__3594\
        );

    \I__653\ : Span12Mux_h
    port map (
            O => \N__3594\,
            I => \N__3591\
        );

    \I__652\ : Odrv12
    port map (
            O => \N__3591\,
            I => \un1_D_LL_AMIGA_5\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__3588\,
            I => \N__3585\
        );

    \I__650\ : InMux
    port map (
            O => \N__3585\,
            I => \N__3582\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__3582\,
            I => \N__3579\
        );

    \I__648\ : Span12Mux_v
    port map (
            O => \N__3579\,
            I => \N__3576\
        );

    \I__647\ : Odrv12
    port map (
            O => \N__3576\,
            I => \D_LL_AMIGA_in_4\
        );

    \I__646\ : IoInMux
    port map (
            O => \N__3573\,
            I => \N__3570\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3570\,
            I => \N__3567\
        );

    \I__644\ : IoSpan4Mux
    port map (
            O => \N__3567\,
            I => \N__3564\
        );

    \I__643\ : Span4Mux_s0_h
    port map (
            O => \N__3564\,
            I => \N__3561\
        );

    \I__642\ : Sp12to4
    port map (
            O => \N__3561\,
            I => \N__3558\
        );

    \I__641\ : Span12Mux_s8_v
    port map (
            O => \N__3558\,
            I => \N__3555\
        );

    \I__640\ : Span12Mux_h
    port map (
            O => \N__3555\,
            I => \N__3552\
        );

    \I__639\ : Odrv12
    port map (
            O => \N__3552\,
            I => \un1_D_LL_AMIGA_4\
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__3549\,
            I => \N__3546\
        );

    \I__637\ : InMux
    port map (
            O => \N__3546\,
            I => \N__3543\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__3543\,
            I => \N__3540\
        );

    \I__635\ : Span12Mux_h
    port map (
            O => \N__3540\,
            I => \N__3537\
        );

    \I__634\ : Odrv12
    port map (
            O => \N__3537\,
            I => \D_UM_040_in_2\
        );

    \I__633\ : IoInMux
    port map (
            O => \N__3534\,
            I => \N__3531\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3531\,
            I => \N__3527\
        );

    \I__631\ : InMux
    port map (
            O => \N__3530\,
            I => \N__3524\
        );

    \I__630\ : IoSpan4Mux
    port map (
            O => \N__3527\,
            I => \N__3521\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3524\,
            I => \N__3518\
        );

    \I__628\ : Span4Mux_s2_h
    port map (
            O => \N__3521\,
            I => \N__3515\
        );

    \I__627\ : Span4Mux_v
    port map (
            O => \N__3518\,
            I => \N__3512\
        );

    \I__626\ : Sp12to4
    port map (
            O => \N__3515\,
            I => \N__3509\
        );

    \I__625\ : Sp12to4
    port map (
            O => \N__3512\,
            I => \N__3506\
        );

    \I__624\ : Span12Mux_h
    port map (
            O => \N__3509\,
            I => \N__3503\
        );

    \I__623\ : Span12Mux_h
    port map (
            O => \N__3506\,
            I => \N__3500\
        );

    \I__622\ : Span12Mux_h
    port map (
            O => \N__3503\,
            I => \N__3495\
        );

    \I__621\ : Span12Mux_v
    port map (
            O => \N__3500\,
            I => \N__3495\
        );

    \I__620\ : Odrv12
    port map (
            O => \N__3495\,
            I => \D_LL_040_in_2\
        );

    \I__619\ : IoInMux
    port map (
            O => \N__3492\,
            I => \N__3489\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3489\,
            I => \N__3486\
        );

    \I__617\ : Span4Mux_s2_h
    port map (
            O => \N__3486\,
            I => \N__3483\
        );

    \I__616\ : Span4Mux_h
    port map (
            O => \N__3483\,
            I => \N__3480\
        );

    \I__615\ : Span4Mux_h
    port map (
            O => \N__3480\,
            I => \N__3477\
        );

    \I__614\ : Span4Mux_v
    port map (
            O => \N__3477\,
            I => \N__3474\
        );

    \I__613\ : Odrv4
    port map (
            O => \N__3474\,
            I => \un1_D_UM_040_2\
        );

    \I__612\ : InMux
    port map (
            O => \N__3471\,
            I => \N__3468\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3468\,
            I => \N__3465\
        );

    \I__610\ : Span12Mux_h
    port map (
            O => \N__3465\,
            I => \N__3462\
        );

    \I__609\ : Odrv12
    port map (
            O => \N__3462\,
            I => \D_LM_AMIGA_in_3\
        );

    \I__608\ : IoInMux
    port map (
            O => \N__3459\,
            I => \N__3456\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3456\,
            I => \N__3453\
        );

    \I__606\ : Span4Mux_s1_h
    port map (
            O => \N__3453\,
            I => \N__3450\
        );

    \I__605\ : Sp12to4
    port map (
            O => \N__3450\,
            I => \N__3447\
        );

    \I__604\ : Span12Mux_v
    port map (
            O => \N__3447\,
            I => \N__3444\
        );

    \I__603\ : Span12Mux_h
    port map (
            O => \N__3444\,
            I => \N__3441\
        );

    \I__602\ : Odrv12
    port map (
            O => \N__3441\,
            I => \un1_D_LM_AMIGA_3\
        );

    \I__601\ : InMux
    port map (
            O => \N__3438\,
            I => \N__3435\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3435\,
            I => \N__3432\
        );

    \I__599\ : Span12Mux_v
    port map (
            O => \N__3432\,
            I => \N__3429\
        );

    \I__598\ : Odrv12
    port map (
            O => \N__3429\,
            I => \D_LM_AMIGA_in_5\
        );

    \I__597\ : IoInMux
    port map (
            O => \N__3426\,
            I => \N__3423\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3423\,
            I => \N__3420\
        );

    \I__595\ : Span4Mux_s2_h
    port map (
            O => \N__3420\,
            I => \N__3417\
        );

    \I__594\ : Sp12to4
    port map (
            O => \N__3417\,
            I => \N__3414\
        );

    \I__593\ : Span12Mux_v
    port map (
            O => \N__3414\,
            I => \N__3411\
        );

    \I__592\ : Span12Mux_h
    port map (
            O => \N__3411\,
            I => \N__3408\
        );

    \I__591\ : Odrv12
    port map (
            O => \N__3408\,
            I => \un1_D_LM_AMIGA_5\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__3405\,
            I => \N__3402\
        );

    \I__589\ : InMux
    port map (
            O => \N__3402\,
            I => \N__3399\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3399\,
            I => \N__3396\
        );

    \I__587\ : Span4Mux_v
    port map (
            O => \N__3396\,
            I => \N__3393\
        );

    \I__586\ : Span4Mux_v
    port map (
            O => \N__3393\,
            I => \N__3390\
        );

    \I__585\ : Sp12to4
    port map (
            O => \N__3390\,
            I => \N__3387\
        );

    \I__584\ : Span12Mux_h
    port map (
            O => \N__3387\,
            I => \N__3384\
        );

    \I__583\ : Odrv12
    port map (
            O => \N__3384\,
            I => \D_UU_040_in_4\
        );

    \I__582\ : IoInMux
    port map (
            O => \N__3381\,
            I => \N__3378\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3378\,
            I => \N__3375\
        );

    \I__580\ : Span4Mux_s1_h
    port map (
            O => \N__3375\,
            I => \N__3372\
        );

    \I__579\ : Sp12to4
    port map (
            O => \N__3372\,
            I => \N__3368\
        );

    \I__578\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3365\
        );

    \I__577\ : Span12Mux_v
    port map (
            O => \N__3368\,
            I => \N__3362\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3365\,
            I => \N__3359\
        );

    \I__575\ : Span12Mux_h
    port map (
            O => \N__3362\,
            I => \N__3356\
        );

    \I__574\ : Span12Mux_h
    port map (
            O => \N__3359\,
            I => \N__3353\
        );

    \I__573\ : Span12Mux_h
    port map (
            O => \N__3356\,
            I => \N__3350\
        );

    \I__572\ : Span12Mux_v
    port map (
            O => \N__3353\,
            I => \N__3347\
        );

    \I__571\ : Odrv12
    port map (
            O => \N__3350\,
            I => \D_LM_040_in_4\
        );

    \I__570\ : Odrv12
    port map (
            O => \N__3347\,
            I => \D_LM_040_in_4\
        );

    \I__569\ : IoInMux
    port map (
            O => \N__3342\,
            I => \N__3339\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3339\,
            I => \N__3336\
        );

    \I__567\ : Span12Mux_s6_v
    port map (
            O => \N__3336\,
            I => \N__3333\
        );

    \I__566\ : Odrv12
    port map (
            O => \N__3333\,
            I => \un1_D_UU_040_4\
        );

    \I__565\ : InMux
    port map (
            O => \N__3330\,
            I => \N__3327\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__3327\,
            I => \N__3324\
        );

    \I__563\ : Span4Mux_v
    port map (
            O => \N__3324\,
            I => \N__3321\
        );

    \I__562\ : Span4Mux_h
    port map (
            O => \N__3321\,
            I => \N__3318\
        );

    \I__561\ : Sp12to4
    port map (
            O => \N__3318\,
            I => \N__3315\
        );

    \I__560\ : Odrv12
    port map (
            O => \N__3315\,
            I => \D_LL_AMIGA_in_0\
        );

    \I__559\ : IoInMux
    port map (
            O => \N__3312\,
            I => \N__3309\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3309\,
            I => \N__3306\
        );

    \I__557\ : IoSpan4Mux
    port map (
            O => \N__3306\,
            I => \N__3303\
        );

    \I__556\ : Sp12to4
    port map (
            O => \N__3303\,
            I => \N__3300\
        );

    \I__555\ : Span12Mux_s7_h
    port map (
            O => \N__3300\,
            I => \N__3297\
        );

    \I__554\ : Span12Mux_h
    port map (
            O => \N__3297\,
            I => \N__3294\
        );

    \I__553\ : Odrv12
    port map (
            O => \N__3294\,
            I => \un1_D_LL_AMIGA_0\
        );

    \I__552\ : IoInMux
    port map (
            O => \N__3291\,
            I => \N__3288\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3288\,
            I => \N__3285\
        );

    \I__550\ : IoSpan4Mux
    port map (
            O => \N__3285\,
            I => \N__3282\
        );

    \I__549\ : Span4Mux_s2_v
    port map (
            O => \N__3282\,
            I => \N__3279\
        );

    \I__548\ : Odrv4
    port map (
            O => \N__3279\,
            I => \TSn_c\
        );

    \I__547\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3273\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3273\,
            I => \N__3270\
        );

    \I__545\ : Span12Mux_h
    port map (
            O => \N__3270\,
            I => \N__3267\
        );

    \I__544\ : Odrv12
    port map (
            O => \N__3267\,
            I => \D_LM_AMIGA_in_2\
        );

    \I__543\ : IoInMux
    port map (
            O => \N__3264\,
            I => \N__3261\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3261\,
            I => \N__3258\
        );

    \I__541\ : Span12Mux_s2_h
    port map (
            O => \N__3258\,
            I => \N__3255\
        );

    \I__540\ : Span12Mux_h
    port map (
            O => \N__3255\,
            I => \N__3252\
        );

    \I__539\ : Span12Mux_v
    port map (
            O => \N__3252\,
            I => \N__3249\
        );

    \I__538\ : Odrv12
    port map (
            O => \N__3249\,
            I => \un1_D_LM_AMIGA_2\
        );

    \I__537\ : InMux
    port map (
            O => \N__3246\,
            I => \N__3243\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3243\,
            I => \N__3240\
        );

    \I__535\ : Sp12to4
    port map (
            O => \N__3240\,
            I => \N__3237\
        );

    \I__534\ : Span12Mux_v
    port map (
            O => \N__3237\,
            I => \N__3234\
        );

    \I__533\ : Span12Mux_h
    port map (
            O => \N__3234\,
            I => \N__3231\
        );

    \I__532\ : Odrv12
    port map (
            O => \N__3231\,
            I => \D_LM_AMIGA_in_6\
        );

    \I__531\ : IoInMux
    port map (
            O => \N__3228\,
            I => \N__3225\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3225\,
            I => \N__3222\
        );

    \I__529\ : IoSpan4Mux
    port map (
            O => \N__3222\,
            I => \N__3219\
        );

    \I__528\ : Span4Mux_s0_h
    port map (
            O => \N__3219\,
            I => \N__3216\
        );

    \I__527\ : Sp12to4
    port map (
            O => \N__3216\,
            I => \N__3213\
        );

    \I__526\ : Span12Mux_s8_h
    port map (
            O => \N__3213\,
            I => \N__3210\
        );

    \I__525\ : Odrv12
    port map (
            O => \N__3210\,
            I => \un1_D_LM_AMIGA_6\
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__3207\,
            I => \N__3204\
        );

    \I__523\ : InMux
    port map (
            O => \N__3204\,
            I => \N__3201\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3201\,
            I => \N__3198\
        );

    \I__521\ : Odrv12
    port map (
            O => \N__3198\,
            I => \D_LM_AMIGA_in_1\
        );

    \I__520\ : IoInMux
    port map (
            O => \N__3195\,
            I => \N__3192\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3192\,
            I => \N__3189\
        );

    \I__518\ : Span4Mux_s2_h
    port map (
            O => \N__3189\,
            I => \N__3186\
        );

    \I__517\ : Span4Mux_h
    port map (
            O => \N__3186\,
            I => \N__3183\
        );

    \I__516\ : Sp12to4
    port map (
            O => \N__3183\,
            I => \N__3180\
        );

    \I__515\ : Span12Mux_v
    port map (
            O => \N__3180\,
            I => \N__3177\
        );

    \I__514\ : Span12Mux_h
    port map (
            O => \N__3177\,
            I => \N__3174\
        );

    \I__513\ : Odrv12
    port map (
            O => \N__3174\,
            I => \un1_D_LM_AMIGA_1\
        );

    \I__512\ : InMux
    port map (
            O => \N__3171\,
            I => \N__3168\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3168\,
            I => \N__3165\
        );

    \I__510\ : Span12Mux_v
    port map (
            O => \N__3165\,
            I => \N__3162\
        );

    \I__509\ : Span12Mux_h
    port map (
            O => \N__3162\,
            I => \N__3159\
        );

    \I__508\ : Odrv12
    port map (
            O => \N__3159\,
            I => \D_UM_040_in_6\
        );

    \I__507\ : IoInMux
    port map (
            O => \N__3156\,
            I => \N__3153\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3153\,
            I => \N__3150\
        );

    \I__505\ : IoSpan4Mux
    port map (
            O => \N__3150\,
            I => \N__3146\
        );

    \I__504\ : CascadeMux
    port map (
            O => \N__3149\,
            I => \N__3143\
        );

    \I__503\ : IoSpan4Mux
    port map (
            O => \N__3146\,
            I => \N__3140\
        );

    \I__502\ : InMux
    port map (
            O => \N__3143\,
            I => \N__3137\
        );

    \I__501\ : Span4Mux_s2_h
    port map (
            O => \N__3140\,
            I => \N__3134\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3137\,
            I => \N__3131\
        );

    \I__499\ : Sp12to4
    port map (
            O => \N__3134\,
            I => \N__3128\
        );

    \I__498\ : Span12Mux_v
    port map (
            O => \N__3131\,
            I => \N__3125\
        );

    \I__497\ : Span12Mux_h
    port map (
            O => \N__3128\,
            I => \N__3122\
        );

    \I__496\ : Span12Mux_v
    port map (
            O => \N__3125\,
            I => \N__3119\
        );

    \I__495\ : Span12Mux_h
    port map (
            O => \N__3122\,
            I => \N__3116\
        );

    \I__494\ : Span12Mux_h
    port map (
            O => \N__3119\,
            I => \N__3113\
        );

    \I__493\ : Odrv12
    port map (
            O => \N__3116\,
            I => \D_LL_040_in_6\
        );

    \I__492\ : Odrv12
    port map (
            O => \N__3113\,
            I => \D_LL_040_in_6\
        );

    \I__491\ : IoInMux
    port map (
            O => \N__3108\,
            I => \N__3105\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3105\,
            I => \N__3102\
        );

    \I__489\ : Span12Mux_s2_h
    port map (
            O => \N__3102\,
            I => \N__3099\
        );

    \I__488\ : Span12Mux_v
    port map (
            O => \N__3099\,
            I => \N__3096\
        );

    \I__487\ : Odrv12
    port map (
            O => \N__3096\,
            I => \un1_D_UM_040_6\
        );

    \I__486\ : CascadeMux
    port map (
            O => \N__3093\,
            I => \N__3090\
        );

    \I__485\ : InMux
    port map (
            O => \N__3090\,
            I => \N__3087\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3087\,
            I => \N__3084\
        );

    \I__483\ : Span4Mux_v
    port map (
            O => \N__3084\,
            I => \N__3081\
        );

    \I__482\ : Sp12to4
    port map (
            O => \N__3081\,
            I => \N__3078\
        );

    \I__481\ : Span12Mux_h
    port map (
            O => \N__3078\,
            I => \N__3075\
        );

    \I__480\ : Span12Mux_h
    port map (
            O => \N__3075\,
            I => \N__3072\
        );

    \I__479\ : Odrv12
    port map (
            O => \N__3072\,
            I => \D_UM_040_in_4\
        );

    \I__478\ : IoInMux
    port map (
            O => \N__3069\,
            I => \N__3066\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3066\,
            I => \N__3062\
        );

    \I__476\ : InMux
    port map (
            O => \N__3065\,
            I => \N__3059\
        );

    \I__475\ : Span4Mux_s2_h
    port map (
            O => \N__3062\,
            I => \N__3056\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3059\,
            I => \N__3053\
        );

    \I__473\ : Span4Mux_v
    port map (
            O => \N__3056\,
            I => \N__3050\
        );

    \I__472\ : Span12Mux_v
    port map (
            O => \N__3053\,
            I => \N__3047\
        );

    \I__471\ : Sp12to4
    port map (
            O => \N__3050\,
            I => \N__3044\
        );

    \I__470\ : Span12Mux_v
    port map (
            O => \N__3047\,
            I => \N__3041\
        );

    \I__469\ : Span12Mux_h
    port map (
            O => \N__3044\,
            I => \N__3038\
        );

    \I__468\ : Span12Mux_h
    port map (
            O => \N__3041\,
            I => \N__3035\
        );

    \I__467\ : Span12Mux_h
    port map (
            O => \N__3038\,
            I => \N__3032\
        );

    \I__466\ : Odrv12
    port map (
            O => \N__3035\,
            I => \D_LL_040_in_4\
        );

    \I__465\ : Odrv12
    port map (
            O => \N__3032\,
            I => \D_LL_040_in_4\
        );

    \I__464\ : IoInMux
    port map (
            O => \N__3027\,
            I => \N__3024\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__3024\,
            I => \N__3021\
        );

    \I__462\ : Span4Mux_s1_h
    port map (
            O => \N__3021\,
            I => \N__3018\
        );

    \I__461\ : Span4Mux_h
    port map (
            O => \N__3018\,
            I => \N__3015\
        );

    \I__460\ : Span4Mux_h
    port map (
            O => \N__3015\,
            I => \N__3012\
        );

    \I__459\ : Odrv4
    port map (
            O => \N__3012\,
            I => \un1_D_UM_040_4\
        );

    \I__458\ : InMux
    port map (
            O => \N__3009\,
            I => \N__3006\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3006\,
            I => \N__3003\
        );

    \I__456\ : Span4Mux_v
    port map (
            O => \N__3003\,
            I => \N__3000\
        );

    \I__455\ : Span4Mux_h
    port map (
            O => \N__3000\,
            I => \N__2997\
        );

    \I__454\ : Span4Mux_h
    port map (
            O => \N__2997\,
            I => \N__2994\
        );

    \I__453\ : Sp12to4
    port map (
            O => \N__2994\,
            I => \N__2991\
        );

    \I__452\ : Span12Mux_h
    port map (
            O => \N__2991\,
            I => \N__2988\
        );

    \I__451\ : Odrv12
    port map (
            O => \N__2988\,
            I => \D_UU_040_in_3\
        );

    \I__450\ : IoInMux
    port map (
            O => \N__2985\,
            I => \N__2982\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2982\,
            I => \N__2979\
        );

    \I__448\ : IoSpan4Mux
    port map (
            O => \N__2979\,
            I => \N__2976\
        );

    \I__447\ : IoSpan4Mux
    port map (
            O => \N__2976\,
            I => \N__2972\
        );

    \I__446\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2969\
        );

    \I__445\ : Span4Mux_s2_h
    port map (
            O => \N__2972\,
            I => \N__2966\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2969\,
            I => \N__2963\
        );

    \I__443\ : Sp12to4
    port map (
            O => \N__2966\,
            I => \N__2960\
        );

    \I__442\ : Span12Mux_s10_v
    port map (
            O => \N__2963\,
            I => \N__2957\
        );

    \I__441\ : Span12Mux_h
    port map (
            O => \N__2960\,
            I => \N__2954\
        );

    \I__440\ : Span12Mux_v
    port map (
            O => \N__2957\,
            I => \N__2951\
        );

    \I__439\ : Span12Mux_h
    port map (
            O => \N__2954\,
            I => \N__2948\
        );

    \I__438\ : Span12Mux_h
    port map (
            O => \N__2951\,
            I => \N__2945\
        );

    \I__437\ : Odrv12
    port map (
            O => \N__2948\,
            I => \D_LM_040_in_3\
        );

    \I__436\ : Odrv12
    port map (
            O => \N__2945\,
            I => \D_LM_040_in_3\
        );

    \I__435\ : IoInMux
    port map (
            O => \N__2940\,
            I => \N__2937\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__2937\,
            I => \N__2934\
        );

    \I__433\ : IoSpan4Mux
    port map (
            O => \N__2934\,
            I => \N__2931\
        );

    \I__432\ : IoSpan4Mux
    port map (
            O => \N__2931\,
            I => \N__2928\
        );

    \I__431\ : Span4Mux_s2_v
    port map (
            O => \N__2928\,
            I => \N__2925\
        );

    \I__430\ : Span4Mux_v
    port map (
            O => \N__2925\,
            I => \N__2922\
        );

    \I__429\ : Odrv4
    port map (
            O => \N__2922\,
            I => \un1_D_UU_040_3\
        );

    \I__428\ : IoInMux
    port map (
            O => \N__2919\,
            I => \N__2916\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2916\,
            I => \N__2913\
        );

    \I__426\ : Span4Mux_s2_h
    port map (
            O => \N__2913\,
            I => \N__2910\
        );

    \I__425\ : Span4Mux_v
    port map (
            O => \N__2910\,
            I => \N__2906\
        );

    \I__424\ : InMux
    port map (
            O => \N__2909\,
            I => \N__2903\
        );

    \I__423\ : Sp12to4
    port map (
            O => \N__2906\,
            I => \N__2900\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2903\,
            I => \N__2897\
        );

    \I__421\ : Span12Mux_h
    port map (
            O => \N__2900\,
            I => \N__2894\
        );

    \I__420\ : Span12Mux_s11_v
    port map (
            O => \N__2897\,
            I => \N__2891\
        );

    \I__419\ : Span12Mux_h
    port map (
            O => \N__2894\,
            I => \N__2888\
        );

    \I__418\ : Span12Mux_h
    port map (
            O => \N__2891\,
            I => \N__2885\
        );

    \I__417\ : Odrv12
    port map (
            O => \N__2888\,
            I => \D_LM_040_in_6\
        );

    \I__416\ : Odrv12
    port map (
            O => \N__2885\,
            I => \D_LM_040_in_6\
        );

    \I__415\ : CascadeMux
    port map (
            O => \N__2880\,
            I => \N__2877\
        );

    \I__414\ : InMux
    port map (
            O => \N__2877\,
            I => \N__2874\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2874\,
            I => \N__2871\
        );

    \I__412\ : Span4Mux_v
    port map (
            O => \N__2871\,
            I => \N__2868\
        );

    \I__411\ : Sp12to4
    port map (
            O => \N__2868\,
            I => \N__2865\
        );

    \I__410\ : Span12Mux_h
    port map (
            O => \N__2865\,
            I => \N__2862\
        );

    \I__409\ : Span12Mux_h
    port map (
            O => \N__2862\,
            I => \N__2859\
        );

    \I__408\ : Odrv12
    port map (
            O => \N__2859\,
            I => \D_UU_040_in_6\
        );

    \I__407\ : IoInMux
    port map (
            O => \N__2856\,
            I => \N__2853\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2853\,
            I => \N__2850\
        );

    \I__405\ : IoSpan4Mux
    port map (
            O => \N__2850\,
            I => \N__2847\
        );

    \I__404\ : Span4Mux_s2_v
    port map (
            O => \N__2847\,
            I => \N__2844\
        );

    \I__403\ : Span4Mux_v
    port map (
            O => \N__2844\,
            I => \N__2841\
        );

    \I__402\ : Odrv4
    port map (
            O => \N__2841\,
            I => \un1_D_UU_040_6\
        );

    \I__401\ : InMux
    port map (
            O => \N__2838\,
            I => \N__2835\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2835\,
            I => \N__2832\
        );

    \I__399\ : Span4Mux_v
    port map (
            O => \N__2832\,
            I => \N__2829\
        );

    \I__398\ : Sp12to4
    port map (
            O => \N__2829\,
            I => \N__2826\
        );

    \I__397\ : Odrv12
    port map (
            O => \N__2826\,
            I => \D_LL_AMIGA_in_7\
        );

    \I__396\ : IoInMux
    port map (
            O => \N__2823\,
            I => \N__2820\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2820\,
            I => \N__2817\
        );

    \I__394\ : IoSpan4Mux
    port map (
            O => \N__2817\,
            I => \N__2814\
        );

    \I__393\ : Sp12to4
    port map (
            O => \N__2814\,
            I => \N__2811\
        );

    \I__392\ : Span12Mux_s9_h
    port map (
            O => \N__2811\,
            I => \N__2808\
        );

    \I__391\ : Span12Mux_h
    port map (
            O => \N__2808\,
            I => \N__2805\
        );

    \I__390\ : Odrv12
    port map (
            O => \N__2805\,
            I => \un1_D_LL_AMIGA_7\
        );

    \I__389\ : IoInMux
    port map (
            O => \N__2802\,
            I => \N__2798\
        );

    \I__388\ : InMux
    port map (
            O => \N__2801\,
            I => \N__2795\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2798\,
            I => \N__2792\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2795\,
            I => \N__2789\
        );

    \I__385\ : Span4Mux_s3_h
    port map (
            O => \N__2792\,
            I => \N__2786\
        );

    \I__384\ : Sp12to4
    port map (
            O => \N__2789\,
            I => \N__2783\
        );

    \I__383\ : Sp12to4
    port map (
            O => \N__2786\,
            I => \N__2780\
        );

    \I__382\ : Span12Mux_v
    port map (
            O => \N__2783\,
            I => \N__2777\
        );

    \I__381\ : Span12Mux_v
    port map (
            O => \N__2780\,
            I => \N__2774\
        );

    \I__380\ : Span12Mux_v
    port map (
            O => \N__2777\,
            I => \N__2771\
        );

    \I__379\ : Span12Mux_h
    port map (
            O => \N__2774\,
            I => \N__2768\
        );

    \I__378\ : Span12Mux_h
    port map (
            O => \N__2771\,
            I => \N__2765\
        );

    \I__377\ : Span12Mux_h
    port map (
            O => \N__2768\,
            I => \N__2762\
        );

    \I__376\ : Odrv12
    port map (
            O => \N__2765\,
            I => \D_LL_040_in_1\
        );

    \I__375\ : Odrv12
    port map (
            O => \N__2762\,
            I => \D_LL_040_in_1\
        );

    \I__374\ : InMux
    port map (
            O => \N__2757\,
            I => \N__2754\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2754\,
            I => \N__2751\
        );

    \I__372\ : Span4Mux_h
    port map (
            O => \N__2751\,
            I => \N__2748\
        );

    \I__371\ : Sp12to4
    port map (
            O => \N__2748\,
            I => \N__2745\
        );

    \I__370\ : Span12Mux_v
    port map (
            O => \N__2745\,
            I => \N__2742\
        );

    \I__369\ : Span12Mux_h
    port map (
            O => \N__2742\,
            I => \N__2739\
        );

    \I__368\ : Odrv12
    port map (
            O => \N__2739\,
            I => \D_UM_040_in_1\
        );

    \I__367\ : IoInMux
    port map (
            O => \N__2736\,
            I => \N__2733\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2733\,
            I => \N__2730\
        );

    \I__365\ : IoSpan4Mux
    port map (
            O => \N__2730\,
            I => \N__2727\
        );

    \I__364\ : Sp12to4
    port map (
            O => \N__2727\,
            I => \N__2724\
        );

    \I__363\ : Odrv12
    port map (
            O => \N__2724\,
            I => \un1_D_UM_040_1\
        );

    \I__362\ : InMux
    port map (
            O => \N__2721\,
            I => \N__2718\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2718\,
            I => \N__2715\
        );

    \I__360\ : Span4Mux_v
    port map (
            O => \N__2715\,
            I => \N__2712\
        );

    \I__359\ : Span4Mux_h
    port map (
            O => \N__2712\,
            I => \N__2709\
        );

    \I__358\ : Sp12to4
    port map (
            O => \N__2709\,
            I => \N__2706\
        );

    \I__357\ : Span12Mux_h
    port map (
            O => \N__2706\,
            I => \N__2703\
        );

    \I__356\ : Odrv12
    port map (
            O => \N__2703\,
            I => \D_UU_040_in_7\
        );

    \I__355\ : IoInMux
    port map (
            O => \N__2700\,
            I => \N__2697\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2697\,
            I => \N__2693\
        );

    \I__353\ : CascadeMux
    port map (
            O => \N__2696\,
            I => \N__2690\
        );

    \I__352\ : IoSpan4Mux
    port map (
            O => \N__2693\,
            I => \N__2687\
        );

    \I__351\ : InMux
    port map (
            O => \N__2690\,
            I => \N__2684\
        );

    \I__350\ : Span4Mux_s2_h
    port map (
            O => \N__2687\,
            I => \N__2681\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2684\,
            I => \N__2678\
        );

    \I__348\ : Sp12to4
    port map (
            O => \N__2681\,
            I => \N__2675\
        );

    \I__347\ : Span4Mux_v
    port map (
            O => \N__2678\,
            I => \N__2672\
        );

    \I__346\ : Span12Mux_h
    port map (
            O => \N__2675\,
            I => \N__2669\
        );

    \I__345\ : Sp12to4
    port map (
            O => \N__2672\,
            I => \N__2666\
        );

    \I__344\ : Span12Mux_h
    port map (
            O => \N__2669\,
            I => \N__2663\
        );

    \I__343\ : Span12Mux_h
    port map (
            O => \N__2666\,
            I => \N__2660\
        );

    \I__342\ : Odrv12
    port map (
            O => \N__2663\,
            I => \D_LM_040_in_7\
        );

    \I__341\ : Odrv12
    port map (
            O => \N__2660\,
            I => \D_LM_040_in_7\
        );

    \I__340\ : IoInMux
    port map (
            O => \N__2655\,
            I => \N__2652\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2652\,
            I => \N__2649\
        );

    \I__338\ : IoSpan4Mux
    port map (
            O => \N__2649\,
            I => \N__2646\
        );

    \I__337\ : Sp12to4
    port map (
            O => \N__2646\,
            I => \N__2643\
        );

    \I__336\ : Span12Mux_s6_v
    port map (
            O => \N__2643\,
            I => \N__2640\
        );

    \I__335\ : Odrv12
    port map (
            O => \N__2640\,
            I => \un1_D_UU_040_7\
        );

    \I__334\ : InMux
    port map (
            O => \N__2637\,
            I => \N__2634\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2634\,
            I => \N__2631\
        );

    \I__332\ : Span4Mux_h
    port map (
            O => \N__2631\,
            I => \N__2628\
        );

    \I__331\ : Span4Mux_v
    port map (
            O => \N__2628\,
            I => \N__2625\
        );

    \I__330\ : Odrv4
    port map (
            O => \N__2625\,
            I => \A_040_c_0\
        );

    \I__329\ : IoInMux
    port map (
            O => \N__2622\,
            I => \N__2619\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2619\,
            I => \N__2616\
        );

    \I__327\ : Span4Mux_s2_v
    port map (
            O => \N__2616\,
            I => \N__2613\
        );

    \I__326\ : Span4Mux_v
    port map (
            O => \N__2613\,
            I => \N__2610\
        );

    \I__325\ : Odrv4
    port map (
            O => \N__2610\,
            I => \A_AMIGA_c_0\
        );

    \I__324\ : InMux
    port map (
            O => \N__2607\,
            I => \N__2604\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2604\,
            I => \N__2601\
        );

    \I__322\ : Span12Mux_h
    port map (
            O => \N__2601\,
            I => \N__2598\
        );

    \I__321\ : Odrv12
    port map (
            O => \N__2598\,
            I => \A_040_c_1\
        );

    \I__320\ : InMux
    port map (
            O => \N__2595\,
            I => \N__2592\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__2592\,
            I => \N__2589\
        );

    \I__318\ : Span12Mux_v
    port map (
            O => \N__2589\,
            I => \N__2586\
        );

    \I__317\ : Odrv12
    port map (
            O => \N__2586\,
            I => \D_LL_AMIGA_in_2\
        );

    \I__316\ : IoInMux
    port map (
            O => \N__2583\,
            I => \N__2580\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2580\,
            I => \N__2577\
        );

    \I__314\ : IoSpan4Mux
    port map (
            O => \N__2577\,
            I => \N__2574\
        );

    \I__313\ : IoSpan4Mux
    port map (
            O => \N__2574\,
            I => \N__2571\
        );

    \I__312\ : Span4Mux_s3_h
    port map (
            O => \N__2571\,
            I => \N__2568\
        );

    \I__311\ : Sp12to4
    port map (
            O => \N__2568\,
            I => \N__2565\
        );

    \I__310\ : Span12Mux_s11_h
    port map (
            O => \N__2565\,
            I => \N__2562\
        );

    \I__309\ : Odrv12
    port map (
            O => \N__2562\,
            I => \un1_D_LL_AMIGA_2\
        );

    \I__308\ : IoInMux
    port map (
            O => \N__2559\,
            I => \N__2552\
        );

    \I__307\ : IoInMux
    port map (
            O => \N__2558\,
            I => \N__2549\
        );

    \I__306\ : IoInMux
    port map (
            O => \N__2557\,
            I => \N__2546\
        );

    \I__305\ : IoInMux
    port map (
            O => \N__2556\,
            I => \N__2539\
        );

    \I__304\ : IoInMux
    port map (
            O => \N__2555\,
            I => \N__2536\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2552\,
            I => \N__2527\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2549\,
            I => \N__2527\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2546\,
            I => \N__2527\
        );

    \I__300\ : IoInMux
    port map (
            O => \N__2545\,
            I => \N__2524\
        );

    \I__299\ : IoInMux
    port map (
            O => \N__2544\,
            I => \N__2521\
        );

    \I__298\ : IoInMux
    port map (
            O => \N__2543\,
            I => \N__2518\
        );

    \I__297\ : IoInMux
    port map (
            O => \N__2542\,
            I => \N__2515\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2539\,
            I => \N__2503\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2536\,
            I => \N__2503\
        );

    \I__294\ : IoInMux
    port map (
            O => \N__2535\,
            I => \N__2500\
        );

    \I__293\ : IoInMux
    port map (
            O => \N__2534\,
            I => \N__2497\
        );

    \I__292\ : IoSpan4Mux
    port map (
            O => \N__2527\,
            I => \N__2486\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2524\,
            I => \N__2486\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2521\,
            I => \N__2486\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2518\,
            I => \N__2486\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2515\,
            I => \N__2486\
        );

    \I__287\ : IoInMux
    port map (
            O => \N__2514\,
            I => \N__2483\
        );

    \I__286\ : IoInMux
    port map (
            O => \N__2513\,
            I => \N__2480\
        );

    \I__285\ : IoInMux
    port map (
            O => \N__2512\,
            I => \N__2477\
        );

    \I__284\ : IoInMux
    port map (
            O => \N__2511\,
            I => \N__2474\
        );

    \I__283\ : IoInMux
    port map (
            O => \N__2510\,
            I => \N__2467\
        );

    \I__282\ : IoInMux
    port map (
            O => \N__2509\,
            I => \N__2464\
        );

    \I__281\ : IoInMux
    port map (
            O => \N__2508\,
            I => \N__2461\
        );

    \I__280\ : IoSpan4Mux
    port map (
            O => \N__2503\,
            I => \N__2454\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2500\,
            I => \N__2454\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2497\,
            I => \N__2451\
        );

    \I__277\ : IoSpan4Mux
    port map (
            O => \N__2486\,
            I => \N__2440\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2483\,
            I => \N__2440\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2480\,
            I => \N__2440\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2477\,
            I => \N__2440\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__2474\,
            I => \N__2440\
        );

    \I__272\ : IoInMux
    port map (
            O => \N__2473\,
            I => \N__2437\
        );

    \I__271\ : IoInMux
    port map (
            O => \N__2472\,
            I => \N__2434\
        );

    \I__270\ : IoInMux
    port map (
            O => \N__2471\,
            I => \N__2431\
        );

    \I__269\ : IoInMux
    port map (
            O => \N__2470\,
            I => \N__2428\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2467\,
            I => \N__2423\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2464\,
            I => \N__2418\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2461\,
            I => \N__2418\
        );

    \I__265\ : IoInMux
    port map (
            O => \N__2460\,
            I => \N__2415\
        );

    \I__264\ : IoInMux
    port map (
            O => \N__2459\,
            I => \N__2412\
        );

    \I__263\ : Span4Mux_s3_v
    port map (
            O => \N__2454\,
            I => \N__2403\
        );

    \I__262\ : Span4Mux_s3_v
    port map (
            O => \N__2451\,
            I => \N__2400\
        );

    \I__261\ : IoSpan4Mux
    port map (
            O => \N__2440\,
            I => \N__2389\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2437\,
            I => \N__2389\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__2434\,
            I => \N__2389\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__2431\,
            I => \N__2389\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2428\,
            I => \N__2389\
        );

    \I__256\ : IoInMux
    port map (
            O => \N__2427\,
            I => \N__2386\
        );

    \I__255\ : IoInMux
    port map (
            O => \N__2426\,
            I => \N__2383\
        );

    \I__254\ : IoSpan4Mux
    port map (
            O => \N__2423\,
            I => \N__2374\
        );

    \I__253\ : IoSpan4Mux
    port map (
            O => \N__2418\,
            I => \N__2374\
        );

    \I__252\ : LocalMux
    port map (
            O => \N__2415\,
            I => \N__2374\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2412\,
            I => \N__2374\
        );

    \I__250\ : IoInMux
    port map (
            O => \N__2411\,
            I => \N__2371\
        );

    \I__249\ : IoInMux
    port map (
            O => \N__2410\,
            I => \N__2368\
        );

    \I__248\ : IoInMux
    port map (
            O => \N__2409\,
            I => \N__2365\
        );

    \I__247\ : IoInMux
    port map (
            O => \N__2408\,
            I => \N__2362\
        );

    \I__246\ : IoInMux
    port map (
            O => \N__2407\,
            I => \N__2359\
        );

    \I__245\ : IoInMux
    port map (
            O => \N__2406\,
            I => \N__2356\
        );

    \I__244\ : Span4Mux_v
    port map (
            O => \N__2403\,
            I => \N__2353\
        );

    \I__243\ : Span4Mux_v
    port map (
            O => \N__2400\,
            I => \N__2350\
        );

    \I__242\ : IoSpan4Mux
    port map (
            O => \N__2389\,
            I => \N__2343\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2386\,
            I => \N__2343\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__2383\,
            I => \N__2343\
        );

    \I__239\ : IoSpan4Mux
    port map (
            O => \N__2374\,
            I => \N__2332\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2371\,
            I => \N__2332\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__2368\,
            I => \N__2332\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2365\,
            I => \N__2332\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__2362\,
            I => \N__2332\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2359\,
            I => \N__2327\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__2356\,
            I => \N__2327\
        );

    \I__232\ : Sp12to4
    port map (
            O => \N__2353\,
            I => \N__2322\
        );

    \I__231\ : Sp12to4
    port map (
            O => \N__2350\,
            I => \N__2322\
        );

    \I__230\ : IoSpan4Mux
    port map (
            O => \N__2343\,
            I => \N__2317\
        );

    \I__229\ : IoSpan4Mux
    port map (
            O => \N__2332\,
            I => \N__2317\
        );

    \I__228\ : Span12Mux_s7_v
    port map (
            O => \N__2327\,
            I => \N__2312\
        );

    \I__227\ : Span12Mux_h
    port map (
            O => \N__2322\,
            I => \N__2312\
        );

    \I__226\ : Span4Mux_s3_h
    port map (
            O => \N__2317\,
            I => \N__2309\
        );

    \I__225\ : Span12Mux_v
    port map (
            O => \N__2312\,
            I => \N__2306\
        );

    \I__224\ : Span4Mux_h
    port map (
            O => \N__2309\,
            I => \N__2303\
        );

    \I__223\ : Odrv12
    port map (
            O => \N__2306\,
            I => \RnW_c_i_0\
        );

    \I__222\ : Odrv4
    port map (
            O => \N__2303\,
            I => \RnW_c_i_0\
        );

    \I__221\ : InMux
    port map (
            O => \N__2298\,
            I => \N__2295\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__2295\,
            I => \N__2292\
        );

    \I__219\ : Span12Mux_h
    port map (
            O => \N__2292\,
            I => \N__2289\
        );

    \I__218\ : Span12Mux_h
    port map (
            O => \N__2289\,
            I => \N__2286\
        );

    \I__217\ : Odrv12
    port map (
            O => \N__2286\,
            I => \D_UM_040_in_0\
        );

    \I__216\ : IoInMux
    port map (
            O => \N__2283\,
            I => \N__2279\
        );

    \I__215\ : CascadeMux
    port map (
            O => \N__2282\,
            I => \N__2276\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__2279\,
            I => \N__2273\
        );

    \I__213\ : InMux
    port map (
            O => \N__2276\,
            I => \N__2270\
        );

    \I__212\ : IoSpan4Mux
    port map (
            O => \N__2273\,
            I => \N__2267\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__2270\,
            I => \N__2264\
        );

    \I__210\ : Span4Mux_s2_h
    port map (
            O => \N__2267\,
            I => \N__2261\
        );

    \I__209\ : Span12Mux_v
    port map (
            O => \N__2264\,
            I => \N__2258\
        );

    \I__208\ : Sp12to4
    port map (
            O => \N__2261\,
            I => \N__2255\
        );

    \I__207\ : Span12Mux_v
    port map (
            O => \N__2258\,
            I => \N__2252\
        );

    \I__206\ : Span12Mux_h
    port map (
            O => \N__2255\,
            I => \N__2249\
        );

    \I__205\ : Span12Mux_h
    port map (
            O => \N__2252\,
            I => \N__2246\
        );

    \I__204\ : Span12Mux_h
    port map (
            O => \N__2249\,
            I => \N__2243\
        );

    \I__203\ : Odrv12
    port map (
            O => \N__2246\,
            I => \D_LL_040_in_0\
        );

    \I__202\ : Odrv12
    port map (
            O => \N__2243\,
            I => \D_LL_040_in_0\
        );

    \I__201\ : IoInMux
    port map (
            O => \N__2238\,
            I => \N__2235\
        );

    \I__200\ : LocalMux
    port map (
            O => \N__2235\,
            I => \N__2232\
        );

    \I__199\ : Span4Mux_s1_h
    port map (
            O => \N__2232\,
            I => \N__2229\
        );

    \I__198\ : Span4Mux_h
    port map (
            O => \N__2229\,
            I => \N__2226\
        );

    \I__197\ : Span4Mux_h
    port map (
            O => \N__2226\,
            I => \N__2223\
        );

    \I__196\ : Odrv4
    port map (
            O => \N__2223\,
            I => \un1_D_UM_040_0\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_5C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net\,
            I => \N__6227\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_2C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_2C_net\,
            I => \N__6231\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            I => \N__6224\
        );

    \INVU111_CYCLE_SM.LW_CYCLEC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.LW_CYCLEC_net\,
            I => \N__6225\
        );

    \INVU111_CYCLE_SM.CYCLE_STATE_0C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.CYCLE_STATE_0C_net\,
            I => \N__6228\
        );

    \INVU111_CYCLE_SM.TS_ENC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TS_ENC_net\,
            I => \N__6229\
        );

    \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            I => \N__6226\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            I => \N__6230\
        );

    \INVU111_CYCLE_SM.A_OUTC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.A_OUTC_net\,
            I => \N__6232\
        );

    \INVU111_CYCLE_SM.TA_ENC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TA_ENC_net\,
            I => \N__6233\
        );

    \INVU111_CYCLE_SM.TSnC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TSnC_net\,
            I => \N__6075\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__2637\,
            in1 => \N__7479\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \A_AMIGA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2607\,
            in1 => \N__7478\,
            in2 => \_gnd_net_\,
            in3 => \N__4134\,
            lcout => \A_AMIGA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__4363\,
            in1 => \N__5386\,
            in2 => \N__6445\,
            in3 => \N__2595\,
            lcout => \un1_D_LL_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RnW_c_sbtinv_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5981\,
            lcout => \RnW_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__2298\,
            in1 => \N__5352\,
            in2 => \N__2282\,
            in3 => \N__4409\,
            lcout => \un1_D_UM_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__5337\,
            in1 => \N__7113\,
            in2 => \N__3207\,
            in3 => \N__4452\,
            lcout => \un1_D_LM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__5368\,
            in1 => \N__3171\,
            in2 => \N__3149\,
            in3 => \N__4453\,
            lcout => \un1_D_UM_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__4449\,
            in1 => \N__5380\,
            in2 => \N__3093\,
            in3 => \N__3065\,
            lcout => \un1_D_UM_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_6_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__5387\,
            in1 => \N__3009\,
            in2 => \N__4554\,
            in3 => \N__2975\,
            lcout => \un1_D_UU_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__2909\,
            in1 => \N__5388\,
            in2 => \N__2880\,
            in3 => \N__4525\,
            lcout => \un1_D_UU_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__2838\,
            in1 => \N__5338\,
            in2 => \N__6776\,
            in3 => \N__4466\,
            lcout => \un1_D_LL_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__2801\,
            in1 => \N__5356\,
            in2 => \N__4560\,
            in3 => \N__2757\,
            lcout => \un1_D_UM_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__5373\,
            in1 => \N__2721\,
            in2 => \N__2696\,
            in3 => \N__4561\,
            lcout => \un1_D_UU_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__5374\,
            in1 => \N__6684\,
            in2 => \N__3588\,
            in3 => \N__4427\,
            lcout => \un1_D_LL_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__4503\,
            in1 => \N__5268\,
            in2 => \N__3549\,
            in3 => \N__3530\,
            lcout => \un1_D_UM_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__4504\,
            in1 => \N__5228\,
            in2 => \N__6540\,
            in3 => \N__3471\,
            lcout => \un1_D_LM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__3438\,
            in1 => \N__5309\,
            in2 => \N__6609\,
            in3 => \N__4539\,
            lcout => \un1_D_LM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__4562\,
            in1 => \N__5379\,
            in2 => \N__3405\,
            in3 => \N__3371\,
            lcout => \un1_D_UU_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__4341\,
            in1 => \N__5372\,
            in2 => \N__4104\,
            in3 => \N__3330\,
            lcout => \un1_D_LL_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TSn_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5601\,
            in2 => \_gnd_net_\,
            in3 => \N__5055\,
            lcout => \TSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TSnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__5307\,
            in1 => \N__3276\,
            in2 => \N__5544\,
            in3 => \N__4492\,
            lcout => \un1_D_LM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__3246\,
            in1 => \N__5308\,
            in2 => \N__4251\,
            in3 => \N__4526\,
            lcout => \un1_D_LM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__5344\,
            in1 => \N__4008\,
            in2 => \N__4566\,
            in3 => \N__3986\,
            lcout => \un1_D_UU_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__4559\,
            in1 => \N__5378\,
            in2 => \N__3927\,
            in3 => \N__3906\,
            lcout => \un1_D_UU_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__6051\,
            in1 => \N__5348\,
            in2 => \N__3846\,
            in3 => \N__4457\,
            lcout => \un1_D_LL_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_RNO_0_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5609\,
            lcout => \U111_CYCLE_SM.RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__5343\,
            in1 => \N__3801\,
            in2 => \N__3756\,
            in3 => \N__4558\,
            lcout => \un1_D_UM_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__5367\,
            in1 => \N__3711\,
            in2 => \N__6861\,
            in3 => \N__4439\,
            lcout => \un1_D_LL_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__4438\,
            in1 => \N__5366\,
            in2 => \N__6135\,
            in3 => \N__3672\,
            lcout => \un1_D_LL_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__5322\,
            in1 => \N__7038\,
            in2 => \N__3633\,
            in3 => \N__4481\,
            lcout => \un1_D_LL_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__5321\,
            in1 => \N__4188\,
            in2 => \N__7185\,
            in3 => \N__4480\,
            lcout => \un1_D_LM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7461\,
            in1 => \N__4059\,
            in2 => \_gnd_net_\,
            in3 => \N__4094\,
            lcout => \un1_D_UM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000011011100"
        )
    port map (
            in0 => \N__5680\,
            in1 => \N__6399\,
            in2 => \N__5445\,
            in3 => \N__6291\,
            lcout => \U111_CYCLE_SM.TA_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TA_ENC_net\,
            ce => 'H',
            sr => \N__4143\
        );

    \U111_CYCLE_SM.A_OUT_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5643\,
            in2 => \_gnd_net_\,
            in3 => \N__4110\,
            lcout => \U111_CYCLE_SM.A_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.A_OUTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_RNO_0_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001110"
        )
    port map (
            in0 => \N__4121\,
            in1 => \N__6392\,
            in2 => \N__5682\,
            in3 => \N__6284\,
            lcout => \U111_CYCLE_SM.A_OUT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6040\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            ce => \N__7272\,
            sr => \N__7243\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4081\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_6C_net\,
            ce => \N__7272\,
            sr => \N__7243\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010101010"
        )
    port map (
            in0 => \N__4050\,
            in1 => \N__5198\,
            in2 => \N__6951\,
            in3 => \N__4448\,
            lcout => \un1_D_LM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5540\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__7273\,
            sr => \N__7236\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4247\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__7273\,
            sr => \N__7236\
        );

    \CONSTANT_ONE_LUT4_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__5275\,
            in1 => \N__7335\,
            in2 => \N__4563\,
            in3 => \N__4938\,
            lcout => \un1_D_LM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011010000"
        )
    port map (
            in0 => \N__4450\,
            in1 => \N__5339\,
            in2 => \N__4899\,
            in3 => \N__4868\,
            lcout => \un1_D_UM_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__5340\,
            in1 => \N__4815\,
            in2 => \N__4796\,
            in3 => \N__4451\,
            lcout => \un1_D_UU_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__4565\,
            in1 => \N__5342\,
            in2 => \N__4724\,
            in3 => \N__4680\,
            lcout => \un1_D_UM_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__5341\,
            in1 => \N__4638\,
            in2 => \N__4613\,
            in3 => \N__4564\,
            lcout => \un1_D_UU_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4263\,
            in1 => \N__4240\,
            in2 => \_gnd_net_\,
            in3 => \N__7467\,
            lcout => \un1_D_UU_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5556\,
            in1 => \N__5527\,
            in2 => \_gnd_net_\,
            in3 => \N__7466\,
            lcout => \un1_D_UU_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_THRU_LUT4_0_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6090\,
            lcout => \GB_BUFFER_CLK40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_RNI1DSB_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__5444\,
            in1 => \N__6341\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM_TAn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__5010\,
            in1 => \N__5004\,
            in2 => \N__5644\,
            in3 => \N__5048\,
            lcout => \U111_CYCLE_SM.TS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TS_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI2RET_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100000111"
        )
    port map (
            in0 => \N__5093\,
            in1 => \N__5111\,
            in2 => \N__7460\,
            in3 => \N__5072\,
            lcout => \U111_CYCLE_SM.un1_LW_TRANS_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000000000"
        )
    port map (
            in0 => \N__5112\,
            in1 => \N__5094\,
            in2 => \N__5076\,
            in3 => \N__5047\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.un3_LW_CYCLE_START_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__7419\,
            in1 => \N__5631\,
            in2 => \N__5031\,
            in3 => \N__5679\,
            lcout => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TS_ENC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_1_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001101010000"
        )
    port map (
            in0 => \N__6283\,
            in1 => \N__5028\,
            in2 => \N__6398\,
            in3 => \N__6088\,
            lcout => \U111_CYCLE_SM.TS_EN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_0_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111011"
        )
    port map (
            in0 => \N__6087\,
            in1 => \N__6388\,
            in2 => \_gnd_net_\,
            in3 => \N__6282\,
            lcout => \U111_CYCLE_SM.N_69_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5678\,
            in1 => \N__6089\,
            in2 => \_gnd_net_\,
            in3 => \N__6393\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_91_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_0_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__5635\,
            in1 => \N__6342\,
            in2 => \N__6054\,
            in3 => \N__6288\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.CYCLE_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_1_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010000001000"
        )
    port map (
            in0 => \N__6289\,
            in1 => \N__5636\,
            in2 => \N__6350\,
            in3 => \N__6394\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.CYCLE_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001010"
        )
    port map (
            in0 => \N__6041\,
            in1 => \N__6015\,
            in2 => \N__7424\,
            in3 => \_gnd_net_\,
            lcout => \un1_D_UM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIFCLM_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6346\,
            in2 => \N__6290\,
            in3 => \N__6385\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1_0_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110101"
        )
    port map (
            in0 => \N__5645\,
            in1 => \_gnd_net_\,
            in2 => \N__5988\,
            in3 => \N__5904\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0\,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_RNI14FL1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGG4C2_0_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5691\,
            in3 => \N__5688\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5681\,
            in2 => \_gnd_net_\,
            in3 => \N__6280\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__5646\,
            in1 => \N__6243\,
            in2 => \N__6402\,
            in3 => \N__6387\,
            lcout => \U111_CYCLE_SM.LW_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.LW_CYCLEC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__6386\,
            in1 => \N__7383\,
            in2 => \N__6351\,
            in3 => \N__6281\,
            lcout => \U111_CYCLE_SM.LW_CYCLE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6854\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__7271\,
            sr => \N__7232\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6674\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__7271\,
            sr => \N__7232\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6533\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__7271\,
            sr => \N__7232\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6128\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__7271\,
            sr => \N__7232\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6777\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__7271\,
            sr => \N__7232\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6608\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__7271\,
            sr => \N__7232\
        );

    \GB_BUFFER_CLK80_THRU_LUT4_0_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6237\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_CLK80_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7425\,
            in1 => \N__6141\,
            in2 => \_gnd_net_\,
            in3 => \N__6127\,
            lcout => \un1_D_UM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6853\,
            in1 => \N__6810\,
            in2 => \_gnd_net_\,
            in3 => \N__7426\,
            lcout => \un1_D_UM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6766\,
            in1 => \N__6726\,
            in2 => \_gnd_net_\,
            in3 => \N__7463\,
            lcout => \un1_D_UM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6693\,
            in1 => \N__6662\,
            in2 => \_gnd_net_\,
            in3 => \N__7462\,
            lcout => \un1_D_UM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7465\,
            in1 => \N__6618\,
            in2 => \_gnd_net_\,
            in3 => \N__6595\,
            lcout => \un1_D_UU_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6526\,
            in1 => \N__7464\,
            in2 => \_gnd_net_\,
            in3 => \N__6495\,
            lcout => \un1_D_UU_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6447\,
            in1 => \N__6408\,
            in2 => \_gnd_net_\,
            in3 => \N__7423\,
            lcout => \un1_D_UM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6446\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_2C_net\,
            ce => \N__7274\,
            sr => \N__7244\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7034\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net\,
            ce => \N__7275\,
            sr => \N__7245\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7109\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net\,
            ce => \N__7275\,
            sr => \N__7245\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6950\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net\,
            ce => \N__7275\,
            sr => \N__7245\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7334\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net\,
            ce => \N__7275\,
            sr => \N__7245\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7178\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_5C_net\,
            ce => \N__7275\,
            sr => \N__7245\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7469\,
            in1 => \N__7194\,
            in2 => \_gnd_net_\,
            in3 => \N__7171\,
            lcout => \un1_D_UU_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7102\,
            in1 => \N__7068\,
            in2 => \_gnd_net_\,
            in3 => \N__7468\,
            lcout => \un1_D_UU_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7030\,
            in1 => \N__6990\,
            in2 => \_gnd_net_\,
            in3 => \N__7470\,
            lcout => \un1_D_UM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7471\,
            in1 => \N__6960\,
            in2 => \_gnd_net_\,
            in3 => \N__6946\,
            lcout => \un1_D_UU_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7472\,
            in1 => \N__7344\,
            in2 => \_gnd_net_\,
            in3 => \N__7327\,
            lcout => \un1_D_UU_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

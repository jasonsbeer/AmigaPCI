// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 23 2024 21:58:13

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    CMA,
    DRA,
    A,
    TSn,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    VBENn,
    CUMBEn,
    CLKRAM,
    C3,
    ASn,
    LDSn,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CASLn,
    RAMSPACEn,
    WEn,
    REGENn,
    DBRn,
    CLK40C,
    CLK40_IN,
    REGSPACEn,
    RAMENn,
    RASn,
    TACKn,
    C1);

    input [1:0] SIZ;
    output [10:0] CMA;
    input [9:0] DRA;
    input [20:0] A;
    input TSn;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    input C3;
    output ASn;
    output LDSn;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    input CASLn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    input DBRn;
    output CLK40C;
    input CLK40_IN;
    input REGSPACEn;
    output RAMENn;
    output RASn;
    output TACKn;
    input C1;

    wire N__10315;
    wire N__10314;
    wire N__10313;
    wire N__10306;
    wire N__10305;
    wire N__10304;
    wire N__10297;
    wire N__10296;
    wire N__10295;
    wire N__10288;
    wire N__10287;
    wire N__10286;
    wire N__10279;
    wire N__10278;
    wire N__10277;
    wire N__10270;
    wire N__10269;
    wire N__10268;
    wire N__10261;
    wire N__10260;
    wire N__10259;
    wire N__10252;
    wire N__10251;
    wire N__10250;
    wire N__10243;
    wire N__10242;
    wire N__10241;
    wire N__10234;
    wire N__10233;
    wire N__10232;
    wire N__10225;
    wire N__10224;
    wire N__10223;
    wire N__10216;
    wire N__10215;
    wire N__10214;
    wire N__10207;
    wire N__10206;
    wire N__10205;
    wire N__10198;
    wire N__10197;
    wire N__10196;
    wire N__10189;
    wire N__10188;
    wire N__10187;
    wire N__10180;
    wire N__10179;
    wire N__10178;
    wire N__10171;
    wire N__10170;
    wire N__10169;
    wire N__10162;
    wire N__10161;
    wire N__10160;
    wire N__10153;
    wire N__10152;
    wire N__10151;
    wire N__10144;
    wire N__10143;
    wire N__10142;
    wire N__10135;
    wire N__10134;
    wire N__10133;
    wire N__10126;
    wire N__10125;
    wire N__10124;
    wire N__10117;
    wire N__10116;
    wire N__10115;
    wire N__10108;
    wire N__10107;
    wire N__10106;
    wire N__10099;
    wire N__10098;
    wire N__10097;
    wire N__10090;
    wire N__10089;
    wire N__10088;
    wire N__10081;
    wire N__10080;
    wire N__10079;
    wire N__10072;
    wire N__10071;
    wire N__10070;
    wire N__10063;
    wire N__10062;
    wire N__10061;
    wire N__10054;
    wire N__10053;
    wire N__10052;
    wire N__10045;
    wire N__10044;
    wire N__10043;
    wire N__10036;
    wire N__10035;
    wire N__10034;
    wire N__10027;
    wire N__10026;
    wire N__10025;
    wire N__10018;
    wire N__10017;
    wire N__10016;
    wire N__10009;
    wire N__10008;
    wire N__10007;
    wire N__10000;
    wire N__9999;
    wire N__9998;
    wire N__9991;
    wire N__9990;
    wire N__9989;
    wire N__9982;
    wire N__9981;
    wire N__9980;
    wire N__9973;
    wire N__9972;
    wire N__9971;
    wire N__9964;
    wire N__9963;
    wire N__9962;
    wire N__9955;
    wire N__9954;
    wire N__9953;
    wire N__9946;
    wire N__9945;
    wire N__9944;
    wire N__9937;
    wire N__9936;
    wire N__9935;
    wire N__9928;
    wire N__9927;
    wire N__9926;
    wire N__9919;
    wire N__9918;
    wire N__9917;
    wire N__9910;
    wire N__9909;
    wire N__9908;
    wire N__9901;
    wire N__9900;
    wire N__9899;
    wire N__9892;
    wire N__9891;
    wire N__9890;
    wire N__9883;
    wire N__9882;
    wire N__9881;
    wire N__9874;
    wire N__9873;
    wire N__9872;
    wire N__9865;
    wire N__9864;
    wire N__9863;
    wire N__9856;
    wire N__9855;
    wire N__9854;
    wire N__9847;
    wire N__9846;
    wire N__9845;
    wire N__9838;
    wire N__9837;
    wire N__9836;
    wire N__9829;
    wire N__9828;
    wire N__9827;
    wire N__9820;
    wire N__9819;
    wire N__9818;
    wire N__9811;
    wire N__9810;
    wire N__9809;
    wire N__9802;
    wire N__9801;
    wire N__9800;
    wire N__9793;
    wire N__9792;
    wire N__9791;
    wire N__9784;
    wire N__9783;
    wire N__9782;
    wire N__9775;
    wire N__9774;
    wire N__9773;
    wire N__9766;
    wire N__9765;
    wire N__9764;
    wire N__9757;
    wire N__9756;
    wire N__9755;
    wire N__9748;
    wire N__9747;
    wire N__9746;
    wire N__9739;
    wire N__9738;
    wire N__9737;
    wire N__9730;
    wire N__9729;
    wire N__9728;
    wire N__9721;
    wire N__9720;
    wire N__9719;
    wire N__9712;
    wire N__9711;
    wire N__9710;
    wire N__9703;
    wire N__9702;
    wire N__9701;
    wire N__9694;
    wire N__9693;
    wire N__9692;
    wire N__9685;
    wire N__9684;
    wire N__9683;
    wire N__9676;
    wire N__9675;
    wire N__9674;
    wire N__9667;
    wire N__9666;
    wire N__9665;
    wire N__9658;
    wire N__9657;
    wire N__9656;
    wire N__9649;
    wire N__9648;
    wire N__9647;
    wire N__9640;
    wire N__9639;
    wire N__9638;
    wire N__9631;
    wire N__9630;
    wire N__9629;
    wire N__9622;
    wire N__9621;
    wire N__9620;
    wire N__9613;
    wire N__9612;
    wire N__9611;
    wire N__9604;
    wire N__9603;
    wire N__9602;
    wire N__9585;
    wire N__9582;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9569;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9555;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9543;
    wire N__9540;
    wire N__9537;
    wire N__9534;
    wire N__9533;
    wire N__9532;
    wire N__9531;
    wire N__9530;
    wire N__9529;
    wire N__9528;
    wire N__9527;
    wire N__9526;
    wire N__9525;
    wire N__9524;
    wire N__9523;
    wire N__9522;
    wire N__9521;
    wire N__9520;
    wire N__9519;
    wire N__9518;
    wire N__9517;
    wire N__9516;
    wire N__9515;
    wire N__9514;
    wire N__9513;
    wire N__9512;
    wire N__9511;
    wire N__9510;
    wire N__9507;
    wire N__9506;
    wire N__9505;
    wire N__9504;
    wire N__9503;
    wire N__9502;
    wire N__9501;
    wire N__9500;
    wire N__9499;
    wire N__9498;
    wire N__9497;
    wire N__9496;
    wire N__9495;
    wire N__9494;
    wire N__9493;
    wire N__9492;
    wire N__9491;
    wire N__9490;
    wire N__9489;
    wire N__9488;
    wire N__9487;
    wire N__9486;
    wire N__9485;
    wire N__9484;
    wire N__9483;
    wire N__9482;
    wire N__9481;
    wire N__9480;
    wire N__9479;
    wire N__9372;
    wire N__9369;
    wire N__9366;
    wire N__9365;
    wire N__9364;
    wire N__9363;
    wire N__9362;
    wire N__9361;
    wire N__9360;
    wire N__9359;
    wire N__9358;
    wire N__9357;
    wire N__9356;
    wire N__9355;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9326;
    wire N__9323;
    wire N__9322;
    wire N__9321;
    wire N__9320;
    wire N__9319;
    wire N__9318;
    wire N__9315;
    wire N__9314;
    wire N__9313;
    wire N__9312;
    wire N__9311;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9303;
    wire N__9302;
    wire N__9301;
    wire N__9298;
    wire N__9297;
    wire N__9296;
    wire N__9295;
    wire N__9294;
    wire N__9293;
    wire N__9292;
    wire N__9289;
    wire N__9286;
    wire N__9285;
    wire N__9284;
    wire N__9283;
    wire N__9280;
    wire N__9279;
    wire N__9278;
    wire N__9277;
    wire N__9276;
    wire N__9273;
    wire N__9272;
    wire N__9271;
    wire N__9270;
    wire N__9269;
    wire N__9268;
    wire N__9267;
    wire N__9266;
    wire N__9265;
    wire N__9264;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9147;
    wire N__9144;
    wire N__9141;
    wire N__9138;
    wire N__9135;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9095;
    wire N__9092;
    wire N__9091;
    wire N__9088;
    wire N__9085;
    wire N__9082;
    wire N__9081;
    wire N__9080;
    wire N__9077;
    wire N__9072;
    wire N__9069;
    wire N__9066;
    wire N__9065;
    wire N__9064;
    wire N__9057;
    wire N__9054;
    wire N__9051;
    wire N__9048;
    wire N__9045;
    wire N__9042;
    wire N__9037;
    wire N__9030;
    wire N__9029;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9021;
    wire N__9020;
    wire N__9019;
    wire N__9018;
    wire N__9017;
    wire N__9014;
    wire N__9009;
    wire N__9006;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8994;
    wire N__8991;
    wire N__8988;
    wire N__8987;
    wire N__8986;
    wire N__8981;
    wire N__8976;
    wire N__8971;
    wire N__8968;
    wire N__8967;
    wire N__8964;
    wire N__8963;
    wire N__8962;
    wire N__8959;
    wire N__8956;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8937;
    wire N__8922;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8900;
    wire N__8899;
    wire N__8898;
    wire N__8897;
    wire N__8896;
    wire N__8895;
    wire N__8892;
    wire N__8891;
    wire N__8890;
    wire N__8887;
    wire N__8882;
    wire N__8881;
    wire N__8878;
    wire N__8875;
    wire N__8872;
    wire N__8869;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8854;
    wire N__8851;
    wire N__8840;
    wire N__8837;
    wire N__8836;
    wire N__8835;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8774;
    wire N__8771;
    wire N__8770;
    wire N__8769;
    wire N__8766;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8736;
    wire N__8731;
    wire N__8728;
    wire N__8725;
    wire N__8718;
    wire N__8717;
    wire N__8716;
    wire N__8715;
    wire N__8714;
    wire N__8711;
    wire N__8710;
    wire N__8709;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8698;
    wire N__8695;
    wire N__8694;
    wire N__8691;
    wire N__8688;
    wire N__8685;
    wire N__8682;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8645;
    wire N__8642;
    wire N__8641;
    wire N__8640;
    wire N__8637;
    wire N__8634;
    wire N__8633;
    wire N__8630;
    wire N__8625;
    wire N__8620;
    wire N__8617;
    wire N__8616;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8591;
    wire N__8586;
    wire N__8583;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8538;
    wire N__8537;
    wire N__8536;
    wire N__8535;
    wire N__8532;
    wire N__8529;
    wire N__8524;
    wire N__8517;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8463;
    wire N__8460;
    wire N__8457;
    wire N__8454;
    wire N__8451;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8380;
    wire N__8379;
    wire N__8378;
    wire N__8377;
    wire N__8376;
    wire N__8375;
    wire N__8374;
    wire N__8373;
    wire N__8372;
    wire N__8371;
    wire N__8370;
    wire N__8369;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8357;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8346;
    wire N__8345;
    wire N__8344;
    wire N__8343;
    wire N__8340;
    wire N__8335;
    wire N__8330;
    wire N__8325;
    wire N__8324;
    wire N__8323;
    wire N__8320;
    wire N__8315;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8298;
    wire N__8295;
    wire N__8288;
    wire N__8285;
    wire N__8278;
    wire N__8273;
    wire N__8272;
    wire N__8267;
    wire N__8264;
    wire N__8253;
    wire N__8250;
    wire N__8241;
    wire N__8240;
    wire N__8239;
    wire N__8236;
    wire N__8233;
    wire N__8228;
    wire N__8225;
    wire N__8220;
    wire N__8215;
    wire N__8202;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8187;
    wire N__8184;
    wire N__8181;
    wire N__8178;
    wire N__8175;
    wire N__8172;
    wire N__8169;
    wire N__8168;
    wire N__8165;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8139;
    wire N__8136;
    wire N__8133;
    wire N__8130;
    wire N__8127;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8094;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8082;
    wire N__8079;
    wire N__8076;
    wire N__8073;
    wire N__8070;
    wire N__8067;
    wire N__8064;
    wire N__8061;
    wire N__8058;
    wire N__8055;
    wire N__8052;
    wire N__8049;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8019;
    wire N__8016;
    wire N__8013;
    wire N__8010;
    wire N__8007;
    wire N__8004;
    wire N__8003;
    wire N__8002;
    wire N__8001;
    wire N__8000;
    wire N__7999;
    wire N__7998;
    wire N__7997;
    wire N__7996;
    wire N__7995;
    wire N__7994;
    wire N__7993;
    wire N__7992;
    wire N__7991;
    wire N__7988;
    wire N__7983;
    wire N__7982;
    wire N__7981;
    wire N__7978;
    wire N__7973;
    wire N__7968;
    wire N__7967;
    wire N__7966;
    wire N__7965;
    wire N__7964;
    wire N__7963;
    wire N__7962;
    wire N__7959;
    wire N__7956;
    wire N__7949;
    wire N__7946;
    wire N__7941;
    wire N__7938;
    wire N__7937;
    wire N__7934;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7912;
    wire N__7909;
    wire N__7906;
    wire N__7901;
    wire N__7900;
    wire N__7899;
    wire N__7898;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7885;
    wire N__7876;
    wire N__7873;
    wire N__7868;
    wire N__7861;
    wire N__7858;
    wire N__7851;
    wire N__7846;
    wire N__7841;
    wire N__7838;
    wire N__7833;
    wire N__7830;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7812;
    wire N__7809;
    wire N__7806;
    wire N__7803;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7788;
    wire N__7785;
    wire N__7782;
    wire N__7779;
    wire N__7776;
    wire N__7773;
    wire N__7770;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7749;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7737;
    wire N__7734;
    wire N__7731;
    wire N__7728;
    wire N__7725;
    wire N__7722;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7710;
    wire N__7707;
    wire N__7704;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7683;
    wire N__7680;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7668;
    wire N__7665;
    wire N__7662;
    wire N__7659;
    wire N__7656;
    wire N__7653;
    wire N__7650;
    wire N__7647;
    wire N__7644;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7614;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7602;
    wire N__7599;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7581;
    wire N__7578;
    wire N__7575;
    wire N__7572;
    wire N__7569;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7551;
    wire N__7548;
    wire N__7545;
    wire N__7542;
    wire N__7539;
    wire N__7536;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7517;
    wire N__7514;
    wire N__7511;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7452;
    wire N__7449;
    wire N__7446;
    wire N__7443;
    wire N__7440;
    wire N__7437;
    wire N__7434;
    wire N__7431;
    wire N__7428;
    wire N__7425;
    wire N__7422;
    wire N__7419;
    wire N__7416;
    wire N__7413;
    wire N__7410;
    wire N__7409;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7392;
    wire N__7389;
    wire N__7386;
    wire N__7385;
    wire N__7382;
    wire N__7379;
    wire N__7378;
    wire N__7373;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7344;
    wire N__7341;
    wire N__7338;
    wire N__7337;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7299;
    wire N__7296;
    wire N__7293;
    wire N__7290;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7278;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7266;
    wire N__7265;
    wire N__7262;
    wire N__7259;
    wire N__7254;
    wire N__7251;
    wire N__7248;
    wire N__7245;
    wire N__7242;
    wire N__7239;
    wire N__7238;
    wire N__7235;
    wire N__7234;
    wire N__7233;
    wire N__7230;
    wire N__7229;
    wire N__7226;
    wire N__7225;
    wire N__7218;
    wire N__7215;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7194;
    wire N__7185;
    wire N__7184;
    wire N__7181;
    wire N__7178;
    wire N__7175;
    wire N__7172;
    wire N__7171;
    wire N__7170;
    wire N__7167;
    wire N__7164;
    wire N__7161;
    wire N__7158;
    wire N__7149;
    wire N__7146;
    wire N__7143;
    wire N__7140;
    wire N__7137;
    wire N__7134;
    wire N__7131;
    wire N__7128;
    wire N__7125;
    wire N__7122;
    wire N__7119;
    wire N__7116;
    wire N__7113;
    wire N__7110;
    wire N__7107;
    wire N__7104;
    wire N__7101;
    wire N__7098;
    wire N__7095;
    wire N__7092;
    wire N__7089;
    wire N__7086;
    wire N__7083;
    wire N__7080;
    wire N__7077;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7047;
    wire N__7044;
    wire N__7041;
    wire N__7038;
    wire N__7035;
    wire N__7032;
    wire N__7029;
    wire N__7026;
    wire N__7023;
    wire N__7020;
    wire N__7017;
    wire N__7014;
    wire N__7011;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6993;
    wire N__6990;
    wire N__6989;
    wire N__6986;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6972;
    wire N__6971;
    wire N__6968;
    wire N__6965;
    wire N__6964;
    wire N__6963;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6953;
    wire N__6950;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6938;
    wire N__6935;
    wire N__6932;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6911;
    wire N__6906;
    wire N__6905;
    wire N__6904;
    wire N__6903;
    wire N__6900;
    wire N__6897;
    wire N__6896;
    wire N__6895;
    wire N__6894;
    wire N__6891;
    wire N__6888;
    wire N__6883;
    wire N__6878;
    wire N__6875;
    wire N__6864;
    wire N__6861;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6831;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6819;
    wire N__6818;
    wire N__6817;
    wire N__6816;
    wire N__6813;
    wire N__6806;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6780;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6768;
    wire N__6765;
    wire N__6762;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6744;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6732;
    wire N__6729;
    wire N__6726;
    wire N__6723;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6708;
    wire N__6705;
    wire N__6702;
    wire N__6699;
    wire N__6696;
    wire N__6693;
    wire N__6690;
    wire N__6687;
    wire N__6684;
    wire N__6681;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6642;
    wire N__6639;
    wire N__6636;
    wire N__6633;
    wire N__6630;
    wire N__6627;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6603;
    wire N__6600;
    wire N__6597;
    wire N__6594;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6569;
    wire N__6564;
    wire N__6563;
    wire N__6562;
    wire N__6561;
    wire N__6558;
    wire N__6555;
    wire N__6550;
    wire N__6543;
    wire N__6540;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6528;
    wire N__6525;
    wire N__6522;
    wire N__6519;
    wire N__6516;
    wire N__6513;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6501;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6493;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6474;
    wire N__6471;
    wire N__6462;
    wire N__6459;
    wire N__6456;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6441;
    wire N__6438;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6420;
    wire N__6419;
    wire N__6414;
    wire N__6411;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6387;
    wire N__6384;
    wire N__6383;
    wire N__6380;
    wire N__6377;
    wire N__6372;
    wire N__6369;
    wire N__6366;
    wire N__6363;
    wire N__6360;
    wire N__6357;
    wire N__6354;
    wire N__6351;
    wire N__6348;
    wire N__6345;
    wire N__6342;
    wire N__6339;
    wire N__6336;
    wire N__6333;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6317;
    wire N__6316;
    wire N__6313;
    wire N__6308;
    wire N__6303;
    wire N__6300;
    wire N__6297;
    wire N__6294;
    wire N__6293;
    wire N__6292;
    wire N__6291;
    wire N__6288;
    wire N__6281;
    wire N__6276;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6264;
    wire N__6263;
    wire N__6260;
    wire N__6259;
    wire N__6258;
    wire N__6257;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6244;
    wire N__6243;
    wire N__6242;
    wire N__6241;
    wire N__6240;
    wire N__6239;
    wire N__6238;
    wire N__6237;
    wire N__6234;
    wire N__6233;
    wire N__6230;
    wire N__6227;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6207;
    wire N__6204;
    wire N__6197;
    wire N__6180;
    wire N__6179;
    wire N__6178;
    wire N__6175;
    wire N__6170;
    wire N__6167;
    wire N__6162;
    wire N__6161;
    wire N__6158;
    wire N__6157;
    wire N__6156;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6129;
    wire N__6128;
    wire N__6127;
    wire N__6126;
    wire N__6125;
    wire N__6120;
    wire N__6117;
    wire N__6112;
    wire N__6109;
    wire N__6104;
    wire N__6101;
    wire N__6096;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6072;
    wire N__6071;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6048;
    wire N__6047;
    wire N__6046;
    wire N__6043;
    wire N__6038;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6018;
    wire N__6015;
    wire N__6012;
    wire N__6011;
    wire N__6010;
    wire N__6009;
    wire N__6008;
    wire N__6007;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5992;
    wire N__5987;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5966;
    wire N__5965;
    wire N__5962;
    wire N__5961;
    wire N__5958;
    wire N__5955;
    wire N__5954;
    wire N__5953;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5941;
    wire N__5938;
    wire N__5933;
    wire N__5922;
    wire N__5919;
    wire N__5918;
    wire N__5917;
    wire N__5916;
    wire N__5915;
    wire N__5914;
    wire N__5913;
    wire N__5912;
    wire N__5911;
    wire N__5906;
    wire N__5903;
    wire N__5902;
    wire N__5901;
    wire N__5898;
    wire N__5897;
    wire N__5894;
    wire N__5889;
    wire N__5888;
    wire N__5887;
    wire N__5886;
    wire N__5881;
    wire N__5878;
    wire N__5875;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5857;
    wire N__5854;
    wire N__5851;
    wire N__5848;
    wire N__5841;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5808;
    wire N__5805;
    wire N__5802;
    wire N__5801;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5756;
    wire N__5751;
    wire N__5748;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5736;
    wire N__5735;
    wire N__5734;
    wire N__5733;
    wire N__5732;
    wire N__5731;
    wire N__5730;
    wire N__5727;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5713;
    wire N__5710;
    wire N__5697;
    wire N__5694;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5682;
    wire N__5681;
    wire N__5680;
    wire N__5679;
    wire N__5678;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5670;
    wire N__5667;
    wire N__5664;
    wire N__5661;
    wire N__5656;
    wire N__5651;
    wire N__5648;
    wire N__5637;
    wire N__5634;
    wire N__5633;
    wire N__5632;
    wire N__5631;
    wire N__5630;
    wire N__5629;
    wire N__5624;
    wire N__5621;
    wire N__5620;
    wire N__5619;
    wire N__5618;
    wire N__5617;
    wire N__5616;
    wire N__5615;
    wire N__5614;
    wire N__5613;
    wire N__5612;
    wire N__5611;
    wire N__5608;
    wire N__5603;
    wire N__5598;
    wire N__5595;
    wire N__5590;
    wire N__5583;
    wire N__5574;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5532;
    wire N__5529;
    wire N__5526;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5504;
    wire N__5499;
    wire N__5496;
    wire N__5495;
    wire N__5494;
    wire N__5493;
    wire N__5490;
    wire N__5483;
    wire N__5478;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5423;
    wire N__5422;
    wire N__5419;
    wire N__5414;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5397;
    wire N__5396;
    wire N__5395;
    wire N__5394;
    wire N__5391;
    wire N__5388;
    wire N__5385;
    wire N__5382;
    wire N__5373;
    wire N__5370;
    wire N__5367;
    wire N__5366;
    wire N__5365;
    wire N__5362;
    wire N__5357;
    wire N__5354;
    wire N__5349;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5337;
    wire N__5334;
    wire N__5331;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5319;
    wire N__5316;
    wire N__5315;
    wire N__5314;
    wire N__5313;
    wire N__5310;
    wire N__5305;
    wire N__5302;
    wire N__5295;
    wire N__5292;
    wire N__5291;
    wire N__5290;
    wire N__5287;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5264;
    wire N__5263;
    wire N__5262;
    wire N__5255;
    wire N__5252;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5234;
    wire N__5233;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5222;
    wire N__5221;
    wire N__5214;
    wire N__5211;
    wire N__5206;
    wire N__5199;
    wire N__5196;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5184;
    wire N__5183;
    wire N__5182;
    wire N__5181;
    wire N__5178;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5137;
    wire N__5134;
    wire N__5129;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5110;
    wire N__5107;
    wire N__5102;
    wire N__5097;
    wire N__5096;
    wire N__5095;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5079;
    wire N__5076;
    wire N__5073;
    wire N__5072;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5064;
    wire N__5061;
    wire N__5056;
    wire N__5051;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5030;
    wire N__5025;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5008;
    wire N__5005;
    wire N__5002;
    wire N__4999;
    wire N__4996;
    wire N__4993;
    wire N__4990;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4923;
    wire N__4920;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4899;
    wire N__4898;
    wire N__4895;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4885;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4869;
    wire N__4868;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4854;
    wire N__4851;
    wire N__4848;
    wire N__4845;
    wire N__4842;
    wire N__4839;
    wire N__4836;
    wire N__4833;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4800;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4785;
    wire N__4784;
    wire N__4781;
    wire N__4778;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4752;
    wire N__4751;
    wire N__4750;
    wire N__4749;
    wire N__4748;
    wire N__4745;
    wire N__4736;
    wire N__4731;
    wire N__4730;
    wire N__4725;
    wire N__4722;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4712;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4695;
    wire N__4692;
    wire N__4689;
    wire N__4686;
    wire N__4683;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4673;
    wire N__4672;
    wire N__4671;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4656;
    wire N__4653;
    wire N__4650;
    wire N__4647;
    wire N__4638;
    wire N__4635;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4608;
    wire N__4605;
    wire N__4602;
    wire N__4599;
    wire N__4596;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4584;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4560;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4548;
    wire N__4547;
    wire N__4546;
    wire N__4545;
    wire N__4544;
    wire N__4541;
    wire N__4532;
    wire N__4527;
    wire N__4524;
    wire N__4523;
    wire N__4522;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4512;
    wire N__4511;
    wire N__4510;
    wire N__4505;
    wire N__4496;
    wire N__4491;
    wire N__4490;
    wire N__4489;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4473;
    wire N__4470;
    wire N__4469;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4459;
    wire N__4452;
    wire N__4449;
    wire N__4446;
    wire N__4445;
    wire N__4444;
    wire N__4443;
    wire N__4442;
    wire N__4437;
    wire N__4430;
    wire N__4425;
    wire N__4424;
    wire N__4421;
    wire N__4420;
    wire N__4417;
    wire N__4416;
    wire N__4415;
    wire N__4410;
    wire N__4403;
    wire N__4398;
    wire N__4395;
    wire N__4392;
    wire N__4389;
    wire N__4388;
    wire N__4387;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4372;
    wire N__4369;
    wire N__4362;
    wire N__4359;
    wire N__4356;
    wire N__4353;
    wire N__4350;
    wire N__4347;
    wire N__4344;
    wire N__4341;
    wire N__4340;
    wire N__4339;
    wire N__4332;
    wire N__4329;
    wire N__4326;
    wire N__4325;
    wire N__4320;
    wire N__4317;
    wire N__4316;
    wire N__4315;
    wire N__4314;
    wire N__4311;
    wire N__4308;
    wire N__4303;
    wire N__4300;
    wire N__4293;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4281;
    wire N__4278;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4270;
    wire N__4269;
    wire N__4264;
    wire N__4259;
    wire N__4254;
    wire N__4251;
    wire N__4250;
    wire N__4245;
    wire N__4242;
    wire N__4241;
    wire N__4240;
    wire N__4239;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4227;
    wire N__4224;
    wire N__4215;
    wire N__4214;
    wire N__4211;
    wire N__4210;
    wire N__4209;
    wire N__4206;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4192;
    wire N__4185;
    wire N__4184;
    wire N__4183;
    wire N__4178;
    wire N__4175;
    wire N__4170;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4155;
    wire N__4152;
    wire N__4151;
    wire N__4150;
    wire N__4147;
    wire N__4142;
    wire N__4137;
    wire N__4134;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4104;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4092;
    wire N__4089;
    wire N__4086;
    wire N__4083;
    wire N__4080;
    wire N__4077;
    wire N__4074;
    wire N__4071;
    wire N__4068;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4049;
    wire N__4048;
    wire N__4045;
    wire N__4038;
    wire N__4035;
    wire N__4034;
    wire N__4029;
    wire N__4026;
    wire N__4023;
    wire N__4020;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4008;
    wire N__4005;
    wire N__4002;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3990;
    wire N__3987;
    wire N__3984;
    wire N__3981;
    wire N__3980;
    wire N__3977;
    wire N__3976;
    wire N__3973;
    wire N__3970;
    wire N__3967;
    wire N__3964;
    wire N__3957;
    wire N__3956;
    wire N__3953;
    wire N__3952;
    wire N__3949;
    wire N__3948;
    wire N__3945;
    wire N__3942;
    wire N__3939;
    wire N__3936;
    wire N__3927;
    wire N__3924;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3916;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire N__3897;
    wire N__3894;
    wire N__3891;
    wire N__3888;
    wire N__3885;
    wire N__3882;
    wire N__3879;
    wire N__3876;
    wire N__3873;
    wire N__3870;
    wire N__3867;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3855;
    wire N__3852;
    wire N__3851;
    wire N__3848;
    wire N__3845;
    wire N__3840;
    wire N__3837;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3825;
    wire N__3822;
    wire N__3821;
    wire N__3818;
    wire N__3815;
    wire N__3812;
    wire N__3807;
    wire N__3804;
    wire N__3801;
    wire N__3798;
    wire N__3795;
    wire N__3792;
    wire N__3789;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3759;
    wire N__3756;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3744;
    wire N__3741;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3717;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3702;
    wire N__3699;
    wire N__3696;
    wire N__3693;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_OUT_i_i;
    wire CLK40_OUT_i_i;
    wire REGSPACEn_c;
    wire \U712_REG_SM.un6_REG_CYCLE_START_cascade_ ;
    wire \U712_REG_SM.REG_CYCLE_GOZ0 ;
    wire C1_c;
    wire C3_c;
    wire \U712_CHIP_RAM.REFRESH_r_1_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ;
    wire bfn_7_7_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH6lto2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire C1_c_g;
    wire \U712_REG_SM.STATE_COUNTZ1Z_0 ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.N_168_0_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_2 ;
    wire \U712_REG_SM.N_175_cascade_ ;
    wire \U712_REG_SM.N_171_0 ;
    wire \U712_REG_SM.N_194_cascade_ ;
    wire \U712_REG_SM.N_169_0 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_1 ;
    wire \U712_REG_SM.N_170_0_cascade_ ;
    wire \U712_REG_SM.N_174_cascade_ ;
    wire \U712_REG_SM.N_162_0_cascade_ ;
    wire \U712_REG_SM.N_172_0 ;
    wire \U712_REG_SM.N_162_0 ;
    wire \U712_REG_SM.N_195 ;
    wire \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_ ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_2 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_163_0 ;
    wire \U712_REG_SM.N_194 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_6 ;
    wire ASn_c;
    wire \U712_REG_SM.N_186_0 ;
    wire N_510_i;
    wire VBENn_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_ ;
    wire \U712_CHIP_RAM.N_43_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_1_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_2_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_a2_0_4_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_a2_0_1 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_cascade_ ;
    wire TACK_OUTn;
    wire \U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1 ;
    wire \U712_REG_SM.DS_EN_7_0 ;
    wire \U712_REG_SM.N_187 ;
    wire \U712_REG_SM.N_157_0 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_2 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.N_159_0 ;
    wire \U712_REG_SM.N_159_0_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_4 ;
    wire \U712_REG_SM.N_165_0 ;
    wire \U712_REG_SM.N_165_0_cascade_ ;
    wire \U712_REG_SM.N_170_0 ;
    wire \U712_REG_SM.N_173_0 ;
    wire \U712_REG_SM.LDS_OUT_2_0_0 ;
    wire \U712_REG_SM.UDS_OUT_2_0_0 ;
    wire \U712_CHIP_RAM.N_105_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_i_1_1_cascade_ ;
    wire \U712_CHIP_RAM.N_105 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER17_1 ;
    wire \U712_CHIP_RAM.N_50_cascade_ ;
    wire \U712_CHIP_RAM.N_43 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_tz_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ;
    wire \U712_CHIP_RAM.N_68 ;
    wire \U712_CHIP_RAM.N_98 ;
    wire \U712_CHIP_RAM.N_55_cascade_ ;
    wire \U712_CHIP_RAM.N_57_cascade_ ;
    wire \U712_CHIP_RAM.N_92_cascade_ ;
    wire \U712_CHIP_RAM.N_44 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.BANK0_0_sqmuxa_3 ;
    wire \U712_CHIP_RAM.N_106_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_cascade_ ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.N_100 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0 ;
    wire \U712_CHIP_RAM.CPU_TACK_6 ;
    wire RAMSPACEn_c;
    wire \U712_CHIP_RAM.un6_CPU_CYCLE_START_cascade_ ;
    wire TSn_c;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire \U712_CYCLE_TERM.N_49 ;
    wire REG_TACK;
    wire CPU_TACKm;
    wire \U712_CYCLE_TERM.TACK_EN6_0_cascade_ ;
    wire CLK40_OUT_i;
    wire \U712_CYCLE_TERM.TACK_STATEZ1Z_2 ;
    wire DBDIR_c;
    wire DRDDIR_0_i;
    wire CLMBEn_c;
    wire \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1 ;
    wire \U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1_cascade_ ;
    wire CLLBEn_c;
    wire DBENn_c;
    wire \U712_REG_SM.STATE_COUNTZ0Z_5 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_3 ;
    wire \U712_REG_SM.N_167_0 ;
    wire \U712_BYTE_ENABLE.LLBE_0 ;
    wire \U712_BYTE_ENABLE.LMBE_0 ;
    wire SIZ_c_0;
    wire A_c_1;
    wire A_c_0;
    wire SIZ_c_1;
    wire A_c_11;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_ ;
    wire A_c_4;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.N_78_cascade_ ;
    wire \U712_CHIP_RAM.N_76_cascade_ ;
    wire \U712_CHIP_RAM.N_58 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c2 ;
    wire \U712_CHIP_RAM.N_46 ;
    wire \U712_CHIP_RAM.N_77 ;
    wire \U712_CHIP_RAM.N_99 ;
    wire \U712_CHIP_RAM.N_99_cascade_ ;
    wire \U712_CHIP_RAM.N_79 ;
    wire \U712_CHIP_RAM.N_93_1 ;
    wire \U712_CHIP_RAM.N_52 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_54 ;
    wire \U712_CHIP_RAM.N_50 ;
    wire \U712_CHIP_RAM.N_54_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire \U712_CHIP_RAM.REFRESH_CYCLE_START_2_2_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.REFRESH_CYCLE_0_sqmuxa_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_0 ;
    wire \U712_CHIP_RAM.REFRESH_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_70_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.N_106 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER53_3_0 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.N_40 ;
    wire \U712_CHIP_RAM.N_40_cascade_ ;
    wire \U712_CHIP_RAM.N_51 ;
    wire \U712_CHIP_RAM.N_59 ;
    wire \U712_CHIP_RAM.N_59_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CYCLE_TERM.N_45_0_0_en ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ;
    wire U712_REG_SM_DBR_SYNC_1;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0 ;
    wire DBRn_c;
    wire U712_REG_SM_DBR_SYNC_0;
    wire \U712_BYTE_ENABLE.UMBE_0 ;
    wire CUMBEn_c;
    wire \U712_BYTE_ENABLE.UUBE_0 ;
    wire \U712_BYTE_ENABLE.un3_CUMBEnZ0Z_0 ;
    wire CUUBEn_c;
    wire \U712_REG_SM.LDS_OUTZ0 ;
    wire U712_REG_SM_un1_LDSn_i;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.N_33 ;
    wire CMA_c_2;
    wire A_c_13;
    wire A_c_6;
    wire \U712_CHIP_RAM.N_35_cascade_ ;
    wire CMA_c_4;
    wire A_c_12;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_ ;
    wire A_c_5;
    wire \U712_CHIP_RAM.N_34 ;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire A_c_10;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_ ;
    wire A_c_3;
    wire \U712_CHIP_RAM.DBENn_7_0_a2_0 ;
    wire AWEn_c;
    wire RnW_c;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0 ;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire TACK_EN_i_ess;
    wire \U712_CYCLE_TERM.N_45_0_0_en_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESS4 ;
    wire CASLn_c;
    wire CASUn_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_REG_SM.UDS_OUTZ0 ;
    wire \U712_REG_SM.DS_ENZ0 ;
    wire U712_REG_SM_un1_UDSn_i;
    wire DMA_CYCLEm;
    wire REG_CYCLEm;
    wire DRDENn_c;
    wire CONSTANT_ONE_NET;
    wire A_c_14;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_5_cascade_ ;
    wire A_c_7;
    wire \U712_CHIP_RAM.un1_CMA31_0_i ;
    wire DRA_c_4;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.N_32 ;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire RESETn_c;
    wire RESETn_c_i;
    wire CMA_c_0;
    wire \U712_CHIP_RAM.N_36 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire A_c_9;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_ ;
    wire A_c_2;
    wire \U712_CHIP_RAM.N_31 ;
    wire A_c_17;
    wire CMA_c_8;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.CMA_5_0_8 ;
    wire A_c_19;
    wire CMA_c_9;
    wire A_c_15;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_6 ;
    wire A_c_8;
    wire \U712_CHIP_RAM.N_37 ;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire CPU_CYCLEm;
    wire A_c_16;
    wire \U712_CHIP_RAM.CMA_5_3_ns_1_7_cascade_ ;
    wire A_c_18;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire DRA_c_7;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_1;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.N_38 ;
    wire CMA_c_7;
    wire CMA_c_10;
    wire \U712_CHIP_RAM.un1_CMA31_0_i_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ;
    wire WEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ;
    wire RASn_c;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire CRCSn_c;
    wire RAS1n_c;
    wire RAS0n_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire _gnd_net_;
    wire CLK80_OUT;
    wire RESETn_c_i_g;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_OUT_i),
            .REFERENCECLK(N__3711),
            .RESETB(N__7125),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_OUT),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__10315),
            .DIN(N__10314),
            .DOUT(N__10313),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__10315),
            .PADOUT(N__10314),
            .PADIN(N__10313),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5436),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__10306),
            .DIN(N__10305),
            .DOUT(N__10304),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__10306),
            .PADOUT(N__10305),
            .PADIN(N__10304),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__10297),
            .DIN(N__10296),
            .DOUT(N__10295),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__10297),
            .PADOUT(N__10296),
            .PADIN(N__10295),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8568),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__10288),
            .DIN(N__10287),
            .DOUT(N__10286),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__10288),
            .PADOUT(N__10287),
            .PADIN(N__10286),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4983),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__10279),
            .DIN(N__10278),
            .DOUT(N__10277),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__10279),
            .PADOUT(N__10278),
            .PADIN(N__10277),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__10270),
            .DIN(N__10269),
            .DOUT(N__10268),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__10270),
            .PADOUT(N__10269),
            .PADIN(N__10268),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__10261),
            .DIN(N__10260),
            .DOUT(N__10259),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__10261),
            .PADOUT(N__10260),
            .PADIN(N__10259),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__10252),
            .DIN(N__10251),
            .DOUT(N__10250),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__10252),
            .PADOUT(N__10251),
            .PADIN(N__10250),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__10243),
            .DIN(N__10242),
            .DOUT(N__10241),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__10243),
            .PADOUT(N__10242),
            .PADIN(N__10241),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__10234),
            .DIN(N__10233),
            .DOUT(N__10232),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__10234),
            .PADOUT(N__10233),
            .PADIN(N__10232),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__10225),
            .DIN(N__10224),
            .DOUT(N__10223),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__10225),
            .PADOUT(N__10224),
            .PADIN(N__10223),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9129),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMENn_obuf_iopad (
            .OE(N__10216),
            .DIN(N__10215),
            .DOUT(N__10214),
            .PACKAGEPIN(RAMENn));
    defparam RAMENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RAMENn_obuf_preio (
            .PADOEN(N__10216),
            .PADOUT(N__10215),
            .PADIN(N__10214),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6989),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__10207),
            .DIN(N__10206),
            .DOUT(N__10205),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__10207),
            .PADOUT(N__10206),
            .PADIN(N__10205),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__10198),
            .DIN(N__10197),
            .DOUT(N__10196),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__10198),
            .PADOUT(N__10197),
            .PADIN(N__10196),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__10189),
            .DIN(N__10188),
            .DOUT(N__10187),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__10189),
            .PADOUT(N__10188),
            .PADIN(N__10187),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4077),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__10180),
            .DIN(N__10179),
            .DOUT(N__10178),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__10180),
            .PADOUT(N__10179),
            .PADIN(N__10178),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__10171),
            .DIN(N__10170),
            .DOUT(N__10169),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__10171),
            .PADOUT(N__10170),
            .PADIN(N__10169),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__10162),
            .DIN(N__10161),
            .DOUT(N__10160),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__10162),
            .PADOUT(N__10161),
            .PADIN(N__10160),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7803),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__10153),
            .DIN(N__10152),
            .DOUT(N__10151),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__10153),
            .PADOUT(N__10152),
            .PADIN(N__10151),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__10144),
            .DIN(N__10143),
            .DOUT(N__10142),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__10144),
            .PADOUT(N__10143),
            .PADIN(N__10142),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8517),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__10135),
            .DIN(N__10134),
            .DOUT(N__10133),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__10135),
            .PADOUT(N__10134),
            .PADIN(N__10133),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__10126),
            .DIN(N__10125),
            .DOUT(N__10124),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__10126),
            .PADOUT(N__10125),
            .PADIN(N__10124),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__10117),
            .DIN(N__10116),
            .DOUT(N__10115),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__10117),
            .PADOUT(N__10116),
            .PADIN(N__10115),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__10108),
            .DIN(N__10107),
            .DOUT(N__10106),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__10108),
            .PADOUT(N__10107),
            .PADIN(N__10106),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__10099),
            .DIN(N__10098),
            .DOUT(N__10097),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__10099),
            .PADOUT(N__10098),
            .PADIN(N__10097),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__10090),
            .DIN(N__10089),
            .DOUT(N__10088),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__10090),
            .PADOUT(N__10089),
            .PADIN(N__10088),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__10081),
            .DIN(N__10080),
            .DOUT(N__10079),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__10081),
            .PADOUT(N__10080),
            .PADIN(N__10079),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__10072),
            .DIN(N__10071),
            .DOUT(N__10070),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__10072),
            .PADOUT(N__10071),
            .PADIN(N__10070),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__10063),
            .DIN(N__10062),
            .DOUT(N__10061),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__10063),
            .PADOUT(N__10062),
            .PADIN(N__10061),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__10054),
            .DIN(N__10053),
            .DOUT(N__10052),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__10054),
            .PADOUT(N__10053),
            .PADIN(N__10052),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7650),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__10045),
            .DIN(N__10044),
            .DOUT(N__10043),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__10045),
            .PADOUT(N__10044),
            .PADIN(N__10043),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__10036),
            .DIN(N__10035),
            .DOUT(N__10034),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__10036),
            .PADOUT(N__10035),
            .PADIN(N__10034),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__10027),
            .DIN(N__10026),
            .DOUT(N__10025),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__10027),
            .PADOUT(N__10026),
            .PADIN(N__10025),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__10018),
            .DIN(N__10017),
            .DOUT(N__10016),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__10018),
            .PADOUT(N__10017),
            .PADIN(N__10016),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_obuf_iopad (
            .OE(N__10009),
            .DIN(N__10008),
            .DOUT(N__10007),
            .PACKAGEPIN(CLK40C));
    defparam CLK40C_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_obuf_preio (
            .PADOEN(N__10009),
            .PADOUT(N__10008),
            .PADIN(N__10007),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3789),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__10000),
            .DIN(N__9999),
            .DOUT(N__9998),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__10000),
            .PADOUT(N__9999),
            .PADIN(N__9998),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6372),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__9991),
            .DIN(N__9990),
            .DOUT(N__9989),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__9991),
            .PADOUT(N__9990),
            .PADIN(N__9989),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__9982),
            .DIN(N__9981),
            .DOUT(N__9980),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__9982),
            .PADOUT(N__9981),
            .PADIN(N__9980),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8793),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__9973),
            .DIN(N__9972),
            .DOUT(N__9971),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__9973),
            .PADOUT(N__9972),
            .PADIN(N__9971),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__9964),
            .DIN(N__9963),
            .DOUT(N__9962),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__9964),
            .PADOUT(N__9963),
            .PADIN(N__9962),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__9955),
            .DIN(N__9954),
            .DOUT(N__9953),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__9955),
            .PADOUT(N__9954),
            .PADIN(N__9953),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3804),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__9946),
            .DIN(N__9945),
            .DOUT(N__9944),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__9946),
            .PADOUT(N__9945),
            .PADIN(N__9944),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__9937),
            .DIN(N__9936),
            .DOUT(N__9935),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__9937),
            .PADOUT(N__9936),
            .PADIN(N__9935),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4137),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__9928),
            .DIN(N__9927),
            .DOUT(N__9926),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__9928),
            .PADOUT(N__9927),
            .PADIN(N__9926),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6348),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__9919),
            .DIN(N__9918),
            .DOUT(N__9917),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__9919),
            .PADOUT(N__9918),
            .PADIN(N__9917),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__9910),
            .DIN(N__9909),
            .DOUT(N__9908),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__9910),
            .PADOUT(N__9909),
            .PADIN(N__9908),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam A_ibuf_0_iopad.PULLUP=1'b1;
    IO_PAD A_ibuf_0_iopad (
            .OE(N__9901),
            .DIN(N__9900),
            .DOUT(N__9899),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__9901),
            .PADOUT(N__9900),
            .PADIN(N__9899),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__9892),
            .DIN(N__9891),
            .DOUT(N__9890),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__9892),
            .PADOUT(N__9891),
            .PADIN(N__9890),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9108),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__9883),
            .DIN(N__9882),
            .DOUT(N__9881),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__9883),
            .PADOUT(N__9882),
            .PADIN(N__9881),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__9874),
            .DIN(N__9873),
            .DOUT(N__9872),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__9874),
            .PADOUT(N__9873),
            .PADIN(N__9872),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6702),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__9865),
            .DIN(N__9864),
            .DOUT(N__9863),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__9865),
            .PADOUT(N__9864),
            .PADIN(N__9863),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7149),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__9856),
            .DIN(N__9855),
            .DOUT(N__9854),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__9856),
            .PADOUT(N__9855),
            .PADIN(N__9854),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5457),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__9847),
            .DIN(N__9846),
            .DOUT(N__9845),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__9847),
            .PADOUT(N__9846),
            .PADIN(N__9845),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7590),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__9838),
            .DIN(N__9837),
            .DOUT(N__9836),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__9838),
            .PADOUT(N__9837),
            .PADIN(N__9836),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4133),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__9829),
            .DIN(N__9828),
            .DOUT(N__9827),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__9829),
            .PADOUT(N__9828),
            .PADIN(N__9827),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__9820),
            .DIN(N__9819),
            .DOUT(N__9818),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__9820),
            .PADOUT(N__9819),
            .PADIN(N__9818),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__9811),
            .DIN(N__9810),
            .DOUT(N__9809),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__9811),
            .PADOUT(N__9810),
            .PADIN(N__9809),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4959),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__9802),
            .DIN(N__9801),
            .DOUT(N__9800),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__9802),
            .PADOUT(N__9801),
            .PADIN(N__9800),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8922),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__9793),
            .DIN(N__9792),
            .DOUT(N__9791),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__9793),
            .PADOUT(N__9792),
            .PADIN(N__9791),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5022),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__9784),
            .DIN(N__9783),
            .DOUT(N__9782),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__9784),
            .PADOUT(N__9783),
            .PADIN(N__9782),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6456),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__9775),
            .DIN(N__9774),
            .DOUT(N__9773),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__9775),
            .PADOUT(N__9774),
            .PADIN(N__9773),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__9766),
            .DIN(N__9765),
            .DOUT(N__9764),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__9766),
            .PADOUT(N__9765),
            .PADIN(N__9764),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__9757),
            .DIN(N__9756),
            .DOUT(N__9755),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__9757),
            .PADOUT(N__9756),
            .PADIN(N__9755),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__9748),
            .DIN(N__9747),
            .DOUT(N__9746),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__9748),
            .PADOUT(N__9747),
            .PADIN(N__9746),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__9739),
            .DIN(N__9738),
            .DOUT(N__9737),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__9739),
            .PADOUT(N__9738),
            .PADIN(N__9737),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7437),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__9730),
            .DIN(N__9729),
            .DOUT(N__9728),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__9730),
            .PADOUT(N__9729),
            .PADIN(N__9728),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__9721),
            .DIN(N__9720),
            .DOUT(N__9719),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__9721),
            .PADOUT(N__9720),
            .PADIN(N__9719),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6411),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__9712),
            .DIN(N__9711),
            .DOUT(N__9710),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__9712),
            .PADOUT(N__9711),
            .PADIN(N__9710),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4089),
            .DIN0(),
            .DOUT0(N__4608),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__9703),
            .DIN(N__9702),
            .DOUT(N__9701),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__9703),
            .PADOUT(N__9702),
            .PADIN(N__9701),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6759),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__9694),
            .DIN(N__9693),
            .DOUT(N__9692),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__9694),
            .PADOUT(N__9693),
            .PADIN(N__9692),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__9685),
            .DIN(N__9684),
            .DOUT(N__9683),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__9685),
            .PADOUT(N__9684),
            .PADIN(N__9683),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__9676),
            .DIN(N__9675),
            .DOUT(N__9674),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__9676),
            .PADOUT(N__9675),
            .PADIN(N__9674),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7671),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__9667),
            .DIN(N__9666),
            .DOUT(N__9665),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__9667),
            .PADOUT(N__9666),
            .PADIN(N__9665),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__9658),
            .DIN(N__9657),
            .DOUT(N__9656),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__9658),
            .PADOUT(N__9657),
            .PADIN(N__9656),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__9649),
            .DIN(N__9648),
            .DOUT(N__9647),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__9649),
            .PADOUT(N__9648),
            .PADIN(N__9647),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__9640),
            .DIN(N__9639),
            .DOUT(N__9638),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__9640),
            .PADOUT(N__9639),
            .PADIN(N__9638),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__9631),
            .DIN(N__9630),
            .DOUT(N__9629),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__9631),
            .PADOUT(N__9630),
            .PADIN(N__9629),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7779),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__9622),
            .DIN(N__9621),
            .DOUT(N__9620),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__9622),
            .PADOUT(N__9621),
            .PADIN(N__9620),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7254),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__9613),
            .DIN(N__9612),
            .DOUT(N__9611),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__9613),
            .PADOUT(N__9612),
            .PADIN(N__9611),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4926),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__9604),
            .DIN(N__9603),
            .DOUT(N__9602),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__9604),
            .PADOUT(N__9603),
            .PADIN(N__9602),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2276 (
            .O(N__9585),
            .I(N__9582));
    LocalMux I__2275 (
            .O(N__9582),
            .I(N__9578));
    InMux I__2274 (
            .O(N__9581),
            .I(N__9575));
    Span4Mux_v I__2273 (
            .O(N__9578),
            .I(N__9572));
    LocalMux I__2272 (
            .O(N__9575),
            .I(N__9569));
    Span4Mux_h I__2271 (
            .O(N__9572),
            .I(N__9564));
    Span4Mux_v I__2270 (
            .O(N__9569),
            .I(N__9564));
    Sp12to4 I__2269 (
            .O(N__9564),
            .I(N__9561));
    Span12Mux_h I__2268 (
            .O(N__9561),
            .I(N__9558));
    Odrv12 I__2267 (
            .O(N__9558),
            .I(RAS0n_c));
    InMux I__2266 (
            .O(N__9555),
            .I(N__9551));
    InMux I__2265 (
            .O(N__9554),
            .I(N__9548));
    LocalMux I__2264 (
            .O(N__9551),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    LocalMux I__2263 (
            .O(N__9548),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2262 (
            .O(N__9543),
            .I(N__9540));
    LocalMux I__2261 (
            .O(N__9540),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__2260 (
            .O(N__9537),
            .I(N__9534));
    LocalMux I__2259 (
            .O(N__9534),
            .I(N__9507));
    ClkMux I__2258 (
            .O(N__9533),
            .I(N__9372));
    ClkMux I__2257 (
            .O(N__9532),
            .I(N__9372));
    ClkMux I__2256 (
            .O(N__9531),
            .I(N__9372));
    ClkMux I__2255 (
            .O(N__9530),
            .I(N__9372));
    ClkMux I__2254 (
            .O(N__9529),
            .I(N__9372));
    ClkMux I__2253 (
            .O(N__9528),
            .I(N__9372));
    ClkMux I__2252 (
            .O(N__9527),
            .I(N__9372));
    ClkMux I__2251 (
            .O(N__9526),
            .I(N__9372));
    ClkMux I__2250 (
            .O(N__9525),
            .I(N__9372));
    ClkMux I__2249 (
            .O(N__9524),
            .I(N__9372));
    ClkMux I__2248 (
            .O(N__9523),
            .I(N__9372));
    ClkMux I__2247 (
            .O(N__9522),
            .I(N__9372));
    ClkMux I__2246 (
            .O(N__9521),
            .I(N__9372));
    ClkMux I__2245 (
            .O(N__9520),
            .I(N__9372));
    ClkMux I__2244 (
            .O(N__9519),
            .I(N__9372));
    ClkMux I__2243 (
            .O(N__9518),
            .I(N__9372));
    ClkMux I__2242 (
            .O(N__9517),
            .I(N__9372));
    ClkMux I__2241 (
            .O(N__9516),
            .I(N__9372));
    ClkMux I__2240 (
            .O(N__9515),
            .I(N__9372));
    ClkMux I__2239 (
            .O(N__9514),
            .I(N__9372));
    ClkMux I__2238 (
            .O(N__9513),
            .I(N__9372));
    ClkMux I__2237 (
            .O(N__9512),
            .I(N__9372));
    ClkMux I__2236 (
            .O(N__9511),
            .I(N__9372));
    ClkMux I__2235 (
            .O(N__9510),
            .I(N__9372));
    Glb2LocalMux I__2234 (
            .O(N__9507),
            .I(N__9372));
    ClkMux I__2233 (
            .O(N__9506),
            .I(N__9372));
    ClkMux I__2232 (
            .O(N__9505),
            .I(N__9372));
    ClkMux I__2231 (
            .O(N__9504),
            .I(N__9372));
    ClkMux I__2230 (
            .O(N__9503),
            .I(N__9372));
    ClkMux I__2229 (
            .O(N__9502),
            .I(N__9372));
    ClkMux I__2228 (
            .O(N__9501),
            .I(N__9372));
    ClkMux I__2227 (
            .O(N__9500),
            .I(N__9372));
    ClkMux I__2226 (
            .O(N__9499),
            .I(N__9372));
    ClkMux I__2225 (
            .O(N__9498),
            .I(N__9372));
    ClkMux I__2224 (
            .O(N__9497),
            .I(N__9372));
    ClkMux I__2223 (
            .O(N__9496),
            .I(N__9372));
    ClkMux I__2222 (
            .O(N__9495),
            .I(N__9372));
    ClkMux I__2221 (
            .O(N__9494),
            .I(N__9372));
    ClkMux I__2220 (
            .O(N__9493),
            .I(N__9372));
    ClkMux I__2219 (
            .O(N__9492),
            .I(N__9372));
    ClkMux I__2218 (
            .O(N__9491),
            .I(N__9372));
    ClkMux I__2217 (
            .O(N__9490),
            .I(N__9372));
    ClkMux I__2216 (
            .O(N__9489),
            .I(N__9372));
    ClkMux I__2215 (
            .O(N__9488),
            .I(N__9372));
    ClkMux I__2214 (
            .O(N__9487),
            .I(N__9372));
    ClkMux I__2213 (
            .O(N__9486),
            .I(N__9372));
    ClkMux I__2212 (
            .O(N__9485),
            .I(N__9372));
    ClkMux I__2211 (
            .O(N__9484),
            .I(N__9372));
    ClkMux I__2210 (
            .O(N__9483),
            .I(N__9372));
    ClkMux I__2209 (
            .O(N__9482),
            .I(N__9372));
    ClkMux I__2208 (
            .O(N__9481),
            .I(N__9372));
    ClkMux I__2207 (
            .O(N__9480),
            .I(N__9372));
    ClkMux I__2206 (
            .O(N__9479),
            .I(N__9372));
    GlobalMux I__2205 (
            .O(N__9372),
            .I(CLK80_OUT));
    CascadeMux I__2204 (
            .O(N__9369),
            .I(N__9366));
    InMux I__2203 (
            .O(N__9366),
            .I(N__9346));
    InMux I__2202 (
            .O(N__9365),
            .I(N__9346));
    InMux I__2201 (
            .O(N__9364),
            .I(N__9346));
    InMux I__2200 (
            .O(N__9363),
            .I(N__9346));
    InMux I__2199 (
            .O(N__9362),
            .I(N__9343));
    InMux I__2198 (
            .O(N__9361),
            .I(N__9340));
    InMux I__2197 (
            .O(N__9360),
            .I(N__9337));
    InMux I__2196 (
            .O(N__9359),
            .I(N__9334));
    InMux I__2195 (
            .O(N__9358),
            .I(N__9331));
    InMux I__2194 (
            .O(N__9357),
            .I(N__9326));
    InMux I__2193 (
            .O(N__9356),
            .I(N__9326));
    InMux I__2192 (
            .O(N__9355),
            .I(N__9323));
    LocalMux I__2191 (
            .O(N__9346),
            .I(N__9315));
    LocalMux I__2190 (
            .O(N__9343),
            .I(N__9307));
    LocalMux I__2189 (
            .O(N__9340),
            .I(N__9304));
    LocalMux I__2188 (
            .O(N__9337),
            .I(N__9298));
    LocalMux I__2187 (
            .O(N__9334),
            .I(N__9289));
    LocalMux I__2186 (
            .O(N__9331),
            .I(N__9286));
    LocalMux I__2185 (
            .O(N__9326),
            .I(N__9280));
    LocalMux I__2184 (
            .O(N__9323),
            .I(N__9273));
    SRMux I__2183 (
            .O(N__9322),
            .I(N__9177));
    SRMux I__2182 (
            .O(N__9321),
            .I(N__9177));
    SRMux I__2181 (
            .O(N__9320),
            .I(N__9177));
    SRMux I__2180 (
            .O(N__9319),
            .I(N__9177));
    SRMux I__2179 (
            .O(N__9318),
            .I(N__9177));
    Glb2LocalMux I__2178 (
            .O(N__9315),
            .I(N__9177));
    SRMux I__2177 (
            .O(N__9314),
            .I(N__9177));
    SRMux I__2176 (
            .O(N__9313),
            .I(N__9177));
    SRMux I__2175 (
            .O(N__9312),
            .I(N__9177));
    SRMux I__2174 (
            .O(N__9311),
            .I(N__9177));
    SRMux I__2173 (
            .O(N__9310),
            .I(N__9177));
    Glb2LocalMux I__2172 (
            .O(N__9307),
            .I(N__9177));
    Glb2LocalMux I__2171 (
            .O(N__9304),
            .I(N__9177));
    SRMux I__2170 (
            .O(N__9303),
            .I(N__9177));
    SRMux I__2169 (
            .O(N__9302),
            .I(N__9177));
    SRMux I__2168 (
            .O(N__9301),
            .I(N__9177));
    Glb2LocalMux I__2167 (
            .O(N__9298),
            .I(N__9177));
    SRMux I__2166 (
            .O(N__9297),
            .I(N__9177));
    SRMux I__2165 (
            .O(N__9296),
            .I(N__9177));
    SRMux I__2164 (
            .O(N__9295),
            .I(N__9177));
    SRMux I__2163 (
            .O(N__9294),
            .I(N__9177));
    SRMux I__2162 (
            .O(N__9293),
            .I(N__9177));
    SRMux I__2161 (
            .O(N__9292),
            .I(N__9177));
    Glb2LocalMux I__2160 (
            .O(N__9289),
            .I(N__9177));
    Glb2LocalMux I__2159 (
            .O(N__9286),
            .I(N__9177));
    SRMux I__2158 (
            .O(N__9285),
            .I(N__9177));
    SRMux I__2157 (
            .O(N__9284),
            .I(N__9177));
    SRMux I__2156 (
            .O(N__9283),
            .I(N__9177));
    Glb2LocalMux I__2155 (
            .O(N__9280),
            .I(N__9177));
    SRMux I__2154 (
            .O(N__9279),
            .I(N__9177));
    SRMux I__2153 (
            .O(N__9278),
            .I(N__9177));
    SRMux I__2152 (
            .O(N__9277),
            .I(N__9177));
    SRMux I__2151 (
            .O(N__9276),
            .I(N__9177));
    Glb2LocalMux I__2150 (
            .O(N__9273),
            .I(N__9177));
    SRMux I__2149 (
            .O(N__9272),
            .I(N__9177));
    SRMux I__2148 (
            .O(N__9271),
            .I(N__9177));
    SRMux I__2147 (
            .O(N__9270),
            .I(N__9177));
    SRMux I__2146 (
            .O(N__9269),
            .I(N__9177));
    SRMux I__2145 (
            .O(N__9268),
            .I(N__9177));
    SRMux I__2144 (
            .O(N__9267),
            .I(N__9177));
    SRMux I__2143 (
            .O(N__9266),
            .I(N__9177));
    SRMux I__2142 (
            .O(N__9265),
            .I(N__9177));
    SRMux I__2141 (
            .O(N__9264),
            .I(N__9177));
    GlobalMux I__2140 (
            .O(N__9177),
            .I(N__9174));
    gio2CtrlBuf I__2139 (
            .O(N__9174),
            .I(RESETn_c_i_g));
    InMux I__2138 (
            .O(N__9171),
            .I(N__9168));
    LocalMux I__2137 (
            .O(N__9168),
            .I(N__9164));
    InMux I__2136 (
            .O(N__9167),
            .I(N__9161));
    Span4Mux_h I__2135 (
            .O(N__9164),
            .I(N__9156));
    LocalMux I__2134 (
            .O(N__9161),
            .I(N__9156));
    Span4Mux_h I__2133 (
            .O(N__9156),
            .I(N__9153));
    Sp12to4 I__2132 (
            .O(N__9153),
            .I(N__9150));
    Span12Mux_v I__2131 (
            .O(N__9150),
            .I(N__9147));
    Odrv12 I__2130 (
            .O(N__9147),
            .I(DRA_c_1));
    InMux I__2129 (
            .O(N__9144),
            .I(N__9141));
    LocalMux I__2128 (
            .O(N__9141),
            .I(N__9138));
    Odrv4 I__2127 (
            .O(N__9138),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__2126 (
            .O(N__9135),
            .I(N__9132));
    LocalMux I__2125 (
            .O(N__9132),
            .I(\U712_CHIP_RAM.N_38 ));
    IoInMux I__2124 (
            .O(N__9129),
            .I(N__9126));
    LocalMux I__2123 (
            .O(N__9126),
            .I(N__9123));
    IoSpan4Mux I__2122 (
            .O(N__9123),
            .I(N__9120));
    Sp12to4 I__2121 (
            .O(N__9120),
            .I(N__9117));
    Span12Mux_s1_h I__2120 (
            .O(N__9117),
            .I(N__9114));
    Span12Mux_h I__2119 (
            .O(N__9114),
            .I(N__9111));
    Odrv12 I__2118 (
            .O(N__9111),
            .I(CMA_c_7));
    IoInMux I__2117 (
            .O(N__9108),
            .I(N__9105));
    LocalMux I__2116 (
            .O(N__9105),
            .I(N__9102));
    Span12Mux_s9_v I__2115 (
            .O(N__9102),
            .I(N__9099));
    Odrv12 I__2114 (
            .O(N__9099),
            .I(CMA_c_10));
    CEMux I__2113 (
            .O(N__9096),
            .I(N__9092));
    CEMux I__2112 (
            .O(N__9095),
            .I(N__9088));
    LocalMux I__2111 (
            .O(N__9092),
            .I(N__9085));
    CEMux I__2110 (
            .O(N__9091),
            .I(N__9082));
    LocalMux I__2109 (
            .O(N__9088),
            .I(N__9077));
    Span4Mux_h I__2108 (
            .O(N__9085),
            .I(N__9072));
    LocalMux I__2107 (
            .O(N__9082),
            .I(N__9072));
    CEMux I__2106 (
            .O(N__9081),
            .I(N__9069));
    CEMux I__2105 (
            .O(N__9080),
            .I(N__9066));
    Span4Mux_v I__2104 (
            .O(N__9077),
            .I(N__9057));
    Span4Mux_v I__2103 (
            .O(N__9072),
            .I(N__9057));
    LocalMux I__2102 (
            .O(N__9069),
            .I(N__9057));
    LocalMux I__2101 (
            .O(N__9066),
            .I(N__9054));
    CEMux I__2100 (
            .O(N__9065),
            .I(N__9051));
    CEMux I__2099 (
            .O(N__9064),
            .I(N__9048));
    Span4Mux_h I__2098 (
            .O(N__9057),
            .I(N__9045));
    Span4Mux_h I__2097 (
            .O(N__9054),
            .I(N__9042));
    LocalMux I__2096 (
            .O(N__9051),
            .I(N__9037));
    LocalMux I__2095 (
            .O(N__9048),
            .I(N__9037));
    Odrv4 I__2094 (
            .O(N__9045),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv4 I__2093 (
            .O(N__9042),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    Odrv12 I__2092 (
            .O(N__9037),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i_0 ));
    CascadeMux I__2091 (
            .O(N__9030),
            .I(N__9025));
    CascadeMux I__2090 (
            .O(N__9029),
            .I(N__9022));
    InMux I__2089 (
            .O(N__9028),
            .I(N__9014));
    InMux I__2088 (
            .O(N__9025),
            .I(N__9009));
    InMux I__2087 (
            .O(N__9022),
            .I(N__9009));
    CascadeMux I__2086 (
            .O(N__9021),
            .I(N__9006));
    InMux I__2085 (
            .O(N__9020),
            .I(N__9002));
    InMux I__2084 (
            .O(N__9019),
            .I(N__8999));
    InMux I__2083 (
            .O(N__9018),
            .I(N__8994));
    InMux I__2082 (
            .O(N__9017),
            .I(N__8994));
    LocalMux I__2081 (
            .O(N__9014),
            .I(N__8991));
    LocalMux I__2080 (
            .O(N__9009),
            .I(N__8988));
    InMux I__2079 (
            .O(N__9006),
            .I(N__8981));
    InMux I__2078 (
            .O(N__9005),
            .I(N__8981));
    LocalMux I__2077 (
            .O(N__9002),
            .I(N__8976));
    LocalMux I__2076 (
            .O(N__8999),
            .I(N__8976));
    LocalMux I__2075 (
            .O(N__8994),
            .I(N__8971));
    Span4Mux_h I__2074 (
            .O(N__8991),
            .I(N__8971));
    Span4Mux_h I__2073 (
            .O(N__8988),
            .I(N__8968));
    CascadeMux I__2072 (
            .O(N__8987),
            .I(N__8964));
    InMux I__2071 (
            .O(N__8986),
            .I(N__8959));
    LocalMux I__2070 (
            .O(N__8981),
            .I(N__8956));
    Span4Mux_v I__2069 (
            .O(N__8976),
            .I(N__8951));
    Span4Mux_v I__2068 (
            .O(N__8971),
            .I(N__8951));
    Span4Mux_h I__2067 (
            .O(N__8968),
            .I(N__8948));
    InMux I__2066 (
            .O(N__8967),
            .I(N__8945));
    InMux I__2065 (
            .O(N__8964),
            .I(N__8942));
    InMux I__2064 (
            .O(N__8963),
            .I(N__8937));
    InMux I__2063 (
            .O(N__8962),
            .I(N__8937));
    LocalMux I__2062 (
            .O(N__8959),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    Odrv4 I__2061 (
            .O(N__8956),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    Odrv4 I__2060 (
            .O(N__8951),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    Odrv4 I__2059 (
            .O(N__8948),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    LocalMux I__2058 (
            .O(N__8945),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    LocalMux I__2057 (
            .O(N__8942),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    LocalMux I__2056 (
            .O(N__8937),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ));
    IoInMux I__2055 (
            .O(N__8922),
            .I(N__8919));
    LocalMux I__2054 (
            .O(N__8919),
            .I(N__8916));
    Span4Mux_s3_h I__2053 (
            .O(N__8916),
            .I(N__8913));
    Span4Mux_v I__2052 (
            .O(N__8913),
            .I(N__8910));
    Span4Mux_h I__2051 (
            .O(N__8910),
            .I(N__8907));
    Span4Mux_h I__2050 (
            .O(N__8907),
            .I(N__8904));
    Odrv4 I__2049 (
            .O(N__8904),
            .I(WEn_c));
    InMux I__2048 (
            .O(N__8901),
            .I(N__8892));
    InMux I__2047 (
            .O(N__8900),
            .I(N__8887));
    InMux I__2046 (
            .O(N__8899),
            .I(N__8882));
    InMux I__2045 (
            .O(N__8898),
            .I(N__8882));
    InMux I__2044 (
            .O(N__8897),
            .I(N__8878));
    InMux I__2043 (
            .O(N__8896),
            .I(N__8875));
    InMux I__2042 (
            .O(N__8895),
            .I(N__8872));
    LocalMux I__2041 (
            .O(N__8892),
            .I(N__8869));
    InMux I__2040 (
            .O(N__8891),
            .I(N__8864));
    InMux I__2039 (
            .O(N__8890),
            .I(N__8864));
    LocalMux I__2038 (
            .O(N__8887),
            .I(N__8861));
    LocalMux I__2037 (
            .O(N__8882),
            .I(N__8858));
    CascadeMux I__2036 (
            .O(N__8881),
            .I(N__8855));
    LocalMux I__2035 (
            .O(N__8878),
            .I(N__8851));
    LocalMux I__2034 (
            .O(N__8875),
            .I(N__8840));
    LocalMux I__2033 (
            .O(N__8872),
            .I(N__8840));
    Span4Mux_v I__2032 (
            .O(N__8869),
            .I(N__8840));
    LocalMux I__2031 (
            .O(N__8864),
            .I(N__8840));
    Span4Mux_h I__2030 (
            .O(N__8861),
            .I(N__8840));
    Span4Mux_h I__2029 (
            .O(N__8858),
            .I(N__8837));
    InMux I__2028 (
            .O(N__8855),
            .I(N__8831));
    InMux I__2027 (
            .O(N__8854),
            .I(N__8828));
    Span4Mux_v I__2026 (
            .O(N__8851),
            .I(N__8825));
    Span4Mux_h I__2025 (
            .O(N__8840),
            .I(N__8822));
    Span4Mux_h I__2024 (
            .O(N__8837),
            .I(N__8819));
    InMux I__2023 (
            .O(N__8836),
            .I(N__8816));
    InMux I__2022 (
            .O(N__8835),
            .I(N__8813));
    InMux I__2021 (
            .O(N__8834),
            .I(N__8810));
    LocalMux I__2020 (
            .O(N__8831),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    LocalMux I__2019 (
            .O(N__8828),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv4 I__2018 (
            .O(N__8825),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv4 I__2017 (
            .O(N__8822),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    Odrv4 I__2016 (
            .O(N__8819),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    LocalMux I__2015 (
            .O(N__8816),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    LocalMux I__2014 (
            .O(N__8813),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    LocalMux I__2013 (
            .O(N__8810),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ));
    IoInMux I__2012 (
            .O(N__8793),
            .I(N__8790));
    LocalMux I__2011 (
            .O(N__8790),
            .I(N__8787));
    Span4Mux_s3_v I__2010 (
            .O(N__8787),
            .I(N__8784));
    Span4Mux_v I__2009 (
            .O(N__8784),
            .I(N__8781));
    Span4Mux_h I__2008 (
            .O(N__8781),
            .I(N__8778));
    Odrv4 I__2007 (
            .O(N__8778),
            .I(RASn_c));
    CEMux I__2006 (
            .O(N__8775),
            .I(N__8771));
    CEMux I__2005 (
            .O(N__8774),
            .I(N__8766));
    LocalMux I__2004 (
            .O(N__8771),
            .I(N__8762));
    CEMux I__2003 (
            .O(N__8770),
            .I(N__8759));
    CEMux I__2002 (
            .O(N__8769),
            .I(N__8756));
    LocalMux I__2001 (
            .O(N__8766),
            .I(N__8753));
    CEMux I__2000 (
            .O(N__8765),
            .I(N__8750));
    Span4Mux_v I__1999 (
            .O(N__8762),
            .I(N__8747));
    LocalMux I__1998 (
            .O(N__8759),
            .I(N__8744));
    LocalMux I__1997 (
            .O(N__8756),
            .I(N__8741));
    Span4Mux_v I__1996 (
            .O(N__8753),
            .I(N__8736));
    LocalMux I__1995 (
            .O(N__8750),
            .I(N__8736));
    Span4Mux_h I__1994 (
            .O(N__8747),
            .I(N__8731));
    Span4Mux_v I__1993 (
            .O(N__8744),
            .I(N__8731));
    Span4Mux_h I__1992 (
            .O(N__8741),
            .I(N__8728));
    Span4Mux_h I__1991 (
            .O(N__8736),
            .I(N__8725));
    Odrv4 I__1990 (
            .O(N__8731),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    Odrv4 I__1989 (
            .O(N__8728),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    Odrv4 I__1988 (
            .O(N__8725),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ));
    CascadeMux I__1987 (
            .O(N__8718),
            .I(N__8711));
    InMux I__1986 (
            .O(N__8717),
            .I(N__8705));
    CascadeMux I__1985 (
            .O(N__8716),
            .I(N__8702));
    CascadeMux I__1984 (
            .O(N__8715),
            .I(N__8699));
    CascadeMux I__1983 (
            .O(N__8714),
            .I(N__8695));
    InMux I__1982 (
            .O(N__8711),
            .I(N__8691));
    CascadeMux I__1981 (
            .O(N__8710),
            .I(N__8688));
    CascadeMux I__1980 (
            .O(N__8709),
            .I(N__8685));
    InMux I__1979 (
            .O(N__8708),
            .I(N__8682));
    LocalMux I__1978 (
            .O(N__8705),
            .I(N__8679));
    InMux I__1977 (
            .O(N__8702),
            .I(N__8676));
    InMux I__1976 (
            .O(N__8699),
            .I(N__8673));
    CascadeMux I__1975 (
            .O(N__8698),
            .I(N__8670));
    InMux I__1974 (
            .O(N__8695),
            .I(N__8667));
    InMux I__1973 (
            .O(N__8694),
            .I(N__8663));
    LocalMux I__1972 (
            .O(N__8691),
            .I(N__8660));
    InMux I__1971 (
            .O(N__8688),
            .I(N__8657));
    InMux I__1970 (
            .O(N__8685),
            .I(N__8654));
    LocalMux I__1969 (
            .O(N__8682),
            .I(N__8645));
    Span4Mux_v I__1968 (
            .O(N__8679),
            .I(N__8645));
    LocalMux I__1967 (
            .O(N__8676),
            .I(N__8645));
    LocalMux I__1966 (
            .O(N__8673),
            .I(N__8645));
    InMux I__1965 (
            .O(N__8670),
            .I(N__8642));
    LocalMux I__1964 (
            .O(N__8667),
            .I(N__8637));
    InMux I__1963 (
            .O(N__8666),
            .I(N__8634));
    LocalMux I__1962 (
            .O(N__8663),
            .I(N__8630));
    Span4Mux_v I__1961 (
            .O(N__8660),
            .I(N__8625));
    LocalMux I__1960 (
            .O(N__8657),
            .I(N__8625));
    LocalMux I__1959 (
            .O(N__8654),
            .I(N__8620));
    Span4Mux_h I__1958 (
            .O(N__8645),
            .I(N__8620));
    LocalMux I__1957 (
            .O(N__8642),
            .I(N__8617));
    CascadeMux I__1956 (
            .O(N__8641),
            .I(N__8612));
    InMux I__1955 (
            .O(N__8640),
            .I(N__8609));
    Span4Mux_v I__1954 (
            .O(N__8637),
            .I(N__8604));
    LocalMux I__1953 (
            .O(N__8634),
            .I(N__8604));
    InMux I__1952 (
            .O(N__8633),
            .I(N__8601));
    Span4Mux_h I__1951 (
            .O(N__8630),
            .I(N__8598));
    Span4Mux_h I__1950 (
            .O(N__8625),
            .I(N__8591));
    Span4Mux_h I__1949 (
            .O(N__8620),
            .I(N__8591));
    Span4Mux_h I__1948 (
            .O(N__8617),
            .I(N__8591));
    InMux I__1947 (
            .O(N__8616),
            .I(N__8586));
    InMux I__1946 (
            .O(N__8615),
            .I(N__8586));
    InMux I__1945 (
            .O(N__8612),
            .I(N__8583));
    LocalMux I__1944 (
            .O(N__8609),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1943 (
            .O(N__8604),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1942 (
            .O(N__8601),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1941 (
            .O(N__8598),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1940 (
            .O(N__8591),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1939 (
            .O(N__8586),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1938 (
            .O(N__8583),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__1937 (
            .O(N__8568),
            .I(N__8565));
    LocalMux I__1936 (
            .O(N__8565),
            .I(N__8562));
    Span4Mux_s2_v I__1935 (
            .O(N__8562),
            .I(N__8559));
    Span4Mux_v I__1934 (
            .O(N__8559),
            .I(N__8556));
    Span4Mux_h I__1933 (
            .O(N__8556),
            .I(N__8553));
    Odrv4 I__1932 (
            .O(N__8553),
            .I(CASn_c));
    InMux I__1931 (
            .O(N__8550),
            .I(N__8546));
    InMux I__1930 (
            .O(N__8549),
            .I(N__8543));
    LocalMux I__1929 (
            .O(N__8546),
            .I(N__8538));
    LocalMux I__1928 (
            .O(N__8543),
            .I(N__8538));
    Span12Mux_h I__1927 (
            .O(N__8538),
            .I(N__8532));
    InMux I__1926 (
            .O(N__8537),
            .I(N__8529));
    InMux I__1925 (
            .O(N__8536),
            .I(N__8524));
    InMux I__1924 (
            .O(N__8535),
            .I(N__8524));
    Odrv12 I__1923 (
            .O(N__8532),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1922 (
            .O(N__8529),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__1921 (
            .O(N__8524),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    IoInMux I__1920 (
            .O(N__8517),
            .I(N__8514));
    LocalMux I__1919 (
            .O(N__8514),
            .I(N__8511));
    Span4Mux_s1_v I__1918 (
            .O(N__8511),
            .I(N__8508));
    Span4Mux_v I__1917 (
            .O(N__8508),
            .I(N__8505));
    Span4Mux_v I__1916 (
            .O(N__8505),
            .I(N__8502));
    Odrv4 I__1915 (
            .O(N__8502),
            .I(CRCSn_c));
    InMux I__1914 (
            .O(N__8499),
            .I(N__8496));
    LocalMux I__1913 (
            .O(N__8496),
            .I(N__8493));
    Span12Mux_h I__1912 (
            .O(N__8493),
            .I(N__8490));
    Odrv12 I__1911 (
            .O(N__8490),
            .I(RAS1n_c));
    InMux I__1910 (
            .O(N__8487),
            .I(N__8484));
    LocalMux I__1909 (
            .O(N__8484),
            .I(N__8480));
    InMux I__1908 (
            .O(N__8483),
            .I(N__8477));
    Span4Mux_h I__1907 (
            .O(N__8480),
            .I(N__8472));
    LocalMux I__1906 (
            .O(N__8477),
            .I(N__8472));
    Sp12to4 I__1905 (
            .O(N__8472),
            .I(N__8469));
    Span12Mux_v I__1904 (
            .O(N__8469),
            .I(N__8466));
    Span12Mux_h I__1903 (
            .O(N__8466),
            .I(N__8463));
    Odrv12 I__1902 (
            .O(N__8463),
            .I(DRA_c_6));
    InMux I__1901 (
            .O(N__8460),
            .I(N__8457));
    LocalMux I__1900 (
            .O(N__8457),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__1899 (
            .O(N__8454),
            .I(N__8451));
    LocalMux I__1898 (
            .O(N__8451),
            .I(N__8447));
    InMux I__1897 (
            .O(N__8450),
            .I(N__8444));
    Span4Mux_v I__1896 (
            .O(N__8447),
            .I(N__8441));
    LocalMux I__1895 (
            .O(N__8444),
            .I(N__8438));
    Sp12to4 I__1894 (
            .O(N__8441),
            .I(N__8435));
    Sp12to4 I__1893 (
            .O(N__8438),
            .I(N__8432));
    Span12Mux_h I__1892 (
            .O(N__8435),
            .I(N__8429));
    Span12Mux_v I__1891 (
            .O(N__8432),
            .I(N__8426));
    Span12Mux_v I__1890 (
            .O(N__8429),
            .I(N__8423));
    Span12Mux_h I__1889 (
            .O(N__8426),
            .I(N__8420));
    Odrv12 I__1888 (
            .O(N__8423),
            .I(DRA_c_3));
    Odrv12 I__1887 (
            .O(N__8420),
            .I(DRA_c_3));
    InMux I__1886 (
            .O(N__8415),
            .I(N__8412));
    LocalMux I__1885 (
            .O(N__8412),
            .I(N__8409));
    Span4Mux_h I__1884 (
            .O(N__8409),
            .I(N__8406));
    Odrv4 I__1883 (
            .O(N__8406),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    InMux I__1882 (
            .O(N__8403),
            .I(N__8400));
    LocalMux I__1881 (
            .O(N__8400),
            .I(N__8397));
    Span4Mux_h I__1880 (
            .O(N__8397),
            .I(N__8394));
    Odrv4 I__1879 (
            .O(N__8394),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    CascadeMux I__1878 (
            .O(N__8391),
            .I(N__8387));
    InMux I__1877 (
            .O(N__8390),
            .I(N__8384));
    InMux I__1876 (
            .O(N__8387),
            .I(N__8381));
    LocalMux I__1875 (
            .O(N__8384),
            .I(N__8364));
    LocalMux I__1874 (
            .O(N__8381),
            .I(N__8364));
    InMux I__1873 (
            .O(N__8380),
            .I(N__8361));
    InMux I__1872 (
            .O(N__8379),
            .I(N__8358));
    CascadeMux I__1871 (
            .O(N__8378),
            .I(N__8353));
    InMux I__1870 (
            .O(N__8377),
            .I(N__8350));
    InMux I__1869 (
            .O(N__8376),
            .I(N__8347));
    CascadeMux I__1868 (
            .O(N__8375),
            .I(N__8340));
    InMux I__1867 (
            .O(N__8374),
            .I(N__8335));
    InMux I__1866 (
            .O(N__8373),
            .I(N__8335));
    InMux I__1865 (
            .O(N__8372),
            .I(N__8330));
    InMux I__1864 (
            .O(N__8371),
            .I(N__8330));
    InMux I__1863 (
            .O(N__8370),
            .I(N__8325));
    InMux I__1862 (
            .O(N__8369),
            .I(N__8325));
    Span4Mux_h I__1861 (
            .O(N__8364),
            .I(N__8320));
    LocalMux I__1860 (
            .O(N__8361),
            .I(N__8315));
    LocalMux I__1859 (
            .O(N__8358),
            .I(N__8315));
    InMux I__1858 (
            .O(N__8357),
            .I(N__8311));
    InMux I__1857 (
            .O(N__8356),
            .I(N__8308));
    InMux I__1856 (
            .O(N__8353),
            .I(N__8305));
    LocalMux I__1855 (
            .O(N__8350),
            .I(N__8302));
    LocalMux I__1854 (
            .O(N__8347),
            .I(N__8299));
    InMux I__1853 (
            .O(N__8346),
            .I(N__8295));
    InMux I__1852 (
            .O(N__8345),
            .I(N__8288));
    InMux I__1851 (
            .O(N__8344),
            .I(N__8288));
    InMux I__1850 (
            .O(N__8343),
            .I(N__8288));
    InMux I__1849 (
            .O(N__8340),
            .I(N__8285));
    LocalMux I__1848 (
            .O(N__8335),
            .I(N__8278));
    LocalMux I__1847 (
            .O(N__8330),
            .I(N__8278));
    LocalMux I__1846 (
            .O(N__8325),
            .I(N__8278));
    InMux I__1845 (
            .O(N__8324),
            .I(N__8273));
    InMux I__1844 (
            .O(N__8323),
            .I(N__8273));
    Span4Mux_v I__1843 (
            .O(N__8320),
            .I(N__8267));
    Span4Mux_v I__1842 (
            .O(N__8315),
            .I(N__8267));
    InMux I__1841 (
            .O(N__8314),
            .I(N__8264));
    LocalMux I__1840 (
            .O(N__8311),
            .I(N__8253));
    LocalMux I__1839 (
            .O(N__8308),
            .I(N__8253));
    LocalMux I__1838 (
            .O(N__8305),
            .I(N__8253));
    Span4Mux_v I__1837 (
            .O(N__8302),
            .I(N__8253));
    Span4Mux_h I__1836 (
            .O(N__8299),
            .I(N__8253));
    InMux I__1835 (
            .O(N__8298),
            .I(N__8250));
    LocalMux I__1834 (
            .O(N__8295),
            .I(N__8241));
    LocalMux I__1833 (
            .O(N__8288),
            .I(N__8241));
    LocalMux I__1832 (
            .O(N__8285),
            .I(N__8241));
    Span4Mux_h I__1831 (
            .O(N__8278),
            .I(N__8241));
    LocalMux I__1830 (
            .O(N__8273),
            .I(N__8236));
    InMux I__1829 (
            .O(N__8272),
            .I(N__8233));
    Sp12to4 I__1828 (
            .O(N__8267),
            .I(N__8228));
    LocalMux I__1827 (
            .O(N__8264),
            .I(N__8228));
    Span4Mux_h I__1826 (
            .O(N__8253),
            .I(N__8225));
    LocalMux I__1825 (
            .O(N__8250),
            .I(N__8220));
    Span4Mux_h I__1824 (
            .O(N__8241),
            .I(N__8220));
    InMux I__1823 (
            .O(N__8240),
            .I(N__8215));
    InMux I__1822 (
            .O(N__8239),
            .I(N__8215));
    Odrv4 I__1821 (
            .O(N__8236),
            .I(CPU_CYCLEm));
    LocalMux I__1820 (
            .O(N__8233),
            .I(CPU_CYCLEm));
    Odrv12 I__1819 (
            .O(N__8228),
            .I(CPU_CYCLEm));
    Odrv4 I__1818 (
            .O(N__8225),
            .I(CPU_CYCLEm));
    Odrv4 I__1817 (
            .O(N__8220),
            .I(CPU_CYCLEm));
    LocalMux I__1816 (
            .O(N__8215),
            .I(CPU_CYCLEm));
    InMux I__1815 (
            .O(N__8202),
            .I(N__8199));
    LocalMux I__1814 (
            .O(N__8199),
            .I(N__8196));
    Span12Mux_v I__1813 (
            .O(N__8196),
            .I(N__8193));
    Span12Mux_h I__1812 (
            .O(N__8193),
            .I(N__8190));
    Odrv12 I__1811 (
            .O(N__8190),
            .I(A_c_16));
    CascadeMux I__1810 (
            .O(N__8187),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_7_cascade_ ));
    InMux I__1809 (
            .O(N__8184),
            .I(N__8181));
    LocalMux I__1808 (
            .O(N__8181),
            .I(N__8178));
    Span12Mux_v I__1807 (
            .O(N__8178),
            .I(N__8175));
    Span12Mux_h I__1806 (
            .O(N__8175),
            .I(N__8172));
    Odrv12 I__1805 (
            .O(N__8172),
            .I(A_c_18));
    InMux I__1804 (
            .O(N__8169),
            .I(N__8165));
    InMux I__1803 (
            .O(N__8168),
            .I(N__8162));
    LocalMux I__1802 (
            .O(N__8165),
            .I(N__8159));
    LocalMux I__1801 (
            .O(N__8162),
            .I(N__8156));
    Span4Mux_v I__1800 (
            .O(N__8159),
            .I(N__8153));
    Span12Mux_v I__1799 (
            .O(N__8156),
            .I(N__8148));
    Sp12to4 I__1798 (
            .O(N__8153),
            .I(N__8148));
    Span12Mux_h I__1797 (
            .O(N__8148),
            .I(N__8145));
    Odrv12 I__1796 (
            .O(N__8145),
            .I(DRA_c_8));
    CascadeMux I__1795 (
            .O(N__8142),
            .I(N__8139));
    InMux I__1794 (
            .O(N__8139),
            .I(N__8136));
    LocalMux I__1793 (
            .O(N__8136),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1792 (
            .O(N__8133),
            .I(N__8130));
    LocalMux I__1791 (
            .O(N__8130),
            .I(N__8127));
    Span4Mux_v I__1790 (
            .O(N__8127),
            .I(N__8123));
    InMux I__1789 (
            .O(N__8126),
            .I(N__8120));
    Span4Mux_v I__1788 (
            .O(N__8123),
            .I(N__8117));
    LocalMux I__1787 (
            .O(N__8120),
            .I(N__8114));
    Sp12to4 I__1786 (
            .O(N__8117),
            .I(N__8109));
    Span12Mux_v I__1785 (
            .O(N__8114),
            .I(N__8109));
    Span12Mux_h I__1784 (
            .O(N__8109),
            .I(N__8106));
    Odrv12 I__1783 (
            .O(N__8106),
            .I(DRA_c_7));
    InMux I__1782 (
            .O(N__8103),
            .I(N__8100));
    LocalMux I__1781 (
            .O(N__8100),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__1780 (
            .O(N__8097),
            .I(N__8094));
    LocalMux I__1779 (
            .O(N__8094),
            .I(N__8090));
    InMux I__1778 (
            .O(N__8093),
            .I(N__8087));
    Span4Mux_v I__1777 (
            .O(N__8090),
            .I(N__8082));
    LocalMux I__1776 (
            .O(N__8087),
            .I(N__8082));
    Span4Mux_h I__1775 (
            .O(N__8082),
            .I(N__8079));
    Span4Mux_v I__1774 (
            .O(N__8079),
            .I(N__8076));
    Sp12to4 I__1773 (
            .O(N__8076),
            .I(N__8073));
    Span12Mux_h I__1772 (
            .O(N__8073),
            .I(N__8070));
    Span12Mux_v I__1771 (
            .O(N__8070),
            .I(N__8067));
    Odrv12 I__1770 (
            .O(N__8067),
            .I(DRA_c_0));
    InMux I__1769 (
            .O(N__8064),
            .I(N__8061));
    LocalMux I__1768 (
            .O(N__8061),
            .I(N__8058));
    Odrv4 I__1767 (
            .O(N__8058),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__1766 (
            .O(N__8055),
            .I(N__8052));
    LocalMux I__1765 (
            .O(N__8052),
            .I(N__8049));
    Span4Mux_v I__1764 (
            .O(N__8049),
            .I(N__8045));
    InMux I__1763 (
            .O(N__8048),
            .I(N__8042));
    Sp12to4 I__1762 (
            .O(N__8045),
            .I(N__8039));
    LocalMux I__1761 (
            .O(N__8042),
            .I(N__8036));
    Span12Mux_h I__1760 (
            .O(N__8039),
            .I(N__8033));
    Span12Mux_v I__1759 (
            .O(N__8036),
            .I(N__8030));
    Span12Mux_v I__1758 (
            .O(N__8033),
            .I(N__8027));
    Span12Mux_h I__1757 (
            .O(N__8030),
            .I(N__8024));
    Odrv12 I__1756 (
            .O(N__8027),
            .I(DRA_c_2));
    Odrv12 I__1755 (
            .O(N__8024),
            .I(DRA_c_2));
    InMux I__1754 (
            .O(N__8019),
            .I(N__8016));
    LocalMux I__1753 (
            .O(N__8016),
            .I(N__8013));
    Span4Mux_h I__1752 (
            .O(N__8013),
            .I(N__8010));
    Odrv4 I__1751 (
            .O(N__8010),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    InMux I__1750 (
            .O(N__8007),
            .I(N__8004));
    LocalMux I__1749 (
            .O(N__8004),
            .I(N__7988));
    InMux I__1748 (
            .O(N__8003),
            .I(N__7983));
    InMux I__1747 (
            .O(N__8002),
            .I(N__7983));
    InMux I__1746 (
            .O(N__8001),
            .I(N__7978));
    InMux I__1745 (
            .O(N__8000),
            .I(N__7973));
    InMux I__1744 (
            .O(N__7999),
            .I(N__7973));
    InMux I__1743 (
            .O(N__7998),
            .I(N__7968));
    InMux I__1742 (
            .O(N__7997),
            .I(N__7968));
    InMux I__1741 (
            .O(N__7996),
            .I(N__7959));
    InMux I__1740 (
            .O(N__7995),
            .I(N__7956));
    InMux I__1739 (
            .O(N__7994),
            .I(N__7949));
    InMux I__1738 (
            .O(N__7993),
            .I(N__7949));
    InMux I__1737 (
            .O(N__7992),
            .I(N__7949));
    InMux I__1736 (
            .O(N__7991),
            .I(N__7946));
    Span4Mux_v I__1735 (
            .O(N__7988),
            .I(N__7941));
    LocalMux I__1734 (
            .O(N__7983),
            .I(N__7941));
    InMux I__1733 (
            .O(N__7982),
            .I(N__7938));
    InMux I__1732 (
            .O(N__7981),
            .I(N__7934));
    LocalMux I__1731 (
            .O(N__7978),
            .I(N__7929));
    LocalMux I__1730 (
            .O(N__7973),
            .I(N__7929));
    LocalMux I__1729 (
            .O(N__7968),
            .I(N__7926));
    InMux I__1728 (
            .O(N__7967),
            .I(N__7923));
    InMux I__1727 (
            .O(N__7966),
            .I(N__7912));
    InMux I__1726 (
            .O(N__7965),
            .I(N__7912));
    InMux I__1725 (
            .O(N__7964),
            .I(N__7912));
    InMux I__1724 (
            .O(N__7963),
            .I(N__7912));
    InMux I__1723 (
            .O(N__7962),
            .I(N__7912));
    LocalMux I__1722 (
            .O(N__7959),
            .I(N__7909));
    LocalMux I__1721 (
            .O(N__7956),
            .I(N__7906));
    LocalMux I__1720 (
            .O(N__7949),
            .I(N__7901));
    LocalMux I__1719 (
            .O(N__7946),
            .I(N__7901));
    Span4Mux_v I__1718 (
            .O(N__7941),
            .I(N__7894));
    LocalMux I__1717 (
            .O(N__7938),
            .I(N__7891));
    InMux I__1716 (
            .O(N__7937),
            .I(N__7888));
    LocalMux I__1715 (
            .O(N__7934),
            .I(N__7885));
    Span4Mux_v I__1714 (
            .O(N__7929),
            .I(N__7876));
    Span4Mux_h I__1713 (
            .O(N__7926),
            .I(N__7876));
    LocalMux I__1712 (
            .O(N__7923),
            .I(N__7876));
    LocalMux I__1711 (
            .O(N__7912),
            .I(N__7876));
    Span4Mux_v I__1710 (
            .O(N__7909),
            .I(N__7873));
    Span4Mux_h I__1709 (
            .O(N__7906),
            .I(N__7868));
    Span4Mux_v I__1708 (
            .O(N__7901),
            .I(N__7868));
    InMux I__1707 (
            .O(N__7900),
            .I(N__7861));
    InMux I__1706 (
            .O(N__7899),
            .I(N__7861));
    InMux I__1705 (
            .O(N__7898),
            .I(N__7861));
    InMux I__1704 (
            .O(N__7897),
            .I(N__7858));
    Span4Mux_h I__1703 (
            .O(N__7894),
            .I(N__7851));
    Span4Mux_v I__1702 (
            .O(N__7891),
            .I(N__7851));
    LocalMux I__1701 (
            .O(N__7888),
            .I(N__7851));
    Span4Mux_v I__1700 (
            .O(N__7885),
            .I(N__7846));
    Span4Mux_v I__1699 (
            .O(N__7876),
            .I(N__7846));
    Span4Mux_h I__1698 (
            .O(N__7873),
            .I(N__7841));
    Span4Mux_v I__1697 (
            .O(N__7868),
            .I(N__7841));
    LocalMux I__1696 (
            .O(N__7861),
            .I(N__7838));
    LocalMux I__1695 (
            .O(N__7858),
            .I(N__7833));
    Sp12to4 I__1694 (
            .O(N__7851),
            .I(N__7833));
    Sp12to4 I__1693 (
            .O(N__7846),
            .I(N__7830));
    Sp12to4 I__1692 (
            .O(N__7841),
            .I(N__7823));
    Span12Mux_h I__1691 (
            .O(N__7838),
            .I(N__7823));
    Span12Mux_v I__1690 (
            .O(N__7833),
            .I(N__7823));
    Span12Mux_h I__1689 (
            .O(N__7830),
            .I(N__7820));
    Span12Mux_h I__1688 (
            .O(N__7823),
            .I(N__7817));
    Odrv12 I__1687 (
            .O(N__7820),
            .I(RESETn_c));
    Odrv12 I__1686 (
            .O(N__7817),
            .I(RESETn_c));
    IoInMux I__1685 (
            .O(N__7812),
            .I(N__7809));
    LocalMux I__1684 (
            .O(N__7809),
            .I(N__7806));
    Odrv12 I__1683 (
            .O(N__7806),
            .I(RESETn_c_i));
    IoInMux I__1682 (
            .O(N__7803),
            .I(N__7800));
    LocalMux I__1681 (
            .O(N__7800),
            .I(N__7797));
    Span4Mux_s2_v I__1680 (
            .O(N__7797),
            .I(N__7794));
    Span4Mux_v I__1679 (
            .O(N__7794),
            .I(N__7791));
    Span4Mux_h I__1678 (
            .O(N__7791),
            .I(N__7788));
    Odrv4 I__1677 (
            .O(N__7788),
            .I(CMA_c_0));
    InMux I__1676 (
            .O(N__7785),
            .I(N__7782));
    LocalMux I__1675 (
            .O(N__7782),
            .I(\U712_CHIP_RAM.N_36 ));
    IoInMux I__1674 (
            .O(N__7779),
            .I(N__7776));
    LocalMux I__1673 (
            .O(N__7776),
            .I(N__7773));
    IoSpan4Mux I__1672 (
            .O(N__7773),
            .I(N__7770));
    IoSpan4Mux I__1671 (
            .O(N__7770),
            .I(N__7767));
    Span4Mux_s3_h I__1670 (
            .O(N__7767),
            .I(N__7764));
    Span4Mux_h I__1669 (
            .O(N__7764),
            .I(N__7761));
    Span4Mux_h I__1668 (
            .O(N__7761),
            .I(N__7758));
    Odrv4 I__1667 (
            .O(N__7758),
            .I(CMA_c_5));
    InMux I__1666 (
            .O(N__7755),
            .I(N__7752));
    LocalMux I__1665 (
            .O(N__7752),
            .I(N__7749));
    Odrv4 I__1664 (
            .O(N__7749),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1663 (
            .O(N__7746),
            .I(N__7743));
    LocalMux I__1662 (
            .O(N__7743),
            .I(N__7740));
    Span4Mux_v I__1661 (
            .O(N__7740),
            .I(N__7737));
    Span4Mux_v I__1660 (
            .O(N__7737),
            .I(N__7734));
    Sp12to4 I__1659 (
            .O(N__7734),
            .I(N__7731));
    Span12Mux_h I__1658 (
            .O(N__7731),
            .I(N__7728));
    Odrv12 I__1657 (
            .O(N__7728),
            .I(A_c_9));
    CascadeMux I__1656 (
            .O(N__7725),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_ ));
    InMux I__1655 (
            .O(N__7722),
            .I(N__7719));
    LocalMux I__1654 (
            .O(N__7719),
            .I(N__7716));
    Span4Mux_v I__1653 (
            .O(N__7716),
            .I(N__7713));
    Span4Mux_v I__1652 (
            .O(N__7713),
            .I(N__7710));
    Sp12to4 I__1651 (
            .O(N__7710),
            .I(N__7707));
    Span12Mux_h I__1650 (
            .O(N__7707),
            .I(N__7704));
    Span12Mux_v I__1649 (
            .O(N__7704),
            .I(N__7701));
    Odrv12 I__1648 (
            .O(N__7701),
            .I(A_c_2));
    InMux I__1647 (
            .O(N__7698),
            .I(N__7695));
    LocalMux I__1646 (
            .O(N__7695),
            .I(\U712_CHIP_RAM.N_31 ));
    InMux I__1645 (
            .O(N__7692),
            .I(N__7689));
    LocalMux I__1644 (
            .O(N__7689),
            .I(N__7686));
    Span4Mux_v I__1643 (
            .O(N__7686),
            .I(N__7683));
    Span4Mux_v I__1642 (
            .O(N__7683),
            .I(N__7680));
    Sp12to4 I__1641 (
            .O(N__7680),
            .I(N__7677));
    Span12Mux_h I__1640 (
            .O(N__7677),
            .I(N__7674));
    Odrv12 I__1639 (
            .O(N__7674),
            .I(A_c_17));
    IoInMux I__1638 (
            .O(N__7671),
            .I(N__7668));
    LocalMux I__1637 (
            .O(N__7668),
            .I(N__7665));
    IoSpan4Mux I__1636 (
            .O(N__7665),
            .I(N__7662));
    Span4Mux_s1_h I__1635 (
            .O(N__7662),
            .I(N__7659));
    Sp12to4 I__1634 (
            .O(N__7659),
            .I(N__7656));
    Span12Mux_h I__1633 (
            .O(N__7656),
            .I(N__7653));
    Odrv12 I__1632 (
            .O(N__7653),
            .I(CMA_c_8));
    IoInMux I__1631 (
            .O(N__7650),
            .I(N__7647));
    LocalMux I__1630 (
            .O(N__7647),
            .I(N__7644));
    Span12Mux_s3_h I__1629 (
            .O(N__7644),
            .I(N__7641));
    Span12Mux_h I__1628 (
            .O(N__7641),
            .I(N__7638));
    Odrv12 I__1627 (
            .O(N__7638),
            .I(CMA_c_6));
    InMux I__1626 (
            .O(N__7635),
            .I(N__7631));
    InMux I__1625 (
            .O(N__7634),
            .I(N__7628));
    LocalMux I__1624 (
            .O(N__7631),
            .I(N__7625));
    LocalMux I__1623 (
            .O(N__7628),
            .I(N__7622));
    Span4Mux_h I__1622 (
            .O(N__7625),
            .I(N__7619));
    Odrv12 I__1621 (
            .O(N__7622),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    Odrv4 I__1620 (
            .O(N__7619),
            .I(\U712_CHIP_RAM.CMA_5_0_8 ));
    CascadeMux I__1619 (
            .O(N__7614),
            .I(N__7611));
    InMux I__1618 (
            .O(N__7611),
            .I(N__7608));
    LocalMux I__1617 (
            .O(N__7608),
            .I(N__7605));
    Span4Mux_v I__1616 (
            .O(N__7605),
            .I(N__7602));
    Span4Mux_v I__1615 (
            .O(N__7602),
            .I(N__7599));
    Sp12to4 I__1614 (
            .O(N__7599),
            .I(N__7596));
    Span12Mux_h I__1613 (
            .O(N__7596),
            .I(N__7593));
    Odrv12 I__1612 (
            .O(N__7593),
            .I(A_c_19));
    IoInMux I__1611 (
            .O(N__7590),
            .I(N__7587));
    LocalMux I__1610 (
            .O(N__7587),
            .I(N__7584));
    Span12Mux_s3_h I__1609 (
            .O(N__7584),
            .I(N__7581));
    Span12Mux_h I__1608 (
            .O(N__7581),
            .I(N__7578));
    Odrv12 I__1607 (
            .O(N__7578),
            .I(CMA_c_9));
    InMux I__1606 (
            .O(N__7575),
            .I(N__7572));
    LocalMux I__1605 (
            .O(N__7572),
            .I(N__7569));
    Span4Mux_v I__1604 (
            .O(N__7569),
            .I(N__7566));
    Span4Mux_v I__1603 (
            .O(N__7566),
            .I(N__7563));
    Sp12to4 I__1602 (
            .O(N__7563),
            .I(N__7560));
    Span12Mux_h I__1601 (
            .O(N__7560),
            .I(N__7557));
    Odrv12 I__1600 (
            .O(N__7557),
            .I(A_c_15));
    InMux I__1599 (
            .O(N__7554),
            .I(N__7551));
    LocalMux I__1598 (
            .O(N__7551),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_6 ));
    CascadeMux I__1597 (
            .O(N__7548),
            .I(N__7545));
    InMux I__1596 (
            .O(N__7545),
            .I(N__7542));
    LocalMux I__1595 (
            .O(N__7542),
            .I(N__7539));
    Span4Mux_h I__1594 (
            .O(N__7539),
            .I(N__7536));
    Span4Mux_v I__1593 (
            .O(N__7536),
            .I(N__7533));
    Sp12to4 I__1592 (
            .O(N__7533),
            .I(N__7530));
    Span12Mux_h I__1591 (
            .O(N__7530),
            .I(N__7527));
    Odrv12 I__1590 (
            .O(N__7527),
            .I(A_c_8));
    InMux I__1589 (
            .O(N__7524),
            .I(N__7521));
    LocalMux I__1588 (
            .O(N__7521),
            .I(\U712_CHIP_RAM.N_37 ));
    InMux I__1587 (
            .O(N__7518),
            .I(N__7514));
    InMux I__1586 (
            .O(N__7517),
            .I(N__7511));
    LocalMux I__1585 (
            .O(N__7514),
            .I(N__7506));
    LocalMux I__1584 (
            .O(N__7511),
            .I(N__7506));
    Sp12to4 I__1583 (
            .O(N__7506),
            .I(N__7503));
    Span12Mux_v I__1582 (
            .O(N__7503),
            .I(N__7500));
    Span12Mux_h I__1581 (
            .O(N__7500),
            .I(N__7497));
    Odrv12 I__1580 (
            .O(N__7497),
            .I(DRA_c_4));
    InMux I__1579 (
            .O(N__7494),
            .I(N__7491));
    LocalMux I__1578 (
            .O(N__7491),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__1577 (
            .O(N__7488),
            .I(N__7484));
    InMux I__1576 (
            .O(N__7487),
            .I(N__7481));
    LocalMux I__1575 (
            .O(N__7484),
            .I(N__7478));
    LocalMux I__1574 (
            .O(N__7481),
            .I(N__7475));
    Span4Mux_v I__1573 (
            .O(N__7478),
            .I(N__7472));
    Span4Mux_h I__1572 (
            .O(N__7475),
            .I(N__7469));
    Sp12to4 I__1571 (
            .O(N__7472),
            .I(N__7466));
    Sp12to4 I__1570 (
            .O(N__7469),
            .I(N__7463));
    Span12Mux_h I__1569 (
            .O(N__7466),
            .I(N__7460));
    Span12Mux_v I__1568 (
            .O(N__7463),
            .I(N__7457));
    Span12Mux_v I__1567 (
            .O(N__7460),
            .I(N__7452));
    Span12Mux_h I__1566 (
            .O(N__7457),
            .I(N__7452));
    Odrv12 I__1565 (
            .O(N__7452),
            .I(DRA_c_5));
    InMux I__1564 (
            .O(N__7449),
            .I(N__7446));
    LocalMux I__1563 (
            .O(N__7446),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1562 (
            .O(N__7443),
            .I(N__7440));
    LocalMux I__1561 (
            .O(N__7440),
            .I(\U712_CHIP_RAM.N_32 ));
    IoInMux I__1560 (
            .O(N__7437),
            .I(N__7434));
    LocalMux I__1559 (
            .O(N__7434),
            .I(N__7431));
    Span12Mux_s8_v I__1558 (
            .O(N__7431),
            .I(N__7428));
    Odrv12 I__1557 (
            .O(N__7428),
            .I(CMA_c_1));
    InMux I__1556 (
            .O(N__7425),
            .I(N__7422));
    LocalMux I__1555 (
            .O(N__7422),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1554 (
            .O(N__7419),
            .I(N__7416));
    LocalMux I__1553 (
            .O(N__7416),
            .I(N__7413));
    Odrv12 I__1552 (
            .O(N__7413),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    CEMux I__1551 (
            .O(N__7410),
            .I(N__7406));
    CEMux I__1550 (
            .O(N__7409),
            .I(N__7403));
    LocalMux I__1549 (
            .O(N__7406),
            .I(N__7400));
    LocalMux I__1548 (
            .O(N__7403),
            .I(N__7397));
    Odrv12 I__1547 (
            .O(N__7400),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    Odrv12 I__1546 (
            .O(N__7397),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ));
    InMux I__1545 (
            .O(N__7392),
            .I(N__7389));
    LocalMux I__1544 (
            .O(N__7389),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__1543 (
            .O(N__7386),
            .I(N__7382));
    InMux I__1542 (
            .O(N__7385),
            .I(N__7379));
    LocalMux I__1541 (
            .O(N__7382),
            .I(N__7373));
    LocalMux I__1540 (
            .O(N__7379),
            .I(N__7373));
    InMux I__1539 (
            .O(N__7378),
            .I(N__7370));
    Span4Mux_v I__1538 (
            .O(N__7373),
            .I(N__7367));
    LocalMux I__1537 (
            .O(N__7370),
            .I(N__7364));
    Sp12to4 I__1536 (
            .O(N__7367),
            .I(N__7361));
    Span12Mux_h I__1535 (
            .O(N__7364),
            .I(N__7358));
    Span12Mux_h I__1534 (
            .O(N__7361),
            .I(N__7355));
    Span12Mux_v I__1533 (
            .O(N__7358),
            .I(N__7352));
    Span12Mux_v I__1532 (
            .O(N__7355),
            .I(N__7349));
    Odrv12 I__1531 (
            .O(N__7352),
            .I(CASLn_c));
    Odrv12 I__1530 (
            .O(N__7349),
            .I(CASLn_c));
    InMux I__1529 (
            .O(N__7344),
            .I(N__7341));
    LocalMux I__1528 (
            .O(N__7341),
            .I(N__7338));
    Span4Mux_v I__1527 (
            .O(N__7338),
            .I(N__7333));
    InMux I__1526 (
            .O(N__7337),
            .I(N__7330));
    InMux I__1525 (
            .O(N__7336),
            .I(N__7327));
    Sp12to4 I__1524 (
            .O(N__7333),
            .I(N__7320));
    LocalMux I__1523 (
            .O(N__7330),
            .I(N__7320));
    LocalMux I__1522 (
            .O(N__7327),
            .I(N__7320));
    Span12Mux_h I__1521 (
            .O(N__7320),
            .I(N__7317));
    Span12Mux_v I__1520 (
            .O(N__7317),
            .I(N__7314));
    Odrv12 I__1519 (
            .O(N__7314),
            .I(CASUn_c));
    InMux I__1518 (
            .O(N__7311),
            .I(N__7307));
    InMux I__1517 (
            .O(N__7310),
            .I(N__7304));
    LocalMux I__1516 (
            .O(N__7307),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    LocalMux I__1515 (
            .O(N__7304),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__1514 (
            .O(N__7299),
            .I(N__7296));
    LocalMux I__1513 (
            .O(N__7296),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    InMux I__1512 (
            .O(N__7293),
            .I(N__7290));
    LocalMux I__1511 (
            .O(N__7290),
            .I(N__7286));
    InMux I__1510 (
            .O(N__7289),
            .I(N__7283));
    Odrv4 I__1509 (
            .O(N__7286),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    LocalMux I__1508 (
            .O(N__7283),
            .I(\U712_REG_SM.UDS_OUTZ0 ));
    InMux I__1507 (
            .O(N__7278),
            .I(N__7274));
    InMux I__1506 (
            .O(N__7277),
            .I(N__7271));
    LocalMux I__1505 (
            .O(N__7274),
            .I(N__7266));
    LocalMux I__1504 (
            .O(N__7271),
            .I(N__7266));
    Span4Mux_v I__1503 (
            .O(N__7266),
            .I(N__7262));
    InMux I__1502 (
            .O(N__7265),
            .I(N__7259));
    Odrv4 I__1501 (
            .O(N__7262),
            .I(\U712_REG_SM.DS_ENZ0 ));
    LocalMux I__1500 (
            .O(N__7259),
            .I(\U712_REG_SM.DS_ENZ0 ));
    IoInMux I__1499 (
            .O(N__7254),
            .I(N__7251));
    LocalMux I__1498 (
            .O(N__7251),
            .I(N__7248));
    Span12Mux_s4_v I__1497 (
            .O(N__7248),
            .I(N__7245));
    Span12Mux_h I__1496 (
            .O(N__7245),
            .I(N__7242));
    Odrv12 I__1495 (
            .O(N__7242),
            .I(U712_REG_SM_un1_UDSn_i));
    InMux I__1494 (
            .O(N__7239),
            .I(N__7235));
    CascadeMux I__1493 (
            .O(N__7238),
            .I(N__7230));
    LocalMux I__1492 (
            .O(N__7235),
            .I(N__7226));
    InMux I__1491 (
            .O(N__7234),
            .I(N__7218));
    InMux I__1490 (
            .O(N__7233),
            .I(N__7218));
    InMux I__1489 (
            .O(N__7230),
            .I(N__7218));
    InMux I__1488 (
            .O(N__7229),
            .I(N__7215));
    Span4Mux_v I__1487 (
            .O(N__7226),
            .I(N__7211));
    InMux I__1486 (
            .O(N__7225),
            .I(N__7208));
    LocalMux I__1485 (
            .O(N__7218),
            .I(N__7205));
    LocalMux I__1484 (
            .O(N__7215),
            .I(N__7202));
    InMux I__1483 (
            .O(N__7214),
            .I(N__7199));
    Span4Mux_v I__1482 (
            .O(N__7211),
            .I(N__7194));
    LocalMux I__1481 (
            .O(N__7208),
            .I(N__7194));
    Odrv12 I__1480 (
            .O(N__7205),
            .I(DMA_CYCLEm));
    Odrv4 I__1479 (
            .O(N__7202),
            .I(DMA_CYCLEm));
    LocalMux I__1478 (
            .O(N__7199),
            .I(DMA_CYCLEm));
    Odrv4 I__1477 (
            .O(N__7194),
            .I(DMA_CYCLEm));
    InMux I__1476 (
            .O(N__7185),
            .I(N__7181));
    InMux I__1475 (
            .O(N__7184),
            .I(N__7178));
    LocalMux I__1474 (
            .O(N__7181),
            .I(N__7175));
    LocalMux I__1473 (
            .O(N__7178),
            .I(N__7172));
    Span4Mux_v I__1472 (
            .O(N__7175),
            .I(N__7167));
    Span4Mux_v I__1471 (
            .O(N__7172),
            .I(N__7164));
    InMux I__1470 (
            .O(N__7171),
            .I(N__7161));
    InMux I__1469 (
            .O(N__7170),
            .I(N__7158));
    Odrv4 I__1468 (
            .O(N__7167),
            .I(REG_CYCLEm));
    Odrv4 I__1467 (
            .O(N__7164),
            .I(REG_CYCLEm));
    LocalMux I__1466 (
            .O(N__7161),
            .I(REG_CYCLEm));
    LocalMux I__1465 (
            .O(N__7158),
            .I(REG_CYCLEm));
    IoInMux I__1464 (
            .O(N__7149),
            .I(N__7146));
    LocalMux I__1463 (
            .O(N__7146),
            .I(N__7143));
    Span4Mux_s3_v I__1462 (
            .O(N__7143),
            .I(N__7140));
    Span4Mux_h I__1461 (
            .O(N__7140),
            .I(N__7137));
    Sp12to4 I__1460 (
            .O(N__7137),
            .I(N__7134));
    Span12Mux_v I__1459 (
            .O(N__7134),
            .I(N__7131));
    Span12Mux_h I__1458 (
            .O(N__7131),
            .I(N__7128));
    Odrv12 I__1457 (
            .O(N__7128),
            .I(DRDENn_c));
    IoInMux I__1456 (
            .O(N__7125),
            .I(N__7122));
    LocalMux I__1455 (
            .O(N__7122),
            .I(N__7119));
    Span4Mux_s2_v I__1454 (
            .O(N__7119),
            .I(N__7116));
    Span4Mux_v I__1453 (
            .O(N__7116),
            .I(N__7113));
    Odrv4 I__1452 (
            .O(N__7113),
            .I(CONSTANT_ONE_NET));
    InMux I__1451 (
            .O(N__7110),
            .I(N__7107));
    LocalMux I__1450 (
            .O(N__7107),
            .I(N__7104));
    Span4Mux_v I__1449 (
            .O(N__7104),
            .I(N__7101));
    Sp12to4 I__1448 (
            .O(N__7101),
            .I(N__7098));
    Span12Mux_h I__1447 (
            .O(N__7098),
            .I(N__7095));
    Odrv12 I__1446 (
            .O(N__7095),
            .I(A_c_14));
    CascadeMux I__1445 (
            .O(N__7092),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_5_cascade_ ));
    InMux I__1444 (
            .O(N__7089),
            .I(N__7086));
    LocalMux I__1443 (
            .O(N__7086),
            .I(N__7083));
    Span12Mux_v I__1442 (
            .O(N__7083),
            .I(N__7080));
    Span12Mux_h I__1441 (
            .O(N__7080),
            .I(N__7077));
    Odrv12 I__1440 (
            .O(N__7077),
            .I(A_c_7));
    InMux I__1439 (
            .O(N__7074),
            .I(N__7071));
    LocalMux I__1438 (
            .O(N__7071),
            .I(N__7068));
    Odrv4 I__1437 (
            .O(N__7068),
            .I(\U712_CHIP_RAM.un1_CMA31_0_i ));
    InMux I__1436 (
            .O(N__7065),
            .I(N__7062));
    LocalMux I__1435 (
            .O(N__7062),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__1434 (
            .O(N__7059),
            .I(N__7056));
    LocalMux I__1433 (
            .O(N__7056),
            .I(N__7053));
    Span4Mux_v I__1432 (
            .O(N__7053),
            .I(N__7050));
    Sp12to4 I__1431 (
            .O(N__7050),
            .I(N__7047));
    Span12Mux_h I__1430 (
            .O(N__7047),
            .I(N__7044));
    Odrv12 I__1429 (
            .O(N__7044),
            .I(A_c_10));
    CascadeMux I__1428 (
            .O(N__7041),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_ ));
    InMux I__1427 (
            .O(N__7038),
            .I(N__7035));
    LocalMux I__1426 (
            .O(N__7035),
            .I(N__7032));
    Span12Mux_h I__1425 (
            .O(N__7032),
            .I(N__7029));
    Span12Mux_v I__1424 (
            .O(N__7029),
            .I(N__7026));
    Odrv12 I__1423 (
            .O(N__7026),
            .I(A_c_3));
    InMux I__1422 (
            .O(N__7023),
            .I(N__7020));
    LocalMux I__1421 (
            .O(N__7020),
            .I(N__7017));
    Odrv12 I__1420 (
            .O(N__7017),
            .I(\U712_CHIP_RAM.DBENn_7_0_a2_0 ));
    InMux I__1419 (
            .O(N__7014),
            .I(N__7011));
    LocalMux I__1418 (
            .O(N__7011),
            .I(N__7007));
    InMux I__1417 (
            .O(N__7010),
            .I(N__7004));
    Span4Mux_v I__1416 (
            .O(N__7007),
            .I(N__7001));
    LocalMux I__1415 (
            .O(N__7004),
            .I(N__6998));
    Span4Mux_h I__1414 (
            .O(N__7001),
            .I(N__6993));
    Span4Mux_v I__1413 (
            .O(N__6998),
            .I(N__6993));
    Span4Mux_h I__1412 (
            .O(N__6993),
            .I(N__6990));
    Sp12to4 I__1411 (
            .O(N__6990),
            .I(N__6986));
    IoInMux I__1410 (
            .O(N__6989),
            .I(N__6983));
    Span12Mux_v I__1409 (
            .O(N__6986),
            .I(N__6980));
    LocalMux I__1408 (
            .O(N__6983),
            .I(N__6977));
    Odrv12 I__1407 (
            .O(N__6980),
            .I(AWEn_c));
    Odrv4 I__1406 (
            .O(N__6977),
            .I(AWEn_c));
    InMux I__1405 (
            .O(N__6972),
            .I(N__6968));
    InMux I__1404 (
            .O(N__6971),
            .I(N__6965));
    LocalMux I__1403 (
            .O(N__6968),
            .I(N__6959));
    LocalMux I__1402 (
            .O(N__6965),
            .I(N__6956));
    CascadeMux I__1401 (
            .O(N__6964),
            .I(N__6953));
    CascadeMux I__1400 (
            .O(N__6963),
            .I(N__6950));
    InMux I__1399 (
            .O(N__6962),
            .I(N__6947));
    Span4Mux_v I__1398 (
            .O(N__6959),
            .I(N__6944));
    Span4Mux_v I__1397 (
            .O(N__6956),
            .I(N__6941));
    InMux I__1396 (
            .O(N__6953),
            .I(N__6938));
    InMux I__1395 (
            .O(N__6950),
            .I(N__6935));
    LocalMux I__1394 (
            .O(N__6947),
            .I(N__6932));
    Sp12to4 I__1393 (
            .O(N__6944),
            .I(N__6923));
    Sp12to4 I__1392 (
            .O(N__6941),
            .I(N__6923));
    LocalMux I__1391 (
            .O(N__6938),
            .I(N__6923));
    LocalMux I__1390 (
            .O(N__6935),
            .I(N__6923));
    Span12Mux_v I__1389 (
            .O(N__6932),
            .I(N__6920));
    Span12Mux_h I__1388 (
            .O(N__6923),
            .I(N__6917));
    Span12Mux_h I__1387 (
            .O(N__6920),
            .I(N__6914));
    Span12Mux_v I__1386 (
            .O(N__6917),
            .I(N__6911));
    Odrv12 I__1385 (
            .O(N__6914),
            .I(RnW_c));
    Odrv12 I__1384 (
            .O(N__6911),
            .I(RnW_c));
    InMux I__1383 (
            .O(N__6906),
            .I(N__6900));
    InMux I__1382 (
            .O(N__6905),
            .I(N__6897));
    InMux I__1381 (
            .O(N__6904),
            .I(N__6891));
    InMux I__1380 (
            .O(N__6903),
            .I(N__6888));
    LocalMux I__1379 (
            .O(N__6900),
            .I(N__6883));
    LocalMux I__1378 (
            .O(N__6897),
            .I(N__6883));
    InMux I__1377 (
            .O(N__6896),
            .I(N__6878));
    InMux I__1376 (
            .O(N__6895),
            .I(N__6878));
    InMux I__1375 (
            .O(N__6894),
            .I(N__6875));
    LocalMux I__1374 (
            .O(N__6891),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1373 (
            .O(N__6888),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1372 (
            .O(N__6883),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1371 (
            .O(N__6878),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1370 (
            .O(N__6875),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    InMux I__1369 (
            .O(N__6864),
            .I(N__6861));
    LocalMux I__1368 (
            .O(N__6861),
            .I(N__6857));
    InMux I__1367 (
            .O(N__6860),
            .I(N__6854));
    Span4Mux_h I__1366 (
            .O(N__6857),
            .I(N__6851));
    LocalMux I__1365 (
            .O(N__6854),
            .I(N__6848));
    Odrv4 I__1364 (
            .O(N__6851),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__1363 (
            .O(N__6848),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    CEMux I__1362 (
            .O(N__6843),
            .I(N__6840));
    LocalMux I__1361 (
            .O(N__6840),
            .I(N__6837));
    Odrv4 I__1360 (
            .O(N__6837),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0 ));
    InMux I__1359 (
            .O(N__6834),
            .I(N__6831));
    LocalMux I__1358 (
            .O(N__6831),
            .I(N__6827));
    InMux I__1357 (
            .O(N__6830),
            .I(N__6824));
    Odrv4 I__1356 (
            .O(N__6827),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    LocalMux I__1355 (
            .O(N__6824),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    InMux I__1354 (
            .O(N__6819),
            .I(N__6813));
    InMux I__1353 (
            .O(N__6818),
            .I(N__6806));
    InMux I__1352 (
            .O(N__6817),
            .I(N__6806));
    InMux I__1351 (
            .O(N__6816),
            .I(N__6806));
    LocalMux I__1350 (
            .O(N__6813),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    LocalMux I__1349 (
            .O(N__6806),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    InMux I__1348 (
            .O(N__6801),
            .I(N__6798));
    LocalMux I__1347 (
            .O(N__6798),
            .I(N__6795));
    Span12Mux_v I__1346 (
            .O(N__6795),
            .I(N__6792));
    Odrv12 I__1345 (
            .O(N__6792),
            .I(TACK_EN_i_ess));
    CEMux I__1344 (
            .O(N__6789),
            .I(N__6786));
    LocalMux I__1343 (
            .O(N__6786),
            .I(\U712_CYCLE_TERM.N_45_0_0_en_0 ));
    CascadeMux I__1342 (
            .O(N__6783),
            .I(N__6780));
    InMux I__1341 (
            .O(N__6780),
            .I(N__6776));
    InMux I__1340 (
            .O(N__6779),
            .I(N__6773));
    LocalMux I__1339 (
            .O(N__6776),
            .I(N__6768));
    LocalMux I__1338 (
            .O(N__6773),
            .I(N__6768));
    Odrv12 I__1337 (
            .O(N__6768),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESS4 ));
    InMux I__1336 (
            .O(N__6765),
            .I(N__6762));
    LocalMux I__1335 (
            .O(N__6762),
            .I(\U712_CHIP_RAM.N_33 ));
    IoInMux I__1334 (
            .O(N__6759),
            .I(N__6756));
    LocalMux I__1333 (
            .O(N__6756),
            .I(N__6753));
    Span12Mux_s2_v I__1332 (
            .O(N__6753),
            .I(N__6750));
    Odrv12 I__1331 (
            .O(N__6750),
            .I(CMA_c_2));
    InMux I__1330 (
            .O(N__6747),
            .I(N__6744));
    LocalMux I__1329 (
            .O(N__6744),
            .I(N__6741));
    Span4Mux_v I__1328 (
            .O(N__6741),
            .I(N__6738));
    Sp12to4 I__1327 (
            .O(N__6738),
            .I(N__6735));
    Span12Mux_h I__1326 (
            .O(N__6735),
            .I(N__6732));
    Odrv12 I__1325 (
            .O(N__6732),
            .I(A_c_13));
    CascadeMux I__1324 (
            .O(N__6729),
            .I(N__6726));
    InMux I__1323 (
            .O(N__6726),
            .I(N__6723));
    LocalMux I__1322 (
            .O(N__6723),
            .I(N__6720));
    Span4Mux_v I__1321 (
            .O(N__6720),
            .I(N__6717));
    Sp12to4 I__1320 (
            .O(N__6717),
            .I(N__6714));
    Span12Mux_h I__1319 (
            .O(N__6714),
            .I(N__6711));
    Span12Mux_v I__1318 (
            .O(N__6711),
            .I(N__6708));
    Odrv12 I__1317 (
            .O(N__6708),
            .I(A_c_6));
    CascadeMux I__1316 (
            .O(N__6705),
            .I(\U712_CHIP_RAM.N_35_cascade_ ));
    IoInMux I__1315 (
            .O(N__6702),
            .I(N__6699));
    LocalMux I__1314 (
            .O(N__6699),
            .I(N__6696));
    IoSpan4Mux I__1313 (
            .O(N__6696),
            .I(N__6693));
    IoSpan4Mux I__1312 (
            .O(N__6693),
            .I(N__6690));
    Span4Mux_s2_h I__1311 (
            .O(N__6690),
            .I(N__6687));
    Span4Mux_h I__1310 (
            .O(N__6687),
            .I(N__6684));
    Sp12to4 I__1309 (
            .O(N__6684),
            .I(N__6681));
    Odrv12 I__1308 (
            .O(N__6681),
            .I(CMA_c_4));
    InMux I__1307 (
            .O(N__6678),
            .I(N__6675));
    LocalMux I__1306 (
            .O(N__6675),
            .I(N__6672));
    Span4Mux_v I__1305 (
            .O(N__6672),
            .I(N__6669));
    Sp12to4 I__1304 (
            .O(N__6669),
            .I(N__6666));
    Span12Mux_h I__1303 (
            .O(N__6666),
            .I(N__6663));
    Odrv12 I__1302 (
            .O(N__6663),
            .I(A_c_12));
    CascadeMux I__1301 (
            .O(N__6660),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_ ));
    InMux I__1300 (
            .O(N__6657),
            .I(N__6654));
    LocalMux I__1299 (
            .O(N__6654),
            .I(N__6651));
    Sp12to4 I__1298 (
            .O(N__6651),
            .I(N__6648));
    Span12Mux_v I__1297 (
            .O(N__6648),
            .I(N__6645));
    Span12Mux_h I__1296 (
            .O(N__6645),
            .I(N__6642));
    Odrv12 I__1295 (
            .O(N__6642),
            .I(A_c_5));
    InMux I__1294 (
            .O(N__6639),
            .I(N__6636));
    LocalMux I__1293 (
            .O(N__6636),
            .I(\U712_CHIP_RAM.N_34 ));
    InMux I__1292 (
            .O(N__6633),
            .I(N__6630));
    LocalMux I__1291 (
            .O(N__6630),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_4 ));
    CascadeMux I__1290 (
            .O(N__6627),
            .I(N__6624));
    InMux I__1289 (
            .O(N__6624),
            .I(N__6621));
    LocalMux I__1288 (
            .O(N__6621),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__1287 (
            .O(N__6618),
            .I(N__6615));
    LocalMux I__1286 (
            .O(N__6615),
            .I(N__6612));
    Odrv4 I__1285 (
            .O(N__6612),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__1284 (
            .O(N__6609),
            .I(N__6606));
    LocalMux I__1283 (
            .O(N__6606),
            .I(N__6603));
    Odrv4 I__1282 (
            .O(N__6603),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1281 (
            .O(N__6600),
            .I(N__6597));
    LocalMux I__1280 (
            .O(N__6597),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ));
    InMux I__1279 (
            .O(N__6594),
            .I(N__6590));
    InMux I__1278 (
            .O(N__6593),
            .I(N__6587));
    LocalMux I__1277 (
            .O(N__6590),
            .I(N__6583));
    LocalMux I__1276 (
            .O(N__6587),
            .I(N__6580));
    InMux I__1275 (
            .O(N__6586),
            .I(N__6577));
    Span4Mux_v I__1274 (
            .O(N__6583),
            .I(N__6574));
    Span4Mux_h I__1273 (
            .O(N__6580),
            .I(N__6569));
    LocalMux I__1272 (
            .O(N__6577),
            .I(N__6569));
    Odrv4 I__1271 (
            .O(N__6574),
            .I(U712_REG_SM_DBR_SYNC_1));
    Odrv4 I__1270 (
            .O(N__6569),
            .I(U712_REG_SM_DBR_SYNC_1));
    InMux I__1269 (
            .O(N__6564),
            .I(N__6558));
    InMux I__1268 (
            .O(N__6563),
            .I(N__6555));
    InMux I__1267 (
            .O(N__6562),
            .I(N__6550));
    InMux I__1266 (
            .O(N__6561),
            .I(N__6550));
    LocalMux I__1265 (
            .O(N__6558),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1264 (
            .O(N__6555),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__1263 (
            .O(N__6550),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    CascadeMux I__1262 (
            .O(N__6543),
            .I(N__6540));
    InMux I__1261 (
            .O(N__6540),
            .I(N__6536));
    InMux I__1260 (
            .O(N__6539),
            .I(N__6533));
    LocalMux I__1259 (
            .O(N__6536),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__1258 (
            .O(N__6533),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__1257 (
            .O(N__6528),
            .I(N__6525));
    LocalMux I__1256 (
            .O(N__6525),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0 ));
    InMux I__1255 (
            .O(N__6522),
            .I(N__6519));
    LocalMux I__1254 (
            .O(N__6519),
            .I(N__6516));
    Span4Mux_v I__1253 (
            .O(N__6516),
            .I(N__6513));
    Sp12to4 I__1252 (
            .O(N__6513),
            .I(N__6510));
    Span12Mux_h I__1251 (
            .O(N__6510),
            .I(N__6507));
    Span12Mux_v I__1250 (
            .O(N__6507),
            .I(N__6504));
    Odrv12 I__1249 (
            .O(N__6504),
            .I(DBRn_c));
    CascadeMux I__1248 (
            .O(N__6501),
            .I(N__6497));
    InMux I__1247 (
            .O(N__6500),
            .I(N__6494));
    InMux I__1246 (
            .O(N__6497),
            .I(N__6489));
    LocalMux I__1245 (
            .O(N__6494),
            .I(N__6486));
    InMux I__1244 (
            .O(N__6493),
            .I(N__6483));
    InMux I__1243 (
            .O(N__6492),
            .I(N__6480));
    LocalMux I__1242 (
            .O(N__6489),
            .I(N__6477));
    Span4Mux_v I__1241 (
            .O(N__6486),
            .I(N__6474));
    LocalMux I__1240 (
            .O(N__6483),
            .I(N__6471));
    LocalMux I__1239 (
            .O(N__6480),
            .I(U712_REG_SM_DBR_SYNC_0));
    Odrv12 I__1238 (
            .O(N__6477),
            .I(U712_REG_SM_DBR_SYNC_0));
    Odrv4 I__1237 (
            .O(N__6474),
            .I(U712_REG_SM_DBR_SYNC_0));
    Odrv4 I__1236 (
            .O(N__6471),
            .I(U712_REG_SM_DBR_SYNC_0));
    InMux I__1235 (
            .O(N__6462),
            .I(N__6459));
    LocalMux I__1234 (
            .O(N__6459),
            .I(\U712_BYTE_ENABLE.UMBE_0 ));
    IoInMux I__1233 (
            .O(N__6456),
            .I(N__6453));
    LocalMux I__1232 (
            .O(N__6453),
            .I(N__6450));
    IoSpan4Mux I__1231 (
            .O(N__6450),
            .I(N__6447));
    Span4Mux_s3_v I__1230 (
            .O(N__6447),
            .I(N__6444));
    Sp12to4 I__1229 (
            .O(N__6444),
            .I(N__6441));
    Span12Mux_v I__1228 (
            .O(N__6441),
            .I(N__6438));
    Span12Mux_h I__1227 (
            .O(N__6438),
            .I(N__6435));
    Odrv12 I__1226 (
            .O(N__6435),
            .I(CUMBEn_c));
    CascadeMux I__1225 (
            .O(N__6432),
            .I(N__6429));
    InMux I__1224 (
            .O(N__6429),
            .I(N__6426));
    LocalMux I__1223 (
            .O(N__6426),
            .I(N__6423));
    Odrv4 I__1222 (
            .O(N__6423),
            .I(\U712_BYTE_ENABLE.UUBE_0 ));
    InMux I__1221 (
            .O(N__6420),
            .I(N__6414));
    InMux I__1220 (
            .O(N__6419),
            .I(N__6414));
    LocalMux I__1219 (
            .O(N__6414),
            .I(\U712_BYTE_ENABLE.un3_CUMBEnZ0Z_0 ));
    IoInMux I__1218 (
            .O(N__6411),
            .I(N__6408));
    LocalMux I__1217 (
            .O(N__6408),
            .I(N__6405));
    IoSpan4Mux I__1216 (
            .O(N__6405),
            .I(N__6402));
    Sp12to4 I__1215 (
            .O(N__6402),
            .I(N__6399));
    Span12Mux_s7_h I__1214 (
            .O(N__6399),
            .I(N__6396));
    Span12Mux_v I__1213 (
            .O(N__6396),
            .I(N__6393));
    Odrv12 I__1212 (
            .O(N__6393),
            .I(CUUBEn_c));
    InMux I__1211 (
            .O(N__6390),
            .I(N__6387));
    LocalMux I__1210 (
            .O(N__6387),
            .I(N__6384));
    Span4Mux_v I__1209 (
            .O(N__6384),
            .I(N__6380));
    InMux I__1208 (
            .O(N__6383),
            .I(N__6377));
    Odrv4 I__1207 (
            .O(N__6380),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    LocalMux I__1206 (
            .O(N__6377),
            .I(\U712_REG_SM.LDS_OUTZ0 ));
    IoInMux I__1205 (
            .O(N__6372),
            .I(N__6369));
    LocalMux I__1204 (
            .O(N__6369),
            .I(N__6366));
    IoSpan4Mux I__1203 (
            .O(N__6366),
            .I(N__6363));
    IoSpan4Mux I__1202 (
            .O(N__6363),
            .I(N__6360));
    Span4Mux_s0_v I__1201 (
            .O(N__6360),
            .I(N__6357));
    Sp12to4 I__1200 (
            .O(N__6357),
            .I(N__6354));
    Span12Mux_v I__1199 (
            .O(N__6354),
            .I(N__6351));
    Odrv12 I__1198 (
            .O(N__6351),
            .I(U712_REG_SM_un1_LDSn_i));
    IoInMux I__1197 (
            .O(N__6348),
            .I(N__6345));
    LocalMux I__1196 (
            .O(N__6345),
            .I(N__6342));
    Span12Mux_s5_h I__1195 (
            .O(N__6342),
            .I(N__6339));
    Span12Mux_h I__1194 (
            .O(N__6339),
            .I(N__6336));
    Odrv12 I__1193 (
            .O(N__6336),
            .I(CMA_c_3));
    InMux I__1192 (
            .O(N__6333),
            .I(N__6330));
    LocalMux I__1191 (
            .O(N__6330),
            .I(N__6327));
    Span4Mux_h I__1190 (
            .O(N__6327),
            .I(N__6324));
    Odrv4 I__1189 (
            .O(N__6324),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    CascadeMux I__1188 (
            .O(N__6321),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_START_2_2_cascade_ ));
    InMux I__1187 (
            .O(N__6318),
            .I(N__6313));
    InMux I__1186 (
            .O(N__6317),
            .I(N__6308));
    InMux I__1185 (
            .O(N__6316),
            .I(N__6308));
    LocalMux I__1184 (
            .O(N__6313),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ));
    LocalMux I__1183 (
            .O(N__6308),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ));
    CascadeMux I__1182 (
            .O(N__6303),
            .I(\U712_CHIP_RAM.REFRESH_CYCLE_0_sqmuxa_cascade_ ));
    InMux I__1181 (
            .O(N__6300),
            .I(N__6297));
    LocalMux I__1180 (
            .O(N__6297),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_0 ));
    InMux I__1179 (
            .O(N__6294),
            .I(N__6288));
    InMux I__1178 (
            .O(N__6293),
            .I(N__6281));
    InMux I__1177 (
            .O(N__6292),
            .I(N__6281));
    InMux I__1176 (
            .O(N__6291),
            .I(N__6281));
    LocalMux I__1175 (
            .O(N__6288),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    LocalMux I__1174 (
            .O(N__6281),
            .I(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ));
    InMux I__1173 (
            .O(N__6276),
            .I(N__6272));
    InMux I__1172 (
            .O(N__6275),
            .I(N__6269));
    LocalMux I__1171 (
            .O(N__6272),
            .I(\U712_CHIP_RAM.N_70_2 ));
    LocalMux I__1170 (
            .O(N__6269),
            .I(\U712_CHIP_RAM.N_70_2 ));
    CascadeMux I__1169 (
            .O(N__6264),
            .I(N__6260));
    CascadeMux I__1168 (
            .O(N__6263),
            .I(N__6253));
    InMux I__1167 (
            .O(N__6260),
            .I(N__6250));
    InMux I__1166 (
            .O(N__6259),
            .I(N__6247));
    InMux I__1165 (
            .O(N__6258),
            .I(N__6244));
    CascadeMux I__1164 (
            .O(N__6257),
            .I(N__6234));
    InMux I__1163 (
            .O(N__6256),
            .I(N__6230));
    InMux I__1162 (
            .O(N__6253),
            .I(N__6227));
    LocalMux I__1161 (
            .O(N__6250),
            .I(N__6220));
    LocalMux I__1160 (
            .O(N__6247),
            .I(N__6220));
    LocalMux I__1159 (
            .O(N__6244),
            .I(N__6220));
    InMux I__1158 (
            .O(N__6243),
            .I(N__6217));
    InMux I__1157 (
            .O(N__6242),
            .I(N__6214));
    InMux I__1156 (
            .O(N__6241),
            .I(N__6207));
    InMux I__1155 (
            .O(N__6240),
            .I(N__6207));
    InMux I__1154 (
            .O(N__6239),
            .I(N__6207));
    InMux I__1153 (
            .O(N__6238),
            .I(N__6204));
    InMux I__1152 (
            .O(N__6237),
            .I(N__6197));
    InMux I__1151 (
            .O(N__6234),
            .I(N__6197));
    InMux I__1150 (
            .O(N__6233),
            .I(N__6197));
    LocalMux I__1149 (
            .O(N__6230),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1148 (
            .O(N__6227),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1147 (
            .O(N__6220),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1146 (
            .O(N__6217),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1145 (
            .O(N__6214),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1144 (
            .O(N__6207),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1143 (
            .O(N__6204),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1142 (
            .O(N__6197),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    CascadeMux I__1141 (
            .O(N__6180),
            .I(N__6175));
    InMux I__1140 (
            .O(N__6179),
            .I(N__6170));
    InMux I__1139 (
            .O(N__6178),
            .I(N__6170));
    InMux I__1138 (
            .O(N__6175),
            .I(N__6167));
    LocalMux I__1137 (
            .O(N__6170),
            .I(\U712_CHIP_RAM.N_106 ));
    LocalMux I__1136 (
            .O(N__6167),
            .I(\U712_CHIP_RAM.N_106 ));
    CascadeMux I__1135 (
            .O(N__6162),
            .I(N__6158));
    InMux I__1134 (
            .O(N__6161),
            .I(N__6152));
    InMux I__1133 (
            .O(N__6158),
            .I(N__6149));
    InMux I__1132 (
            .O(N__6157),
            .I(N__6145));
    InMux I__1131 (
            .O(N__6156),
            .I(N__6142));
    CascadeMux I__1130 (
            .O(N__6155),
            .I(N__6139));
    LocalMux I__1129 (
            .O(N__6152),
            .I(N__6136));
    LocalMux I__1128 (
            .O(N__6149),
            .I(N__6133));
    CascadeMux I__1127 (
            .O(N__6148),
            .I(N__6130));
    LocalMux I__1126 (
            .O(N__6145),
            .I(N__6120));
    LocalMux I__1125 (
            .O(N__6142),
            .I(N__6120));
    InMux I__1124 (
            .O(N__6139),
            .I(N__6117));
    Span4Mux_h I__1123 (
            .O(N__6136),
            .I(N__6112));
    Span4Mux_v I__1122 (
            .O(N__6133),
            .I(N__6112));
    InMux I__1121 (
            .O(N__6130),
            .I(N__6109));
    InMux I__1120 (
            .O(N__6129),
            .I(N__6104));
    InMux I__1119 (
            .O(N__6128),
            .I(N__6104));
    InMux I__1118 (
            .O(N__6127),
            .I(N__6101));
    InMux I__1117 (
            .O(N__6126),
            .I(N__6096));
    InMux I__1116 (
            .O(N__6125),
            .I(N__6096));
    Odrv4 I__1115 (
            .O(N__6120),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1114 (
            .O(N__6117),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1113 (
            .O(N__6112),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1112 (
            .O(N__6109),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1111 (
            .O(N__6104),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1110 (
            .O(N__6101),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1109 (
            .O(N__6096),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    CascadeMux I__1108 (
            .O(N__6081),
            .I(N__6078));
    InMux I__1107 (
            .O(N__6078),
            .I(N__6075));
    LocalMux I__1106 (
            .O(N__6075),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_3_0 ));
    InMux I__1105 (
            .O(N__6072),
            .I(N__6067));
    CascadeMux I__1104 (
            .O(N__6071),
            .I(N__6064));
    InMux I__1103 (
            .O(N__6070),
            .I(N__6061));
    LocalMux I__1102 (
            .O(N__6067),
            .I(N__6058));
    InMux I__1101 (
            .O(N__6064),
            .I(N__6055));
    LocalMux I__1100 (
            .O(N__6061),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    Odrv4 I__1099 (
            .O(N__6058),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__1098 (
            .O(N__6055),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    InMux I__1097 (
            .O(N__6048),
            .I(N__6043));
    InMux I__1096 (
            .O(N__6047),
            .I(N__6038));
    InMux I__1095 (
            .O(N__6046),
            .I(N__6038));
    LocalMux I__1094 (
            .O(N__6043),
            .I(N__6034));
    LocalMux I__1093 (
            .O(N__6038),
            .I(N__6031));
    InMux I__1092 (
            .O(N__6037),
            .I(N__6028));
    Span4Mux_h I__1091 (
            .O(N__6034),
            .I(N__6025));
    Odrv4 I__1090 (
            .O(N__6031),
            .I(\U712_CHIP_RAM.N_40 ));
    LocalMux I__1089 (
            .O(N__6028),
            .I(\U712_CHIP_RAM.N_40 ));
    Odrv4 I__1088 (
            .O(N__6025),
            .I(\U712_CHIP_RAM.N_40 ));
    CascadeMux I__1087 (
            .O(N__6018),
            .I(\U712_CHIP_RAM.N_40_cascade_ ));
    CascadeMux I__1086 (
            .O(N__6015),
            .I(N__6012));
    InMux I__1085 (
            .O(N__6012),
            .I(N__6003));
    InMux I__1084 (
            .O(N__6011),
            .I(N__6000));
    InMux I__1083 (
            .O(N__6010),
            .I(N__5997));
    InMux I__1082 (
            .O(N__6009),
            .I(N__5992));
    InMux I__1081 (
            .O(N__6008),
            .I(N__5992));
    InMux I__1080 (
            .O(N__6007),
            .I(N__5987));
    InMux I__1079 (
            .O(N__6006),
            .I(N__5987));
    LocalMux I__1078 (
            .O(N__6003),
            .I(\U712_CHIP_RAM.N_51 ));
    LocalMux I__1077 (
            .O(N__6000),
            .I(\U712_CHIP_RAM.N_51 ));
    LocalMux I__1076 (
            .O(N__5997),
            .I(\U712_CHIP_RAM.N_51 ));
    LocalMux I__1075 (
            .O(N__5992),
            .I(\U712_CHIP_RAM.N_51 ));
    LocalMux I__1074 (
            .O(N__5987),
            .I(\U712_CHIP_RAM.N_51 ));
    InMux I__1073 (
            .O(N__5976),
            .I(N__5973));
    LocalMux I__1072 (
            .O(N__5973),
            .I(\U712_CHIP_RAM.N_59 ));
    CascadeMux I__1071 (
            .O(N__5970),
            .I(\U712_CHIP_RAM.N_59_cascade_ ));
    InMux I__1070 (
            .O(N__5967),
            .I(N__5962));
    InMux I__1069 (
            .O(N__5966),
            .I(N__5958));
    InMux I__1068 (
            .O(N__5965),
            .I(N__5955));
    LocalMux I__1067 (
            .O(N__5962),
            .I(N__5949));
    InMux I__1066 (
            .O(N__5961),
            .I(N__5946));
    LocalMux I__1065 (
            .O(N__5958),
            .I(N__5941));
    LocalMux I__1064 (
            .O(N__5955),
            .I(N__5941));
    InMux I__1063 (
            .O(N__5954),
            .I(N__5938));
    InMux I__1062 (
            .O(N__5953),
            .I(N__5933));
    InMux I__1061 (
            .O(N__5952),
            .I(N__5933));
    Odrv4 I__1060 (
            .O(N__5949),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0 ));
    LocalMux I__1059 (
            .O(N__5946),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0 ));
    Odrv4 I__1058 (
            .O(N__5941),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0 ));
    LocalMux I__1057 (
            .O(N__5938),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0 ));
    LocalMux I__1056 (
            .O(N__5933),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0 ));
    CascadeMux I__1055 (
            .O(N__5922),
            .I(N__5919));
    InMux I__1054 (
            .O(N__5919),
            .I(N__5906));
    InMux I__1053 (
            .O(N__5918),
            .I(N__5906));
    CascadeMux I__1052 (
            .O(N__5917),
            .I(N__5903));
    InMux I__1051 (
            .O(N__5916),
            .I(N__5898));
    InMux I__1050 (
            .O(N__5915),
            .I(N__5894));
    InMux I__1049 (
            .O(N__5914),
            .I(N__5889));
    InMux I__1048 (
            .O(N__5913),
            .I(N__5889));
    InMux I__1047 (
            .O(N__5912),
            .I(N__5881));
    InMux I__1046 (
            .O(N__5911),
            .I(N__5881));
    LocalMux I__1045 (
            .O(N__5906),
            .I(N__5878));
    InMux I__1044 (
            .O(N__5903),
            .I(N__5875));
    InMux I__1043 (
            .O(N__5902),
            .I(N__5870));
    InMux I__1042 (
            .O(N__5901),
            .I(N__5870));
    LocalMux I__1041 (
            .O(N__5898),
            .I(N__5867));
    InMux I__1040 (
            .O(N__5897),
            .I(N__5864));
    LocalMux I__1039 (
            .O(N__5894),
            .I(N__5861));
    LocalMux I__1038 (
            .O(N__5889),
            .I(N__5858));
    InMux I__1037 (
            .O(N__5888),
            .I(N__5854));
    InMux I__1036 (
            .O(N__5887),
            .I(N__5851));
    InMux I__1035 (
            .O(N__5886),
            .I(N__5848));
    LocalMux I__1034 (
            .O(N__5881),
            .I(N__5841));
    Span4Mux_v I__1033 (
            .O(N__5878),
            .I(N__5841));
    LocalMux I__1032 (
            .O(N__5875),
            .I(N__5841));
    LocalMux I__1031 (
            .O(N__5870),
            .I(N__5834));
    Span4Mux_h I__1030 (
            .O(N__5867),
            .I(N__5834));
    LocalMux I__1029 (
            .O(N__5864),
            .I(N__5834));
    Span4Mux_h I__1028 (
            .O(N__5861),
            .I(N__5831));
    Span4Mux_h I__1027 (
            .O(N__5858),
            .I(N__5828));
    InMux I__1026 (
            .O(N__5857),
            .I(N__5825));
    LocalMux I__1025 (
            .O(N__5854),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1024 (
            .O(N__5851),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1023 (
            .O(N__5848),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1022 (
            .O(N__5841),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1021 (
            .O(N__5834),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1020 (
            .O(N__5831),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1019 (
            .O(N__5828),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1018 (
            .O(N__5825),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1017 (
            .O(N__5808),
            .I(N__5805));
    LocalMux I__1016 (
            .O(N__5805),
            .I(\U712_CYCLE_TERM.N_45_0_0_en ));
    InMux I__1015 (
            .O(N__5802),
            .I(N__5797));
    InMux I__1014 (
            .O(N__5801),
            .I(N__5794));
    InMux I__1013 (
            .O(N__5800),
            .I(N__5791));
    LocalMux I__1012 (
            .O(N__5797),
            .I(\U712_CHIP_RAM.N_46 ));
    LocalMux I__1011 (
            .O(N__5794),
            .I(\U712_CHIP_RAM.N_46 ));
    LocalMux I__1010 (
            .O(N__5791),
            .I(\U712_CHIP_RAM.N_46 ));
    InMux I__1009 (
            .O(N__5784),
            .I(N__5781));
    LocalMux I__1008 (
            .O(N__5781),
            .I(\U712_CHIP_RAM.N_77 ));
    InMux I__1007 (
            .O(N__5778),
            .I(N__5774));
    InMux I__1006 (
            .O(N__5777),
            .I(N__5771));
    LocalMux I__1005 (
            .O(N__5774),
            .I(\U712_CHIP_RAM.N_99 ));
    LocalMux I__1004 (
            .O(N__5771),
            .I(\U712_CHIP_RAM.N_99 ));
    CascadeMux I__1003 (
            .O(N__5766),
            .I(\U712_CHIP_RAM.N_99_cascade_ ));
    InMux I__1002 (
            .O(N__5763),
            .I(N__5760));
    LocalMux I__1001 (
            .O(N__5760),
            .I(\U712_CHIP_RAM.N_79 ));
    InMux I__1000 (
            .O(N__5757),
            .I(N__5751));
    InMux I__999 (
            .O(N__5756),
            .I(N__5751));
    LocalMux I__998 (
            .O(N__5751),
            .I(\U712_CHIP_RAM.N_93_1 ));
    InMux I__997 (
            .O(N__5748),
            .I(N__5744));
    InMux I__996 (
            .O(N__5747),
            .I(N__5741));
    LocalMux I__995 (
            .O(N__5744),
            .I(\U712_CHIP_RAM.N_52 ));
    LocalMux I__994 (
            .O(N__5741),
            .I(\U712_CHIP_RAM.N_52 ));
    InMux I__993 (
            .O(N__5736),
            .I(N__5727));
    InMux I__992 (
            .O(N__5735),
            .I(N__5724));
    InMux I__991 (
            .O(N__5734),
            .I(N__5721));
    InMux I__990 (
            .O(N__5733),
            .I(N__5718));
    InMux I__989 (
            .O(N__5732),
            .I(N__5713));
    InMux I__988 (
            .O(N__5731),
            .I(N__5713));
    InMux I__987 (
            .O(N__5730),
            .I(N__5710));
    LocalMux I__986 (
            .O(N__5727),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__985 (
            .O(N__5724),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__984 (
            .O(N__5721),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__983 (
            .O(N__5718),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__982 (
            .O(N__5713),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__981 (
            .O(N__5710),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__980 (
            .O(N__5697),
            .I(N__5694));
    LocalMux I__979 (
            .O(N__5694),
            .I(N__5690));
    InMux I__978 (
            .O(N__5693),
            .I(N__5687));
    Odrv4 I__977 (
            .O(N__5690),
            .I(\U712_CHIP_RAM.N_54 ));
    LocalMux I__976 (
            .O(N__5687),
            .I(\U712_CHIP_RAM.N_54 ));
    CascadeMux I__975 (
            .O(N__5682),
            .I(N__5674));
    CascadeMux I__974 (
            .O(N__5681),
            .I(N__5671));
    InMux I__973 (
            .O(N__5680),
            .I(N__5667));
    InMux I__972 (
            .O(N__5679),
            .I(N__5664));
    InMux I__971 (
            .O(N__5678),
            .I(N__5661));
    InMux I__970 (
            .O(N__5677),
            .I(N__5656));
    InMux I__969 (
            .O(N__5674),
            .I(N__5656));
    InMux I__968 (
            .O(N__5671),
            .I(N__5651));
    InMux I__967 (
            .O(N__5670),
            .I(N__5651));
    LocalMux I__966 (
            .O(N__5667),
            .I(N__5648));
    LocalMux I__965 (
            .O(N__5664),
            .I(\U712_CHIP_RAM.N_50 ));
    LocalMux I__964 (
            .O(N__5661),
            .I(\U712_CHIP_RAM.N_50 ));
    LocalMux I__963 (
            .O(N__5656),
            .I(\U712_CHIP_RAM.N_50 ));
    LocalMux I__962 (
            .O(N__5651),
            .I(\U712_CHIP_RAM.N_50 ));
    Odrv4 I__961 (
            .O(N__5648),
            .I(\U712_CHIP_RAM.N_50 ));
    CascadeMux I__960 (
            .O(N__5637),
            .I(\U712_CHIP_RAM.N_54_cascade_ ));
    InMux I__959 (
            .O(N__5634),
            .I(N__5624));
    InMux I__958 (
            .O(N__5633),
            .I(N__5624));
    InMux I__957 (
            .O(N__5632),
            .I(N__5621));
    InMux I__956 (
            .O(N__5631),
            .I(N__5608));
    InMux I__955 (
            .O(N__5630),
            .I(N__5603));
    InMux I__954 (
            .O(N__5629),
            .I(N__5603));
    LocalMux I__953 (
            .O(N__5624),
            .I(N__5598));
    LocalMux I__952 (
            .O(N__5621),
            .I(N__5598));
    InMux I__951 (
            .O(N__5620),
            .I(N__5595));
    InMux I__950 (
            .O(N__5619),
            .I(N__5590));
    InMux I__949 (
            .O(N__5618),
            .I(N__5590));
    InMux I__948 (
            .O(N__5617),
            .I(N__5583));
    InMux I__947 (
            .O(N__5616),
            .I(N__5583));
    InMux I__946 (
            .O(N__5615),
            .I(N__5583));
    InMux I__945 (
            .O(N__5614),
            .I(N__5574));
    InMux I__944 (
            .O(N__5613),
            .I(N__5574));
    InMux I__943 (
            .O(N__5612),
            .I(N__5574));
    InMux I__942 (
            .O(N__5611),
            .I(N__5574));
    LocalMux I__941 (
            .O(N__5608),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__940 (
            .O(N__5603),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__939 (
            .O(N__5598),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__938 (
            .O(N__5595),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__937 (
            .O(N__5590),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__936 (
            .O(N__5583),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__935 (
            .O(N__5574),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__934 (
            .O(N__5559),
            .I(N__5556));
    LocalMux I__933 (
            .O(N__5556),
            .I(N__5553));
    Span4Mux_v I__932 (
            .O(N__5553),
            .I(N__5550));
    Sp12to4 I__931 (
            .O(N__5550),
            .I(N__5547));
    Span12Mux_h I__930 (
            .O(N__5547),
            .I(N__5544));
    Odrv12 I__929 (
            .O(N__5544),
            .I(A_c_11));
    CascadeMux I__928 (
            .O(N__5541),
            .I(\U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_ ));
    InMux I__927 (
            .O(N__5538),
            .I(N__5535));
    LocalMux I__926 (
            .O(N__5535),
            .I(N__5532));
    Span12Mux_v I__925 (
            .O(N__5532),
            .I(N__5529));
    Span12Mux_h I__924 (
            .O(N__5529),
            .I(N__5526));
    Odrv12 I__923 (
            .O(N__5526),
            .I(A_c_4));
    SRMux I__922 (
            .O(N__5523),
            .I(N__5520));
    LocalMux I__921 (
            .O(N__5520),
            .I(N__5517));
    Span4Mux_h I__920 (
            .O(N__5517),
            .I(N__5514));
    Odrv4 I__919 (
            .O(N__5514),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    CascadeMux I__918 (
            .O(N__5511),
            .I(\U712_CHIP_RAM.N_78_cascade_ ));
    CascadeMux I__917 (
            .O(N__5508),
            .I(\U712_CHIP_RAM.N_76_cascade_ ));
    InMux I__916 (
            .O(N__5505),
            .I(N__5499));
    InMux I__915 (
            .O(N__5504),
            .I(N__5499));
    LocalMux I__914 (
            .O(N__5499),
            .I(\U712_CHIP_RAM.N_58 ));
    InMux I__913 (
            .O(N__5496),
            .I(N__5490));
    InMux I__912 (
            .O(N__5495),
            .I(N__5483));
    InMux I__911 (
            .O(N__5494),
            .I(N__5483));
    InMux I__910 (
            .O(N__5493),
            .I(N__5483));
    LocalMux I__909 (
            .O(N__5490),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ));
    LocalMux I__908 (
            .O(N__5483),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ));
    InMux I__907 (
            .O(N__5478),
            .I(N__5474));
    InMux I__906 (
            .O(N__5477),
            .I(N__5471));
    LocalMux I__905 (
            .O(N__5474),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c2 ));
    LocalMux I__904 (
            .O(N__5471),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c2 ));
    InMux I__903 (
            .O(N__5466),
            .I(N__5463));
    LocalMux I__902 (
            .O(N__5463),
            .I(\U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1 ));
    CascadeMux I__901 (
            .O(N__5460),
            .I(\U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1_cascade_ ));
    IoInMux I__900 (
            .O(N__5457),
            .I(N__5454));
    LocalMux I__899 (
            .O(N__5454),
            .I(N__5451));
    IoSpan4Mux I__898 (
            .O(N__5451),
            .I(N__5448));
    Span4Mux_s2_v I__897 (
            .O(N__5448),
            .I(N__5445));
    Sp12to4 I__896 (
            .O(N__5445),
            .I(N__5442));
    Span12Mux_v I__895 (
            .O(N__5442),
            .I(N__5439));
    Odrv12 I__894 (
            .O(N__5439),
            .I(CLLBEn_c));
    IoInMux I__893 (
            .O(N__5436),
            .I(N__5433));
    LocalMux I__892 (
            .O(N__5433),
            .I(N__5430));
    Span4Mux_s1_v I__891 (
            .O(N__5430),
            .I(N__5427));
    Sp12to4 I__890 (
            .O(N__5427),
            .I(N__5424));
    Span12Mux_h I__889 (
            .O(N__5424),
            .I(N__5419));
    InMux I__888 (
            .O(N__5423),
            .I(N__5414));
    InMux I__887 (
            .O(N__5422),
            .I(N__5414));
    Span12Mux_v I__886 (
            .O(N__5419),
            .I(N__5410));
    LocalMux I__885 (
            .O(N__5414),
            .I(N__5407));
    InMux I__884 (
            .O(N__5413),
            .I(N__5404));
    Odrv12 I__883 (
            .O(N__5410),
            .I(DBENn_c));
    Odrv4 I__882 (
            .O(N__5407),
            .I(DBENn_c));
    LocalMux I__881 (
            .O(N__5404),
            .I(DBENn_c));
    InMux I__880 (
            .O(N__5397),
            .I(N__5391));
    InMux I__879 (
            .O(N__5396),
            .I(N__5388));
    InMux I__878 (
            .O(N__5395),
            .I(N__5385));
    InMux I__877 (
            .O(N__5394),
            .I(N__5382));
    LocalMux I__876 (
            .O(N__5391),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    LocalMux I__875 (
            .O(N__5388),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    LocalMux I__874 (
            .O(N__5385),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    LocalMux I__873 (
            .O(N__5382),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_5 ));
    CascadeMux I__872 (
            .O(N__5373),
            .I(N__5370));
    InMux I__871 (
            .O(N__5370),
            .I(N__5367));
    LocalMux I__870 (
            .O(N__5367),
            .I(N__5362));
    InMux I__869 (
            .O(N__5366),
            .I(N__5357));
    InMux I__868 (
            .O(N__5365),
            .I(N__5357));
    Span4Mux_h I__867 (
            .O(N__5362),
            .I(N__5354));
    LocalMux I__866 (
            .O(N__5357),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    Odrv4 I__865 (
            .O(N__5354),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_3 ));
    InMux I__864 (
            .O(N__5349),
            .I(N__5345));
    InMux I__863 (
            .O(N__5348),
            .I(N__5342));
    LocalMux I__862 (
            .O(N__5345),
            .I(\U712_REG_SM.N_167_0 ));
    LocalMux I__861 (
            .O(N__5342),
            .I(\U712_REG_SM.N_167_0 ));
    InMux I__860 (
            .O(N__5337),
            .I(N__5334));
    LocalMux I__859 (
            .O(N__5334),
            .I(N__5331));
    Odrv12 I__858 (
            .O(N__5331),
            .I(\U712_BYTE_ENABLE.LLBE_0 ));
    CascadeMux I__857 (
            .O(N__5328),
            .I(N__5325));
    InMux I__856 (
            .O(N__5325),
            .I(N__5322));
    LocalMux I__855 (
            .O(N__5322),
            .I(N__5319));
    Odrv4 I__854 (
            .O(N__5319),
            .I(\U712_BYTE_ENABLE.LMBE_0 ));
    InMux I__853 (
            .O(N__5316),
            .I(N__5310));
    InMux I__852 (
            .O(N__5315),
            .I(N__5305));
    InMux I__851 (
            .O(N__5314),
            .I(N__5305));
    InMux I__850 (
            .O(N__5313),
            .I(N__5302));
    LocalMux I__849 (
            .O(N__5310),
            .I(N__5295));
    LocalMux I__848 (
            .O(N__5305),
            .I(N__5295));
    LocalMux I__847 (
            .O(N__5302),
            .I(N__5295));
    Span4Mux_v I__846 (
            .O(N__5295),
            .I(N__5292));
    Span4Mux_v I__845 (
            .O(N__5292),
            .I(N__5287));
    InMux I__844 (
            .O(N__5291),
            .I(N__5282));
    InMux I__843 (
            .O(N__5290),
            .I(N__5282));
    Span4Mux_v I__842 (
            .O(N__5287),
            .I(N__5279));
    LocalMux I__841 (
            .O(N__5282),
            .I(N__5276));
    Sp12to4 I__840 (
            .O(N__5279),
            .I(N__5271));
    Span12Mux_v I__839 (
            .O(N__5276),
            .I(N__5271));
    Odrv12 I__838 (
            .O(N__5271),
            .I(SIZ_c_0));
    CascadeMux I__837 (
            .O(N__5268),
            .I(N__5265));
    InMux I__836 (
            .O(N__5265),
            .I(N__5255));
    InMux I__835 (
            .O(N__5264),
            .I(N__5255));
    InMux I__834 (
            .O(N__5263),
            .I(N__5255));
    InMux I__833 (
            .O(N__5262),
            .I(N__5252));
    LocalMux I__832 (
            .O(N__5255),
            .I(N__5247));
    LocalMux I__831 (
            .O(N__5252),
            .I(N__5247));
    Span4Mux_v I__830 (
            .O(N__5247),
            .I(N__5244));
    Span4Mux_v I__829 (
            .O(N__5244),
            .I(N__5241));
    Sp12to4 I__828 (
            .O(N__5241),
            .I(N__5238));
    Odrv12 I__827 (
            .O(N__5238),
            .I(A_c_1));
    CascadeMux I__826 (
            .O(N__5235),
            .I(N__5229));
    CascadeMux I__825 (
            .O(N__5234),
            .I(N__5226));
    CascadeMux I__824 (
            .O(N__5233),
            .I(N__5223));
    InMux I__823 (
            .O(N__5232),
            .I(N__5214));
    InMux I__822 (
            .O(N__5229),
            .I(N__5214));
    InMux I__821 (
            .O(N__5226),
            .I(N__5214));
    InMux I__820 (
            .O(N__5223),
            .I(N__5211));
    InMux I__819 (
            .O(N__5222),
            .I(N__5206));
    InMux I__818 (
            .O(N__5221),
            .I(N__5206));
    LocalMux I__817 (
            .O(N__5214),
            .I(N__5199));
    LocalMux I__816 (
            .O(N__5211),
            .I(N__5199));
    LocalMux I__815 (
            .O(N__5206),
            .I(N__5199));
    Span4Mux_v I__814 (
            .O(N__5199),
            .I(N__5196));
    Sp12to4 I__813 (
            .O(N__5196),
            .I(N__5193));
    Odrv12 I__812 (
            .O(N__5193),
            .I(A_c_0));
    InMux I__811 (
            .O(N__5190),
            .I(N__5187));
    LocalMux I__810 (
            .O(N__5187),
            .I(N__5184));
    Span4Mux_v I__809 (
            .O(N__5184),
            .I(N__5178));
    InMux I__808 (
            .O(N__5183),
            .I(N__5173));
    InMux I__807 (
            .O(N__5182),
            .I(N__5173));
    InMux I__806 (
            .O(N__5181),
            .I(N__5170));
    Span4Mux_v I__805 (
            .O(N__5178),
            .I(N__5167));
    LocalMux I__804 (
            .O(N__5173),
            .I(N__5162));
    LocalMux I__803 (
            .O(N__5170),
            .I(N__5162));
    Span4Mux_v I__802 (
            .O(N__5167),
            .I(N__5159));
    Sp12to4 I__801 (
            .O(N__5162),
            .I(N__5156));
    Sp12to4 I__800 (
            .O(N__5159),
            .I(N__5151));
    Span12Mux_v I__799 (
            .O(N__5156),
            .I(N__5151));
    Span12Mux_h I__798 (
            .O(N__5151),
            .I(N__5148));
    Odrv12 I__797 (
            .O(N__5148),
            .I(SIZ_c_1));
    CascadeMux I__796 (
            .O(N__5145),
            .I(N__5141));
    CascadeMux I__795 (
            .O(N__5144),
            .I(N__5138));
    InMux I__794 (
            .O(N__5141),
            .I(N__5134));
    InMux I__793 (
            .O(N__5138),
            .I(N__5129));
    InMux I__792 (
            .O(N__5137),
            .I(N__5129));
    LocalMux I__791 (
            .O(N__5134),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__790 (
            .O(N__5129),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    InMux I__789 (
            .O(N__5124),
            .I(N__5121));
    LocalMux I__788 (
            .O(N__5121),
            .I(\U712_CYCLE_TERM.N_49 ));
    CascadeMux I__787 (
            .O(N__5118),
            .I(N__5114));
    CascadeMux I__786 (
            .O(N__5117),
            .I(N__5111));
    InMux I__785 (
            .O(N__5114),
            .I(N__5107));
    InMux I__784 (
            .O(N__5111),
            .I(N__5102));
    InMux I__783 (
            .O(N__5110),
            .I(N__5102));
    LocalMux I__782 (
            .O(N__5107),
            .I(REG_TACK));
    LocalMux I__781 (
            .O(N__5102),
            .I(REG_TACK));
    InMux I__780 (
            .O(N__5097),
            .I(N__5090));
    InMux I__779 (
            .O(N__5096),
            .I(N__5090));
    InMux I__778 (
            .O(N__5095),
            .I(N__5087));
    LocalMux I__777 (
            .O(N__5090),
            .I(N__5084));
    LocalMux I__776 (
            .O(N__5087),
            .I(CPU_TACKm));
    Odrv4 I__775 (
            .O(N__5084),
            .I(CPU_TACKm));
    CascadeMux I__774 (
            .O(N__5079),
            .I(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ));
    InMux I__773 (
            .O(N__5076),
            .I(N__5073));
    LocalMux I__772 (
            .O(N__5073),
            .I(N__5068));
    InMux I__771 (
            .O(N__5072),
            .I(N__5065));
    CascadeMux I__770 (
            .O(N__5071),
            .I(N__5061));
    Span4Mux_h I__769 (
            .O(N__5068),
            .I(N__5056));
    LocalMux I__768 (
            .O(N__5065),
            .I(N__5056));
    InMux I__767 (
            .O(N__5064),
            .I(N__5051));
    InMux I__766 (
            .O(N__5061),
            .I(N__5051));
    Span4Mux_h I__765 (
            .O(N__5056),
            .I(N__5046));
    LocalMux I__764 (
            .O(N__5051),
            .I(N__5046));
    Span4Mux_h I__763 (
            .O(N__5046),
            .I(N__5043));
    Span4Mux_v I__762 (
            .O(N__5043),
            .I(N__5040));
    Span4Mux_v I__761 (
            .O(N__5040),
            .I(N__5037));
    Span4Mux_v I__760 (
            .O(N__5037),
            .I(N__5034));
    Odrv4 I__759 (
            .O(N__5034),
            .I(CLK40_OUT_i));
    InMux I__758 (
            .O(N__5031),
            .I(N__5025));
    InMux I__757 (
            .O(N__5030),
            .I(N__5025));
    LocalMux I__756 (
            .O(N__5025),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    IoInMux I__755 (
            .O(N__5022),
            .I(N__5019));
    LocalMux I__754 (
            .O(N__5019),
            .I(N__5016));
    IoSpan4Mux I__753 (
            .O(N__5016),
            .I(N__5012));
    InMux I__752 (
            .O(N__5015),
            .I(N__5009));
    Sp12to4 I__751 (
            .O(N__5012),
            .I(N__5005));
    LocalMux I__750 (
            .O(N__5009),
            .I(N__5002));
    CascadeMux I__749 (
            .O(N__5008),
            .I(N__4999));
    Span12Mux_s9_v I__748 (
            .O(N__5005),
            .I(N__4996));
    Span4Mux_v I__747 (
            .O(N__5002),
            .I(N__4993));
    InMux I__746 (
            .O(N__4999),
            .I(N__4990));
    Odrv12 I__745 (
            .O(N__4996),
            .I(DBDIR_c));
    Odrv4 I__744 (
            .O(N__4993),
            .I(DBDIR_c));
    LocalMux I__743 (
            .O(N__4990),
            .I(DBDIR_c));
    IoInMux I__742 (
            .O(N__4983),
            .I(N__4980));
    LocalMux I__741 (
            .O(N__4980),
            .I(N__4977));
    Span4Mux_s3_h I__740 (
            .O(N__4977),
            .I(N__4974));
    Span4Mux_h I__739 (
            .O(N__4974),
            .I(N__4971));
    Sp12to4 I__738 (
            .O(N__4971),
            .I(N__4968));
    Span12Mux_s6_v I__737 (
            .O(N__4968),
            .I(N__4965));
    Span12Mux_h I__736 (
            .O(N__4965),
            .I(N__4962));
    Odrv12 I__735 (
            .O(N__4962),
            .I(DRDDIR_0_i));
    IoInMux I__734 (
            .O(N__4959),
            .I(N__4956));
    LocalMux I__733 (
            .O(N__4956),
            .I(N__4953));
    IoSpan4Mux I__732 (
            .O(N__4953),
            .I(N__4950));
    Span4Mux_s0_h I__731 (
            .O(N__4950),
            .I(N__4947));
    Sp12to4 I__730 (
            .O(N__4947),
            .I(N__4944));
    Span12Mux_h I__729 (
            .O(N__4944),
            .I(N__4941));
    Span12Mux_v I__728 (
            .O(N__4941),
            .I(N__4938));
    Odrv12 I__727 (
            .O(N__4938),
            .I(CLMBEn_c));
    CascadeMux I__726 (
            .O(N__4935),
            .I(\U712_CHIP_RAM.N_106_cascade_ ));
    CascadeMux I__725 (
            .O(N__4932),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_ ));
    CascadeMux I__724 (
            .O(N__4929),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_cascade_ ));
    IoInMux I__723 (
            .O(N__4926),
            .I(N__4923));
    LocalMux I__722 (
            .O(N__4923),
            .I(N__4920));
    IoSpan4Mux I__721 (
            .O(N__4920),
            .I(N__4917));
    Sp12to4 I__720 (
            .O(N__4917),
            .I(N__4914));
    Span12Mux_s7_h I__719 (
            .O(N__4914),
            .I(N__4911));
    Span12Mux_h I__718 (
            .O(N__4911),
            .I(N__4907));
    InMux I__717 (
            .O(N__4910),
            .I(N__4904));
    Odrv12 I__716 (
            .O(N__4907),
            .I(CLK_EN_c));
    LocalMux I__715 (
            .O(N__4904),
            .I(CLK_EN_c));
    InMux I__714 (
            .O(N__4899),
            .I(N__4895));
    InMux I__713 (
            .O(N__4898),
            .I(N__4891));
    LocalMux I__712 (
            .O(N__4895),
            .I(N__4888));
    InMux I__711 (
            .O(N__4894),
            .I(N__4885));
    LocalMux I__710 (
            .O(N__4891),
            .I(\U712_CHIP_RAM.N_100 ));
    Odrv4 I__709 (
            .O(N__4888),
            .I(\U712_CHIP_RAM.N_100 ));
    LocalMux I__708 (
            .O(N__4885),
            .I(\U712_CHIP_RAM.N_100 ));
    CascadeMux I__707 (
            .O(N__4878),
            .I(N__4875));
    InMux I__706 (
            .O(N__4875),
            .I(N__4872));
    LocalMux I__705 (
            .O(N__4872),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0 ));
    InMux I__704 (
            .O(N__4869),
            .I(N__4863));
    InMux I__703 (
            .O(N__4868),
            .I(N__4863));
    LocalMux I__702 (
            .O(N__4863),
            .I(N__4860));
    Odrv4 I__701 (
            .O(N__4860),
            .I(\U712_CHIP_RAM.CPU_TACK_6 ));
    InMux I__700 (
            .O(N__4857),
            .I(N__4854));
    LocalMux I__699 (
            .O(N__4854),
            .I(N__4851));
    Span12Mux_h I__698 (
            .O(N__4851),
            .I(N__4848));
    Span12Mux_v I__697 (
            .O(N__4848),
            .I(N__4845));
    Span12Mux_h I__696 (
            .O(N__4845),
            .I(N__4842));
    Odrv12 I__695 (
            .O(N__4842),
            .I(RAMSPACEn_c));
    CascadeMux I__694 (
            .O(N__4839),
            .I(\U712_CHIP_RAM.un6_CPU_CYCLE_START_cascade_ ));
    InMux I__693 (
            .O(N__4836),
            .I(N__4833));
    LocalMux I__692 (
            .O(N__4833),
            .I(N__4829));
    InMux I__691 (
            .O(N__4832),
            .I(N__4826));
    Span4Mux_v I__690 (
            .O(N__4829),
            .I(N__4823));
    LocalMux I__689 (
            .O(N__4826),
            .I(N__4820));
    Span4Mux_h I__688 (
            .O(N__4823),
            .I(N__4817));
    Span12Mux_h I__687 (
            .O(N__4820),
            .I(N__4814));
    Sp12to4 I__686 (
            .O(N__4817),
            .I(N__4811));
    Span12Mux_v I__685 (
            .O(N__4814),
            .I(N__4808));
    Span12Mux_v I__684 (
            .O(N__4811),
            .I(N__4805));
    Odrv12 I__683 (
            .O(N__4808),
            .I(TSn_c));
    Odrv12 I__682 (
            .O(N__4805),
            .I(TSn_c));
    InMux I__681 (
            .O(N__4800),
            .I(N__4796));
    InMux I__680 (
            .O(N__4799),
            .I(N__4793));
    LocalMux I__679 (
            .O(N__4796),
            .I(N__4790));
    LocalMux I__678 (
            .O(N__4793),
            .I(\U712_CHIP_RAM.N_68 ));
    Odrv4 I__677 (
            .O(N__4790),
            .I(\U712_CHIP_RAM.N_68 ));
    InMux I__676 (
            .O(N__4785),
            .I(N__4781));
    InMux I__675 (
            .O(N__4784),
            .I(N__4778));
    LocalMux I__674 (
            .O(N__4781),
            .I(\U712_CHIP_RAM.N_98 ));
    LocalMux I__673 (
            .O(N__4778),
            .I(\U712_CHIP_RAM.N_98 ));
    CascadeMux I__672 (
            .O(N__4773),
            .I(\U712_CHIP_RAM.N_55_cascade_ ));
    CascadeMux I__671 (
            .O(N__4770),
            .I(\U712_CHIP_RAM.N_57_cascade_ ));
    CascadeMux I__670 (
            .O(N__4767),
            .I(\U712_CHIP_RAM.N_92_cascade_ ));
    InMux I__669 (
            .O(N__4764),
            .I(N__4760));
    InMux I__668 (
            .O(N__4763),
            .I(N__4757));
    LocalMux I__667 (
            .O(N__4760),
            .I(\U712_CHIP_RAM.N_44 ));
    LocalMux I__666 (
            .O(N__4757),
            .I(\U712_CHIP_RAM.N_44 ));
    InMux I__665 (
            .O(N__4752),
            .I(N__4745));
    InMux I__664 (
            .O(N__4751),
            .I(N__4736));
    InMux I__663 (
            .O(N__4750),
            .I(N__4736));
    InMux I__662 (
            .O(N__4749),
            .I(N__4736));
    InMux I__661 (
            .O(N__4748),
            .I(N__4736));
    LocalMux I__660 (
            .O(N__4745),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__659 (
            .O(N__4736),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__658 (
            .O(N__4731),
            .I(N__4725));
    InMux I__657 (
            .O(N__4730),
            .I(N__4725));
    LocalMux I__656 (
            .O(N__4725),
            .I(\U712_CHIP_RAM.BANK0_0_sqmuxa_3 ));
    InMux I__655 (
            .O(N__4722),
            .I(N__4719));
    LocalMux I__654 (
            .O(N__4719),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER17_1 ));
    CascadeMux I__653 (
            .O(N__4716),
            .I(\U712_CHIP_RAM.N_50_cascade_ ));
    InMux I__652 (
            .O(N__4713),
            .I(N__4708));
    InMux I__651 (
            .O(N__4712),
            .I(N__4705));
    InMux I__650 (
            .O(N__4711),
            .I(N__4702));
    LocalMux I__649 (
            .O(N__4708),
            .I(\U712_CHIP_RAM.N_43 ));
    LocalMux I__648 (
            .O(N__4705),
            .I(\U712_CHIP_RAM.N_43 ));
    LocalMux I__647 (
            .O(N__4702),
            .I(\U712_CHIP_RAM.N_43 ));
    CascadeMux I__646 (
            .O(N__4695),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_tz_1_cascade_ ));
    CascadeMux I__645 (
            .O(N__4692),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_ ));
    InMux I__644 (
            .O(N__4689),
            .I(N__4686));
    LocalMux I__643 (
            .O(N__4686),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ));
    CascadeMux I__642 (
            .O(N__4683),
            .I(\U712_REG_SM.N_165_0_cascade_ ));
    InMux I__641 (
            .O(N__4680),
            .I(N__4677));
    LocalMux I__640 (
            .O(N__4677),
            .I(\U712_REG_SM.N_170_0 ));
    CascadeMux I__639 (
            .O(N__4674),
            .I(N__4667));
    InMux I__638 (
            .O(N__4673),
            .I(N__4664));
    InMux I__637 (
            .O(N__4672),
            .I(N__4661));
    InMux I__636 (
            .O(N__4671),
            .I(N__4656));
    InMux I__635 (
            .O(N__4670),
            .I(N__4656));
    InMux I__634 (
            .O(N__4667),
            .I(N__4653));
    LocalMux I__633 (
            .O(N__4664),
            .I(N__4650));
    LocalMux I__632 (
            .O(N__4661),
            .I(N__4647));
    LocalMux I__631 (
            .O(N__4656),
            .I(\U712_REG_SM.N_173_0 ));
    LocalMux I__630 (
            .O(N__4653),
            .I(\U712_REG_SM.N_173_0 ));
    Odrv4 I__629 (
            .O(N__4650),
            .I(\U712_REG_SM.N_173_0 ));
    Odrv4 I__628 (
            .O(N__4647),
            .I(\U712_REG_SM.N_173_0 ));
    InMux I__627 (
            .O(N__4638),
            .I(N__4635));
    LocalMux I__626 (
            .O(N__4635),
            .I(\U712_REG_SM.LDS_OUT_2_0_0 ));
    InMux I__625 (
            .O(N__4632),
            .I(N__4629));
    LocalMux I__624 (
            .O(N__4629),
            .I(\U712_REG_SM.UDS_OUT_2_0_0 ));
    CascadeMux I__623 (
            .O(N__4626),
            .I(\U712_CHIP_RAM.N_105_cascade_ ));
    CascadeMux I__622 (
            .O(N__4623),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_1_1_cascade_ ));
    InMux I__621 (
            .O(N__4620),
            .I(N__4617));
    LocalMux I__620 (
            .O(N__4617),
            .I(\U712_CHIP_RAM.N_105 ));
    CascadeMux I__619 (
            .O(N__4614),
            .I(\U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_1_cascade_ ));
    CascadeMux I__618 (
            .O(N__4611),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_cascade_ ));
    IoInMux I__617 (
            .O(N__4608),
            .I(N__4605));
    LocalMux I__616 (
            .O(N__4605),
            .I(N__4602));
    Span4Mux_s2_h I__615 (
            .O(N__4602),
            .I(N__4599));
    Sp12to4 I__614 (
            .O(N__4599),
            .I(N__4596));
    Span12Mux_v I__613 (
            .O(N__4596),
            .I(N__4592));
    InMux I__612 (
            .O(N__4595),
            .I(N__4589));
    Odrv12 I__611 (
            .O(N__4592),
            .I(TACK_OUTn));
    LocalMux I__610 (
            .O(N__4589),
            .I(TACK_OUTn));
    InMux I__609 (
            .O(N__4584),
            .I(N__4581));
    LocalMux I__608 (
            .O(N__4581),
            .I(N__4578));
    Odrv4 I__607 (
            .O(N__4578),
            .I(\U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1 ));
    CascadeMux I__606 (
            .O(N__4575),
            .I(N__4572));
    InMux I__605 (
            .O(N__4572),
            .I(N__4569));
    LocalMux I__604 (
            .O(N__4569),
            .I(\U712_REG_SM.DS_EN_7_0 ));
    InMux I__603 (
            .O(N__4566),
            .I(N__4563));
    LocalMux I__602 (
            .O(N__4563),
            .I(\U712_REG_SM.N_187 ));
    InMux I__601 (
            .O(N__4560),
            .I(N__4556));
    InMux I__600 (
            .O(N__4559),
            .I(N__4553));
    LocalMux I__599 (
            .O(N__4556),
            .I(\U712_REG_SM.N_157_0 ));
    LocalMux I__598 (
            .O(N__4553),
            .I(\U712_REG_SM.N_157_0 ));
    InMux I__597 (
            .O(N__4548),
            .I(N__4541));
    InMux I__596 (
            .O(N__4547),
            .I(N__4532));
    InMux I__595 (
            .O(N__4546),
            .I(N__4532));
    InMux I__594 (
            .O(N__4545),
            .I(N__4532));
    InMux I__593 (
            .O(N__4544),
            .I(N__4532));
    LocalMux I__592 (
            .O(N__4541),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    LocalMux I__591 (
            .O(N__4532),
            .I(\U712_REG_SM.C3_SYNCZ0Z_2 ));
    InMux I__590 (
            .O(N__4527),
            .I(N__4524));
    LocalMux I__589 (
            .O(N__4524),
            .I(N__4519));
    InMux I__588 (
            .O(N__4523),
            .I(N__4516));
    CascadeMux I__587 (
            .O(N__4522),
            .I(N__4513));
    Span4Mux_v I__586 (
            .O(N__4519),
            .I(N__4505));
    LocalMux I__585 (
            .O(N__4516),
            .I(N__4505));
    InMux I__584 (
            .O(N__4513),
            .I(N__4496));
    InMux I__583 (
            .O(N__4512),
            .I(N__4496));
    InMux I__582 (
            .O(N__4511),
            .I(N__4496));
    InMux I__581 (
            .O(N__4510),
            .I(N__4496));
    Odrv4 I__580 (
            .O(N__4505),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__579 (
            .O(N__4496),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__578 (
            .O(N__4491),
            .I(N__4486));
    InMux I__577 (
            .O(N__4490),
            .I(N__4483));
    InMux I__576 (
            .O(N__4489),
            .I(N__4480));
    LocalMux I__575 (
            .O(N__4486),
            .I(\U712_REG_SM.N_159_0 ));
    LocalMux I__574 (
            .O(N__4483),
            .I(\U712_REG_SM.N_159_0 ));
    LocalMux I__573 (
            .O(N__4480),
            .I(\U712_REG_SM.N_159_0 ));
    CascadeMux I__572 (
            .O(N__4473),
            .I(\U712_REG_SM.N_159_0_cascade_ ));
    InMux I__571 (
            .O(N__4470),
            .I(N__4465));
    InMux I__570 (
            .O(N__4469),
            .I(N__4462));
    InMux I__569 (
            .O(N__4468),
            .I(N__4459));
    LocalMux I__568 (
            .O(N__4465),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__567 (
            .O(N__4462),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    LocalMux I__566 (
            .O(N__4459),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_4 ));
    InMux I__565 (
            .O(N__4452),
            .I(N__4449));
    LocalMux I__564 (
            .O(N__4449),
            .I(\U712_REG_SM.N_165_0 ));
    InMux I__563 (
            .O(N__4446),
            .I(N__4437));
    InMux I__562 (
            .O(N__4445),
            .I(N__4437));
    InMux I__561 (
            .O(N__4444),
            .I(N__4430));
    InMux I__560 (
            .O(N__4443),
            .I(N__4430));
    InMux I__559 (
            .O(N__4442),
            .I(N__4430));
    LocalMux I__558 (
            .O(N__4437),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__557 (
            .O(N__4430),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    CascadeMux I__556 (
            .O(N__4425),
            .I(N__4421));
    CascadeMux I__555 (
            .O(N__4424),
            .I(N__4417));
    InMux I__554 (
            .O(N__4421),
            .I(N__4410));
    InMux I__553 (
            .O(N__4420),
            .I(N__4410));
    InMux I__552 (
            .O(N__4417),
            .I(N__4403));
    InMux I__551 (
            .O(N__4416),
            .I(N__4403));
    InMux I__550 (
            .O(N__4415),
            .I(N__4403));
    LocalMux I__549 (
            .O(N__4410),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__548 (
            .O(N__4403),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    CascadeMux I__547 (
            .O(N__4398),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_1_cascade_ ));
    CascadeMux I__546 (
            .O(N__4395),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_2_cascade_ ));
    CascadeMux I__545 (
            .O(N__4392),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_0_cascade_ ));
    CascadeMux I__544 (
            .O(N__4389),
            .I(N__4383));
    CascadeMux I__543 (
            .O(N__4388),
            .I(N__4380));
    InMux I__542 (
            .O(N__4387),
            .I(N__4377));
    InMux I__541 (
            .O(N__4386),
            .I(N__4372));
    InMux I__540 (
            .O(N__4383),
            .I(N__4372));
    InMux I__539 (
            .O(N__4380),
            .I(N__4369));
    LocalMux I__538 (
            .O(N__4377),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__537 (
            .O(N__4372),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__536 (
            .O(N__4369),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    CascadeMux I__535 (
            .O(N__4362),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_a2_0_4_cascade_ ));
    InMux I__534 (
            .O(N__4359),
            .I(N__4356));
    LocalMux I__533 (
            .O(N__4356),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_a2_0_1 ));
    CascadeMux I__532 (
            .O(N__4353),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_ ));
    CascadeMux I__531 (
            .O(N__4350),
            .I(\U712_CHIP_RAM.N_43_cascade_ ));
    InMux I__530 (
            .O(N__4347),
            .I(N__4344));
    LocalMux I__529 (
            .O(N__4344),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6 ));
    InMux I__528 (
            .O(N__4341),
            .I(N__4332));
    InMux I__527 (
            .O(N__4340),
            .I(N__4332));
    InMux I__526 (
            .O(N__4339),
            .I(N__4332));
    LocalMux I__525 (
            .O(N__4332),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4 ));
    CascadeMux I__524 (
            .O(N__4329),
            .I(\U712_REG_SM.N_162_0_cascade_ ));
    InMux I__523 (
            .O(N__4326),
            .I(N__4320));
    InMux I__522 (
            .O(N__4325),
            .I(N__4320));
    LocalMux I__521 (
            .O(N__4320),
            .I(\U712_REG_SM.N_172_0 ));
    CascadeMux I__520 (
            .O(N__4317),
            .I(N__4311));
    InMux I__519 (
            .O(N__4316),
            .I(N__4308));
    InMux I__518 (
            .O(N__4315),
            .I(N__4303));
    InMux I__517 (
            .O(N__4314),
            .I(N__4303));
    InMux I__516 (
            .O(N__4311),
            .I(N__4300));
    LocalMux I__515 (
            .O(N__4308),
            .I(\U712_REG_SM.N_162_0 ));
    LocalMux I__514 (
            .O(N__4303),
            .I(\U712_REG_SM.N_162_0 ));
    LocalMux I__513 (
            .O(N__4300),
            .I(\U712_REG_SM.N_162_0 ));
    InMux I__512 (
            .O(N__4293),
            .I(N__4289));
    InMux I__511 (
            .O(N__4292),
            .I(N__4286));
    LocalMux I__510 (
            .O(N__4289),
            .I(\U712_REG_SM.N_195 ));
    LocalMux I__509 (
            .O(N__4286),
            .I(\U712_REG_SM.N_195 ));
    CascadeMux I__508 (
            .O(N__4281),
            .I(\U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_ ));
    InMux I__507 (
            .O(N__4278),
            .I(N__4274));
    InMux I__506 (
            .O(N__4277),
            .I(N__4271));
    LocalMux I__505 (
            .O(N__4274),
            .I(N__4264));
    LocalMux I__504 (
            .O(N__4271),
            .I(N__4264));
    InMux I__503 (
            .O(N__4270),
            .I(N__4259));
    InMux I__502 (
            .O(N__4269),
            .I(N__4259));
    Odrv4 I__501 (
            .O(N__4264),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    LocalMux I__500 (
            .O(N__4259),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    CascadeMux I__499 (
            .O(N__4254),
            .I(N__4251));
    InMux I__498 (
            .O(N__4251),
            .I(N__4245));
    InMux I__497 (
            .O(N__4250),
            .I(N__4245));
    LocalMux I__496 (
            .O(N__4245),
            .I(\U712_REG_SM.C1_SYNCZ0Z_2 ));
    InMux I__495 (
            .O(N__4242),
            .I(N__4235));
    InMux I__494 (
            .O(N__4241),
            .I(N__4232));
    InMux I__493 (
            .O(N__4240),
            .I(N__4227));
    InMux I__492 (
            .O(N__4239),
            .I(N__4227));
    InMux I__491 (
            .O(N__4238),
            .I(N__4224));
    LocalMux I__490 (
            .O(N__4235),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__489 (
            .O(N__4232),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__488 (
            .O(N__4227),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    LocalMux I__487 (
            .O(N__4224),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    CascadeMux I__486 (
            .O(N__4215),
            .I(N__4211));
    InMux I__485 (
            .O(N__4214),
            .I(N__4206));
    InMux I__484 (
            .O(N__4211),
            .I(N__4203));
    InMux I__483 (
            .O(N__4210),
            .I(N__4200));
    InMux I__482 (
            .O(N__4209),
            .I(N__4197));
    LocalMux I__481 (
            .O(N__4206),
            .I(N__4192));
    LocalMux I__480 (
            .O(N__4203),
            .I(N__4192));
    LocalMux I__479 (
            .O(N__4200),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__478 (
            .O(N__4197),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__477 (
            .O(N__4192),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    InMux I__476 (
            .O(N__4185),
            .I(N__4178));
    InMux I__475 (
            .O(N__4184),
            .I(N__4178));
    InMux I__474 (
            .O(N__4183),
            .I(N__4175));
    LocalMux I__473 (
            .O(N__4178),
            .I(\U712_REG_SM.N_163_0 ));
    LocalMux I__472 (
            .O(N__4175),
            .I(\U712_REG_SM.N_163_0 ));
    InMux I__471 (
            .O(N__4170),
            .I(N__4166));
    InMux I__470 (
            .O(N__4169),
            .I(N__4163));
    LocalMux I__469 (
            .O(N__4166),
            .I(N__4160));
    LocalMux I__468 (
            .O(N__4163),
            .I(\U712_REG_SM.N_194 ));
    Odrv4 I__467 (
            .O(N__4160),
            .I(\U712_REG_SM.N_194 ));
    InMux I__466 (
            .O(N__4155),
            .I(N__4152));
    LocalMux I__465 (
            .O(N__4152),
            .I(N__4147));
    InMux I__464 (
            .O(N__4151),
            .I(N__4142));
    InMux I__463 (
            .O(N__4150),
            .I(N__4142));
    Odrv4 I__462 (
            .O(N__4147),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    LocalMux I__461 (
            .O(N__4142),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_6 ));
    IoInMux I__460 (
            .O(N__4137),
            .I(N__4134));
    LocalMux I__459 (
            .O(N__4134),
            .I(N__4130));
    IoInMux I__458 (
            .O(N__4133),
            .I(N__4127));
    IoSpan4Mux I__457 (
            .O(N__4130),
            .I(N__4124));
    LocalMux I__456 (
            .O(N__4127),
            .I(N__4121));
    Sp12to4 I__455 (
            .O(N__4124),
            .I(N__4118));
    IoSpan4Mux I__454 (
            .O(N__4121),
            .I(N__4115));
    Span12Mux_v I__453 (
            .O(N__4118),
            .I(N__4112));
    Sp12to4 I__452 (
            .O(N__4115),
            .I(N__4109));
    Span12Mux_h I__451 (
            .O(N__4112),
            .I(N__4104));
    Span12Mux_v I__450 (
            .O(N__4109),
            .I(N__4104));
    Odrv12 I__449 (
            .O(N__4104),
            .I(ASn_c));
    CEMux I__448 (
            .O(N__4101),
            .I(N__4098));
    LocalMux I__447 (
            .O(N__4098),
            .I(N__4095));
    Span4Mux_v I__446 (
            .O(N__4095),
            .I(N__4092));
    Odrv4 I__445 (
            .O(N__4092),
            .I(\U712_REG_SM.N_186_0 ));
    IoInMux I__444 (
            .O(N__4089),
            .I(N__4086));
    LocalMux I__443 (
            .O(N__4086),
            .I(N__4083));
    Span12Mux_s10_h I__442 (
            .O(N__4083),
            .I(N__4080));
    Odrv12 I__441 (
            .O(N__4080),
            .I(N_510_i));
    IoInMux I__440 (
            .O(N__4077),
            .I(N__4074));
    LocalMux I__439 (
            .O(N__4074),
            .I(N__4071));
    Span12Mux_s8_v I__438 (
            .O(N__4071),
            .I(N__4068));
    Odrv12 I__437 (
            .O(N__4068),
            .I(VBENn_c));
    CascadeMux I__436 (
            .O(N__4065),
            .I(\U712_REG_SM.N_175_cascade_ ));
    InMux I__435 (
            .O(N__4062),
            .I(N__4059));
    LocalMux I__434 (
            .O(N__4059),
            .I(N__4056));
    Odrv4 I__433 (
            .O(N__4056),
            .I(\U712_REG_SM.N_171_0 ));
    CascadeMux I__432 (
            .O(N__4053),
            .I(\U712_REG_SM.N_194_cascade_ ));
    CascadeMux I__431 (
            .O(N__4050),
            .I(N__4045));
    InMux I__430 (
            .O(N__4049),
            .I(N__4038));
    InMux I__429 (
            .O(N__4048),
            .I(N__4038));
    InMux I__428 (
            .O(N__4045),
            .I(N__4038));
    LocalMux I__427 (
            .O(N__4038),
            .I(\U712_REG_SM.N_169_0 ));
    InMux I__426 (
            .O(N__4035),
            .I(N__4029));
    InMux I__425 (
            .O(N__4034),
            .I(N__4029));
    LocalMux I__424 (
            .O(N__4029),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_1 ));
    CascadeMux I__423 (
            .O(N__4026),
            .I(\U712_REG_SM.N_170_0_cascade_ ));
    CascadeMux I__422 (
            .O(N__4023),
            .I(\U712_REG_SM.N_174_cascade_ ));
    InMux I__421 (
            .O(N__4020),
            .I(N__4016));
    InMux I__420 (
            .O(N__4019),
            .I(N__4013));
    LocalMux I__419 (
            .O(N__4016),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__418 (
            .O(N__4013),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__417 (
            .O(N__4008),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__416 (
            .O(N__4005),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    InMux I__415 (
            .O(N__4002),
            .I(N__3998));
    InMux I__414 (
            .O(N__4001),
            .I(N__3995));
    LocalMux I__413 (
            .O(N__3998),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    LocalMux I__412 (
            .O(N__3995),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    ClkMux I__411 (
            .O(N__3990),
            .I(N__3987));
    GlobalMux I__410 (
            .O(N__3987),
            .I(N__3984));
    gio2CtrlBuf I__409 (
            .O(N__3984),
            .I(C1_c_g));
    CascadeMux I__408 (
            .O(N__3981),
            .I(N__3977));
    InMux I__407 (
            .O(N__3980),
            .I(N__3973));
    InMux I__406 (
            .O(N__3977),
            .I(N__3970));
    InMux I__405 (
            .O(N__3976),
            .I(N__3967));
    LocalMux I__404 (
            .O(N__3973),
            .I(N__3964));
    LocalMux I__403 (
            .O(N__3970),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    LocalMux I__402 (
            .O(N__3967),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    Odrv4 I__401 (
            .O(N__3964),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_0 ));
    CascadeMux I__400 (
            .O(N__3957),
            .I(N__3953));
    InMux I__399 (
            .O(N__3956),
            .I(N__3949));
    InMux I__398 (
            .O(N__3953),
            .I(N__3945));
    InMux I__397 (
            .O(N__3952),
            .I(N__3942));
    LocalMux I__396 (
            .O(N__3949),
            .I(N__3939));
    InMux I__395 (
            .O(N__3948),
            .I(N__3936));
    LocalMux I__394 (
            .O(N__3945),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__393 (
            .O(N__3942),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    Odrv4 I__392 (
            .O(N__3939),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__391 (
            .O(N__3936),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    CascadeMux I__390 (
            .O(N__3927),
            .I(\U712_REG_SM.N_168_0_cascade_ ));
    CascadeMux I__389 (
            .O(N__3924),
            .I(N__3920));
    CascadeMux I__388 (
            .O(N__3923),
            .I(N__3917));
    InMux I__387 (
            .O(N__3920),
            .I(N__3909));
    InMux I__386 (
            .O(N__3917),
            .I(N__3909));
    InMux I__385 (
            .O(N__3916),
            .I(N__3909));
    LocalMux I__384 (
            .O(N__3909),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_2 ));
    InMux I__383 (
            .O(N__3906),
            .I(N__3903));
    LocalMux I__382 (
            .O(N__3903),
            .I(N__3900));
    Span4Mux_v I__381 (
            .O(N__3900),
            .I(N__3897));
    Sp12to4 I__380 (
            .O(N__3897),
            .I(N__3894));
    Span12Mux_h I__379 (
            .O(N__3894),
            .I(N__3891));
    Odrv12 I__378 (
            .O(N__3891),
            .I(C3_c));
    CascadeMux I__377 (
            .O(N__3888),
            .I(\U712_CHIP_RAM.REFRESH_r_1_cascade_ ));
    InMux I__376 (
            .O(N__3885),
            .I(N__3882));
    LocalMux I__375 (
            .O(N__3882),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ));
    InMux I__374 (
            .O(N__3879),
            .I(bfn_7_7_0_));
    InMux I__373 (
            .O(N__3876),
            .I(N__3873));
    LocalMux I__372 (
            .O(N__3873),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    InMux I__371 (
            .O(N__3870),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__370 (
            .O(N__3867),
            .I(N__3863));
    InMux I__369 (
            .O(N__3866),
            .I(N__3860));
    LocalMux I__368 (
            .O(N__3863),
            .I(\U712_CHIP_RAM.REFRESH6lto2 ));
    LocalMux I__367 (
            .O(N__3860),
            .I(\U712_CHIP_RAM.REFRESH6lto2 ));
    InMux I__366 (
            .O(N__3855),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__365 (
            .O(N__3852),
            .I(N__3848));
    InMux I__364 (
            .O(N__3851),
            .I(N__3845));
    LocalMux I__363 (
            .O(N__3848),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__362 (
            .O(N__3845),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__361 (
            .O(N__3840),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__360 (
            .O(N__3837),
            .I(N__3833));
    InMux I__359 (
            .O(N__3836),
            .I(N__3830));
    LocalMux I__358 (
            .O(N__3833),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__357 (
            .O(N__3830),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__356 (
            .O(N__3825),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    CascadeMux I__355 (
            .O(N__3822),
            .I(N__3818));
    InMux I__354 (
            .O(N__3821),
            .I(N__3815));
    InMux I__353 (
            .O(N__3818),
            .I(N__3812));
    LocalMux I__352 (
            .O(N__3815),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__351 (
            .O(N__3812),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    InMux I__350 (
            .O(N__3807),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    IoInMux I__349 (
            .O(N__3804),
            .I(N__3801));
    LocalMux I__348 (
            .O(N__3801),
            .I(N__3798));
    Span4Mux_s2_v I__347 (
            .O(N__3798),
            .I(N__3795));
    Span4Mux_v I__346 (
            .O(N__3795),
            .I(N__3792));
    Odrv4 I__345 (
            .O(N__3792),
            .I(CLK80_OUT_i_i));
    IoInMux I__344 (
            .O(N__3789),
            .I(N__3786));
    LocalMux I__343 (
            .O(N__3786),
            .I(N__3783));
    Odrv12 I__342 (
            .O(N__3783),
            .I(CLK40_OUT_i_i));
    InMux I__341 (
            .O(N__3780),
            .I(N__3777));
    LocalMux I__340 (
            .O(N__3777),
            .I(N__3774));
    Span4Mux_v I__339 (
            .O(N__3774),
            .I(N__3771));
    Span4Mux_h I__338 (
            .O(N__3771),
            .I(N__3768));
    Sp12to4 I__337 (
            .O(N__3768),
            .I(N__3765));
    Span12Mux_v I__336 (
            .O(N__3765),
            .I(N__3762));
    Odrv12 I__335 (
            .O(N__3762),
            .I(REGSPACEn_c));
    CascadeMux I__334 (
            .O(N__3759),
            .I(\U712_REG_SM.un6_REG_CYCLE_START_cascade_ ));
    InMux I__333 (
            .O(N__3756),
            .I(N__3752));
    InMux I__332 (
            .O(N__3755),
            .I(N__3749));
    LocalMux I__331 (
            .O(N__3752),
            .I(\U712_REG_SM.REG_CYCLE_GOZ0 ));
    LocalMux I__330 (
            .O(N__3749),
            .I(\U712_REG_SM.REG_CYCLE_GOZ0 ));
    InMux I__329 (
            .O(N__3744),
            .I(N__3741));
    LocalMux I__328 (
            .O(N__3741),
            .I(N__3737));
    IoInMux I__327 (
            .O(N__3740),
            .I(N__3734));
    Span4Mux_v I__326 (
            .O(N__3737),
            .I(N__3731));
    LocalMux I__325 (
            .O(N__3734),
            .I(N__3728));
    Sp12to4 I__324 (
            .O(N__3731),
            .I(N__3725));
    Span4Mux_s3_h I__323 (
            .O(N__3728),
            .I(N__3722));
    Span12Mux_h I__322 (
            .O(N__3725),
            .I(N__3717));
    Sp12to4 I__321 (
            .O(N__3722),
            .I(N__3717));
    Span12Mux_v I__320 (
            .O(N__3717),
            .I(N__3714));
    Odrv12 I__319 (
            .O(N__3714),
            .I(C1_c));
    IoInMux I__318 (
            .O(N__3711),
            .I(N__3708));
    LocalMux I__317 (
            .O(N__3708),
            .I(N__3705));
    IoSpan4Mux I__316 (
            .O(N__3705),
            .I(N__3702));
    Span4Mux_s2_v I__315 (
            .O(N__3702),
            .I(N__3699));
    Sp12to4 I__314 (
            .O(N__3699),
            .I(N__3696));
    Span12Mux_v I__313 (
            .O(N__3696),
            .I(N__3693));
    Odrv12 I__312 (
            .O(N__3693),
            .I(CLK40_IN_c));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__7812),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__3740),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_2_1_1.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_2_1_1.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_2_1_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 CLKRAM_obuf_RNO_LC_2_1_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9537),
            .lcout(CLK80_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CLK40C_obuf_RNO_LC_3_10_3.C_ON=1'b0;
    defparam CLK40C_obuf_RNO_LC_3_10_3.SEQ_MODE=4'b0000;
    defparam CLK40C_obuf_RNO_LC_3_10_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLK40C_obuf_RNO_LC_3_10_3 (
            .in0(N__5076),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_OUT_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_10_6 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_10_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(N__3755),
            .in2(_gnd_net_),
            .in3(N__3952),
            .lcout(),
            .ltout(\U712_REG_SM.un6_REG_CYCLE_START_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_6_10_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_6_10_7 .LUT_INIT=16'b1010000010100010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_6_10_7  (
            .in0(N__7996),
            .in1(N__3780),
            .in2(N__3759),
            .in3(N__4836),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9524),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_6_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_GO_LC_6_11_3 .LUT_INIT=16'b1010000011101100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_GO_LC_6_11_3  (
            .in0(N__3976),
            .in1(N__3756),
            .in2(N__3957),
            .in3(N__4673),
            .lcout(\U712_REG_SM.REG_CYCLE_GOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9527),
            .ce(),
            .sr(N__9293));
    defparam \U712_REG_SM.C3_SYNC_1_LC_6_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_6_12_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_6_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4278),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9530),
            .ce(),
            .sr(N__9284));
    defparam \U712_REG_SM.C1_SYNC_0_LC_6_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_6_12_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_6_12_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_6_12_5  (
            .in0(N__3744),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9530),
            .ce(),
            .sr(N__9284));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_6_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_6_12_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_6_12_6 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_6_12_6  (
            .in0(N__3956),
            .in1(N__4316),
            .in2(N__3981),
            .in3(N__4293),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9530),
            .ce(),
            .sr(N__9284));
    defparam \U712_REG_SM.C1_SYNC_2_LC_6_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_2_LC_6_13_5 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_2_LC_6_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_2_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4210),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9531),
            .ce(),
            .sr(N__9277));
    defparam \U712_REG_SM.C1_SYNC_1_LC_6_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_6_13_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_6_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4242),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9531),
            .ce(),
            .sr(N__9277));
    defparam \U712_REG_SM.C3_SYNC_0_LC_6_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_6_14_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_6_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_6_14_1  (
            .in0(N__3906),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9533),
            .ce(),
            .sr(N__9270));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_7_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_7_6_1 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_7_6_1  (
            .in0(N__3836),
            .in1(N__3851),
            .in2(N__3822),
            .in3(N__3866),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH_r_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_7_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_7_6_2 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_7_6_2  (
            .in0(N__8007),
            .in1(N__4001),
            .in2(N__3888),
            .in3(N__4019),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9510),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__3885),
            .in2(_gnd_net_),
            .in3(N__3879),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__3990),
            .ce(),
            .sr(N__5523));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__3876),
            .in2(_gnd_net_),
            .in3(N__3870),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__3990),
            .ce(),
            .sr(N__5523));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__3867),
            .in2(_gnd_net_),
            .in3(N__3855),
            .lcout(\U712_CHIP_RAM.REFRESH6lto2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__3990),
            .ce(),
            .sr(N__5523));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__3852),
            .in2(_gnd_net_),
            .in3(N__3840),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__3990),
            .ce(),
            .sr(N__5523));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__3837),
            .in2(_gnd_net_),
            .in3(N__3825),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__3990),
            .ce(),
            .sr(N__5523));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__3821),
            .in2(_gnd_net_),
            .in3(N__3807),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__3990),
            .ce(),
            .sr(N__5523));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__4020),
            .in2(_gnd_net_),
            .in3(N__4008),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__3990),
            .ce(),
            .sr(N__5523));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(N__4002),
            .in2(_gnd_net_),
            .in3(N__4005),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__3990),
            .ce(),
            .sr(N__5523));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_10_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__3980),
            .in2(_gnd_net_),
            .in3(N__3948),
            .lcout(\U712_REG_SM.N_171_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_7_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_0_LC_7_11_0 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_0_LC_7_11_0  (
            .in0(N__6971),
            .in1(N__4277),
            .in2(_gnd_net_),
            .in3(N__4241),
            .lcout(\U712_REG_SM.DS_EN_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_7_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_7_11_1 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_7_11_1  (
            .in0(N__4672),
            .in1(N__7898),
            .in2(N__3924),
            .in3(N__4049),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9525),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_4_LC_7_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_4_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_4_LC_7_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_4_LC_7_11_2  (
            .in0(N__5366),
            .in1(N__6593),
            .in2(N__6501),
            .in3(N__4490),
            .lcout(),
            .ltout(\U712_REG_SM.N_168_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_7_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_7_11_3 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_7_11_3  (
            .in0(N__4470),
            .in1(N__7900),
            .in2(N__3927),
            .in3(N__4452),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9525),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_7_11_4 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DS_EN_RNO_1_LC_7_11_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_REG_SM.DS_EN_RNO_1_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4050),
            .in3(N__3916),
            .lcout(\U712_REG_SM.N_187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_7_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_7_11_5 .LUT_INIT=16'b0000001111110011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__5365),
            .in2(N__3923),
            .in3(N__4048),
            .lcout(),
            .ltout(\U712_REG_SM.N_175_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_7_11_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_7_11_6 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_7_11_6  (
            .in0(N__7899),
            .in1(_gnd_net_),
            .in2(N__4065),
            .in3(N__5349),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9525),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_7_12_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_7_12_0 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_7_12_0  (
            .in0(N__8002),
            .in1(N__4062),
            .in2(N__4674),
            .in3(N__4035),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9528),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNICU4F1_1_LC_7_12_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNICU4F1_1_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNICU4F1_1_LC_7_12_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNICU4F1_1_LC_7_12_1  (
            .in0(N__4510),
            .in1(N__4544),
            .in2(N__4215),
            .in3(N__4238),
            .lcout(\U712_REG_SM.N_194 ),
            .ltout(\U712_REG_SM.N_194_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_7_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_7_12_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNISG3L1_6_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4053),
            .in3(N__4150),
            .lcout(\U712_REG_SM.N_195 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_7_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_7_12_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_0_2_LC_7_12_3  (
            .in0(N__4512),
            .in1(N__4560),
            .in2(_gnd_net_),
            .in3(N__4546),
            .lcout(\U712_REG_SM.N_169_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_7_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_7_12_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIKD9V_1_LC_7_12_4  (
            .in0(N__4545),
            .in1(N__4034),
            .in2(_gnd_net_),
            .in3(N__4511),
            .lcout(\U712_REG_SM.N_172_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_7_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_7_12_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_1_2_LC_7_12_5  (
            .in0(N__4314),
            .in1(N__4183),
            .in2(N__4522),
            .in3(N__4547),
            .lcout(\U712_REG_SM.N_170_0 ),
            .ltout(\U712_REG_SM.N_170_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_7_12_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_7_12_6 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_7_12_6  (
            .in0(_gnd_net_),
            .in1(N__5394),
            .in2(N__4026),
            .in3(N__4151),
            .lcout(),
            .ltout(\U712_REG_SM.N_174_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_7_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_7_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_7_12_7 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_7_12_7  (
            .in0(N__4315),
            .in1(N__8003),
            .in2(N__4023),
            .in3(N__4169),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9528),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_7_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_7_13_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI6FIN_2_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__4270),
            .in2(_gnd_net_),
            .in3(N__4250),
            .lcout(\U712_REG_SM.N_162_0 ),
            .ltout(\U712_REG_SM.N_162_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_7_13_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_7_13_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_7_13_2  (
            .in0(N__4185),
            .in1(_gnd_net_),
            .in2(N__4329),
            .in3(N__4326),
            .lcout(\U712_REG_SM.N_173_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_7_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_7_13_4 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIPBP14_1_LC_7_13_4  (
            .in0(N__4184),
            .in1(N__4325),
            .in2(N__4317),
            .in3(N__4292),
            .lcout(\U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1 ),
            .ltout(\U712_REG_SM.STATE_COUNT_RNIPBP14Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_1_ess_RNO_LC_7_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_1_ess_RNO_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REGENn_1_ess_RNO_LC_7_13_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_REG_SM.REGENn_1_ess_RNO_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4281),
            .in3(N__9355),
            .lcout(\U712_REG_SM.N_186_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_7_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_7_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_7_13_6  (
            .in0(N__4269),
            .in1(N__4209),
            .in2(N__4254),
            .in3(N__4239),
            .lcout(\U712_REG_SM.N_157_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_7_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_7_13_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_REG_SM.C1_SYNC_RNI3UPL_1_LC_7_13_7  (
            .in0(N__4240),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4214),
            .lcout(\U712_REG_SM.N_163_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_1_ess_LC_7_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_1_ess_LC_7_14_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_1_ess_LC_7_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_REG_SM.REGENn_1_ess_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__4170),
            .in2(_gnd_net_),
            .in3(N__4155),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9532),
            .ce(N__4101),
            .sr(N__9265));
    defparam TACKn_obuft_RNO_LC_7_15_6.C_ON=1'b0;
    defparam TACKn_obuft_RNO_LC_7_15_6.SEQ_MODE=4'b0000;
    defparam TACKn_obuft_RNO_LC_7_15_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 TACKn_obuft_RNO_LC_7_15_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6801),
            .lcout(N_510_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_LC_8_5_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_LC_8_5_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_BUFFERS.un1_VBENn_LC_8_5_2  (
            .in0(_gnd_net_),
            .in1(N__7185),
            .in2(_gnd_net_),
            .in3(N__8298),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_8_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_8_5_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_8_5_7  (
            .in0(N__6242),
            .in1(N__5916),
            .in2(N__6162),
            .in3(N__5632),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_6_0 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_6_0  (
            .in0(N__4751),
            .in1(N__9364),
            .in2(N__4424),
            .in3(N__4341),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9503),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_4_LC_8_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_4_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_4_LC_8_6_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_4_LC_8_6_1  (
            .in0(N__4339),
            .in1(N__4416),
            .in2(_gnd_net_),
            .in3(N__4749),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_6_2 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(N__9365),
            .in2(N__4353),
            .in3(N__4443),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9503),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_6_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_8_6_3  (
            .in0(N__4442),
            .in1(N__4415),
            .in2(N__4388),
            .in3(N__4748),
            .lcout(\U712_CHIP_RAM.N_43 ),
            .ltout(\U712_CHIP_RAM.N_43_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_8_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_8_6_4 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI74LA2_0_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4350),
            .in3(N__5915),
            .lcout(\U712_CHIP_RAM.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_6_5 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_6_5  (
            .in0(N__4444),
            .in1(N__4347),
            .in2(N__9369),
            .in3(N__4387),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9503),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_6_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_6_6  (
            .in0(N__4750),
            .in1(N__9363),
            .in2(_gnd_net_),
            .in3(N__4340),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9503),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_6_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_8_6_7  (
            .in0(N__4898),
            .in1(N__6161),
            .in2(N__6263),
            .in3(N__5735),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_0_LC_8_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_0_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_0_LC_8_7_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5RIP2_0_LC_8_7_0  (
            .in0(N__5616),
            .in1(N__5913),
            .in2(_gnd_net_),
            .in3(N__4712),
            .lcout(\U712_CHIP_RAM.N_100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3EPC1_5_LC_8_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3EPC1_5_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI3EPC1_5_LC_8_7_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI3EPC1_5_LC_8_7_1  (
            .in0(N__4445),
            .in1(N__4420),
            .in2(_gnd_net_),
            .in3(N__5615),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_7_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_7_2  (
            .in0(N__4386),
            .in1(N__4446),
            .in2(N__4425),
            .in3(N__4731),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_7_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_7_3  (
            .in0(N__6009),
            .in1(_gnd_net_),
            .in2(N__4398),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_7_4 .LUT_INIT=16'b0110000000100000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_7_4  (
            .in0(N__5617),
            .in1(N__5914),
            .in2(N__4395),
            .in3(N__6256),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_7_5 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_8_7_5  (
            .in0(N__4869),
            .in1(N__7995),
            .in2(N__4392),
            .in3(N__5095),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9511),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6F3C2_7_LC_8_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6F3C2_7_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6F3C2_7_LC_8_7_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6F3C2_7_LC_8_7_6  (
            .in0(N__6238),
            .in1(N__4730),
            .in2(N__4389),
            .in3(N__6008),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_a2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAB4_5_LC_8_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAB4_5_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAB4_5_LC_8_7_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAB4_5_LC_8_7_7  (
            .in0(N__4868),
            .in1(_gnd_net_),
            .in2(N__4362),
            .in3(N__4359),
            .lcout(\U712_CHIP_RAM.N_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBDIR_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_8_8_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_8_8_0 .LUT_INIT=16'b0111001011110000;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_8_8_0  (
            .in0(N__6047),
            .in1(N__7010),
            .in2(N__5008),
            .in3(N__6179),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9514),
            .ce(),
            .sr(N__9301));
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_8_1 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_8_8_1  (
            .in0(N__6178),
            .in1(N__6046),
            .in2(_gnd_net_),
            .in3(N__4799),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_8_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_LC_8_8_2 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_LC_8_8_2  (
            .in0(N__5965),
            .in1(N__6905),
            .in2(N__4611),
            .in3(N__8272),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9514),
            .ce(),
            .sr(N__9301));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_10_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_10_5 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_8_10_5 .LUT_INIT=16'b1111100011111010;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_8_10_5  (
            .in0(N__4595),
            .in1(N__5072),
            .in2(N__5145),
            .in3(N__6564),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9521),
            .ce(),
            .sr(N__9285));
    defparam \U712_REG_SM.DS_EN_LC_8_11_0 .C_ON=1'b0;
    defparam \U712_REG_SM.DS_EN_LC_8_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.DS_EN_LC_8_11_0 .LUT_INIT=16'b0000111100101110;
    LogicCell40 \U712_REG_SM.DS_EN_LC_8_11_0  (
            .in0(N__7265),
            .in1(N__4584),
            .in2(N__4575),
            .in3(N__4566),
            .lcout(\U712_REG_SM.DS_ENZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9522),
            .ce(),
            .sr(N__9278));
    defparam \U712_REG_SM.C3_SYNC_2_LC_8_11_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_2_LC_8_11_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_2_LC_8_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_2_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4527),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9522),
            .ce(),
            .sr(N__9278));
    defparam \U712_REG_SM.REG_TACK_LC_8_11_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_8_11_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_8_11_5 .LUT_INIT=16'b1011101010111000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_8_11_5  (
            .in0(N__4469),
            .in1(N__5397),
            .in2(N__5118),
            .in3(N__4491),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9522),
            .ce(),
            .sr(N__9278));
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_8_12_2 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_8_12_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_RNI3QN13_1_LC_8_12_2  (
            .in0(N__4489),
            .in1(N__6594),
            .in2(_gnd_net_),
            .in3(N__6500),
            .lcout(\U712_REG_SM.N_167_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_8_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_8_12_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_8_12_3  (
            .in0(N__4559),
            .in1(N__4548),
            .in2(_gnd_net_),
            .in3(N__4523),
            .lcout(\U712_REG_SM.N_159_0 ),
            .ltout(\U712_REG_SM.N_159_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI0ULC2_4_LC_8_12_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI0ULC2_4_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI0ULC2_4_LC_8_12_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI0ULC2_4_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4473),
            .in3(N__4468),
            .lcout(\U712_REG_SM.N_165_0 ),
            .ltout(\U712_REG_SM.N_165_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_8_12_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_8_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_8_12_5 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_8_12_5  (
            .in0(N__7981),
            .in1(N__5395),
            .in2(N__4683),
            .in3(N__4680),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9526),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDS_OUT_LC_8_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.UDS_OUT_LC_8_13_1 .LUT_INIT=16'b1111010111001100;
    LogicCell40 \U712_REG_SM.UDS_OUT_LC_8_13_1  (
            .in0(N__4632),
            .in1(N__7289),
            .in2(N__6964),
            .in3(N__4671),
            .lcout(\U712_REG_SM.UDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9529),
            .ce(),
            .sr(N__9266));
    defparam \U712_REG_SM.LDS_OUT_LC_8_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.LDS_OUT_LC_8_13_6 .LUT_INIT=16'b1111011110100010;
    LogicCell40 \U712_REG_SM.LDS_OUT_LC_8_13_6  (
            .in0(N__4670),
            .in1(N__4638),
            .in2(N__6963),
            .in3(N__6383),
            .lcout(\U712_REG_SM.LDS_OUTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9529),
            .ce(),
            .sr(N__9266));
    defparam \U712_REG_SM.LDS_OUT_RNO_0_LC_8_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_RNO_0_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_RNO_0_LC_8_14_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_REG_SM.LDS_OUT_RNO_0_LC_8_14_4  (
            .in0(N__5221),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5290),
            .lcout(\U712_REG_SM.LDS_OUT_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.UDS_OUT_RNO_0_LC_8_14_5 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_RNO_0_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDS_OUT_RNO_0_LC_8_14_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \U712_REG_SM.UDS_OUT_RNO_0_LC_8_14_5  (
            .in0(N__5291),
            .in1(N__5222),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.UDS_OUT_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_9_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_9_5_1 .LUT_INIT=16'b0000000011001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_9_5_1  (
            .in0(N__6243),
            .in1(N__4899),
            .in2(N__6155),
            .in3(N__5734),
            .lcout(\U712_CHIP_RAM.N_105 ),
            .ltout(\U712_CHIP_RAM.N_105_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI264TB_LC_9_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI264TB_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI264TB_LC_9_5_2 .LUT_INIT=16'b1111001011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI264TB_LC_9_5_2  (
            .in0(N__5747),
            .in1(N__5670),
            .in2(N__4626),
            .in3(N__5952),
            .lcout(\U712_CHIP_RAM.N_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_5_3 .LUT_INIT=16'b0001110100010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_5_3  (
            .in0(N__5953),
            .in1(N__5697),
            .in2(N__5681),
            .in3(N__4722),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_cnst_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_5_4 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__8001),
            .in2(N__4623),
            .in3(N__4620),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_5_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_5_5  (
            .in0(N__5496),
            .in1(_gnd_net_),
            .in2(N__4614),
            .in3(N__8640),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9494),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_LC_9_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_LC_9_5_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRCRT_0_LC_9_5_6  (
            .in0(N__5634),
            .in1(_gnd_net_),
            .in2(N__5922),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(N__5918),
            .in2(_gnd_net_),
            .in3(N__5633),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_9_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_9_6_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_3_LC_9_6_1  (
            .in0(N__6233),
            .in1(N__6125),
            .in2(_gnd_net_),
            .in3(N__4711),
            .lcout(\U712_CHIP_RAM.N_50 ),
            .ltout(\U712_CHIP_RAM.N_50_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_9_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_9_6_2 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_9_6_2  (
            .in0(N__5901),
            .in1(_gnd_net_),
            .in2(N__4716),
            .in3(N__5629),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRB433_2_LC_9_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRB433_2_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIRB433_2_LC_9_6_3 .LUT_INIT=16'b0000111101011110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIRB433_2_LC_9_6_3  (
            .in0(N__5630),
            .in1(N__6048),
            .in2(N__6257),
            .in3(N__5902),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_0_tz_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIT32E6_3_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIT32E6_3_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIT32E6_3_LC_9_6_4 .LUT_INIT=16'b0001000011111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIT32E6_3_LC_9_6_4  (
            .in0(N__6126),
            .in1(N__4713),
            .in2(N__4695),
            .in3(N__5777),
            .lcout(),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHPUTC_3_LC_9_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHPUTC_3_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIHPUTC_3_LC_9_6_5 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIHPUTC_3_LC_9_6_5  (
            .in0(N__4785),
            .in1(N__8000),
            .in2(N__4692),
            .in3(N__4764),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_6_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_9_6_6  (
            .in0(N__7999),
            .in1(N__4689),
            .in2(_gnd_net_),
            .in3(N__5736),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9497),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_6_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_9_6_7  (
            .in0(N__6237),
            .in1(N__5477),
            .in2(_gnd_net_),
            .in3(N__5801),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9497),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMMGI5_2_LC_9_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMMGI5_2_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMMGI5_2_LC_9_7_0 .LUT_INIT=16'b1111111100000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIMMGI5_2_LC_9_7_0  (
            .in0(N__5757),
            .in1(N__6241),
            .in2(N__6015),
            .in3(N__4763),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIP5G8C_2_LC_9_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIP5G8C_2_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIP5G8C_2_LC_9_7_1 .LUT_INIT=16'b1110101011101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIP5G8C_2_LC_9_7_1  (
            .in0(N__4800),
            .in1(N__4784),
            .in2(N__4773),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_57_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIM9IMI_0_LC_9_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIM9IMI_0_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIM9IMI_0_LC_9_7_2 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIM9IMI_0_LC_9_7_2  (
            .in0(N__9362),
            .in1(N__5976),
            .in2(N__4770),
            .in3(N__5954),
            .lcout(\U712_CHIP_RAM.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_3_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_3_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_3_LC_9_7_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_3_LC_9_7_3  (
            .in0(N__6239),
            .in1(N__5618),
            .in2(N__6148),
            .in3(N__5693),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_92_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN7BL3_LC_9_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN7BL3_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN7BL3_LC_9_7_4 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN7BL3_LC_9_7_4  (
            .in0(N__5756),
            .in1(N__6240),
            .in2(N__4767),
            .in3(N__5732),
            .lcout(\U712_CHIP_RAM.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_4_LC_9_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_4_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_4_LC_9_7_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI1JRT_4_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__6127),
            .in2(_gnd_net_),
            .in3(N__4752),
            .lcout(\U712_CHIP_RAM.BANK0_0_sqmuxa_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_7_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_7_6  (
            .in0(N__5619),
            .in1(N__5887),
            .in2(_gnd_net_),
            .in3(N__5800),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9504),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_9_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_9_7_7 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_9_7_7  (
            .in0(N__5731),
            .in1(N__6318),
            .in2(_gnd_net_),
            .in3(N__6294),
            .lcout(\U712_CHIP_RAM.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_9_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_9_8_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_9_8_1  (
            .in0(N__5680),
            .in1(N__6006),
            .in2(N__5917),
            .in3(N__5620),
            .lcout(\U712_CHIP_RAM.N_106 ),
            .ltout(\U712_CHIP_RAM.N_106_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7Q5U5_0_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7Q5U5_0_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI7Q5U5_0_LC_9_8_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI7Q5U5_0_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4935),
            .in3(N__6037),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_3_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_3_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_3_LC_9_8_3 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIDD06A_3_LC_9_8_3  (
            .in0(N__6275),
            .in1(N__6258),
            .in2(N__4932),
            .in3(N__6157),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_9_8_4 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_9_8_4 .LUT_INIT=16'b1010110011111100;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_9_8_4  (
            .in0(N__5911),
            .in1(N__5413),
            .in2(N__4929),
            .in3(N__7023),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9512),
            .ce(),
            .sr(N__9294));
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_8_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_LC_9_8_5 .LUT_INIT=16'b1011111110110000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_LC_9_8_5  (
            .in0(N__6864),
            .in1(N__5912),
            .in2(N__6081),
            .in3(N__4910),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9512),
            .ce(),
            .sr(N__9294));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI72V93_0_LC_9_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI72V93_0_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI72V93_0_LC_9_8_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI72V93_0_LC_9_8_6  (
            .in0(N__6007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4894),
            .lcout(\U712_CHIP_RAM.N_70_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_9_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_LC_9_8_7 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_LC_9_8_7  (
            .in0(N__7214),
            .in1(N__5966),
            .in2(N__4878),
            .in3(N__6906),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9512),
            .ce(),
            .sr(N__9294));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJDDI_0_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJDDI_0_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIJDDI_0_LC_9_9_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIJDDI_0_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__5857),
            .in2(_gnd_net_),
            .in3(N__8239),
            .lcout(\U712_CHIP_RAM.CPU_TACK_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_1  (
            .in0(N__8240),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6070),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un6_CPU_CYCLE_START_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_2 .LUT_INIT=16'b1100000011000100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_2  (
            .in0(N__4857),
            .in1(N__7967),
            .in2(N__4839),
            .in3(N__4832),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9515),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_10_0 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_9_10_0  (
            .in0(N__7963),
            .in1(N__5124),
            .in2(N__5071),
            .in3(N__6818),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9517),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_10_1 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__7965),
            .in2(_gnd_net_),
            .in3(N__5031),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9517),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_10_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_9_10_2  (
            .in0(N__7966),
            .in1(_gnd_net_),
            .in2(N__5144),
            .in3(_gnd_net_),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9517),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_10_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_10_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__5137),
            .in2(_gnd_net_),
            .in3(N__5030),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_10_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_10_4 .LUT_INIT=16'b0000000000110111;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_10_4  (
            .in0(N__5097),
            .in1(N__6817),
            .in2(N__5117),
            .in3(N__6561),
            .lcout(\U712_CYCLE_TERM.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_10_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN6_LC_9_10_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN6_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__5110),
            .in2(_gnd_net_),
            .in3(N__5096),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(\U712_CYCLE_TERM.TACK_EN6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_6 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_10_6  (
            .in0(N__7962),
            .in1(N__6539),
            .in2(N__5079),
            .in3(N__6816),
            .lcout(\U712_CYCLE_TERM.N_45_0_0_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_10_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_9_10_7  (
            .in0(N__6562),
            .in1(N__7964),
            .in2(_gnd_net_),
            .in3(N__5064),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9517),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_0_i_LC_9_11_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_0_i_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_0_i_LC_9_11_1 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \U712_BUFFERS.DRDDIR_0_i_LC_9_11_1  (
            .in0(N__7171),
            .in1(N__6972),
            .in2(N__7238),
            .in3(N__5015),
            .lcout(DRDDIR_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_LC_9_11_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_LC_9_11_2 .LUT_INIT=16'b1101000011011101;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_LC_9_11_2  (
            .in0(N__5466),
            .in1(N__7344),
            .in2(N__5328),
            .in3(N__8324),
            .lcout(CLMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un3_CLLBEn_1_LC_9_11_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un3_CLLBEn_1_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un3_CLLBEn_1_LC_9_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_BYTE_ENABLE.un3_CLLBEn_1_LC_9_11_3  (
            .in0(N__7233),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5422),
            .lcout(\U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1 ),
            .ltout(\U712_BYTE_ENABLE.un3_CLLBEnZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_LC_9_11_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_LC_9_11_4 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_LC_9_11_4  (
            .in0(N__7378),
            .in1(N__5337),
            .in2(N__5460),
            .in3(N__8323),
            .lcout(CLLBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un3_CUMBEn_0_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un3_CUMBEn_0_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un3_CUMBEn_0_LC_9_11_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_BYTE_ENABLE.un3_CUMBEn_0_LC_9_11_7  (
            .in0(N__7234),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5423),
            .lcout(\U712_BYTE_ENABLE.un3_CUMBEnZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_9_12_3 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_9_12_3 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_9_12_3  (
            .in0(N__5396),
            .in1(N__7170),
            .in2(N__5373),
            .in3(N__5348),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9523),
            .ce(),
            .sr(N__9267));
    defparam \U712_BYTE_ENABLE.LLBE_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_LC_9_13_0 .LUT_INIT=16'b0001010100100010;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_LC_9_13_0  (
            .in0(N__5182),
            .in1(N__5263),
            .in2(N__5234),
            .in3(N__5314),
            .lcout(\U712_BYTE_ENABLE.LLBE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.LMBE_LC_9_13_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LMBE_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LMBE_LC_9_13_4 .LUT_INIT=16'b0101000110100010;
    LogicCell40 \U712_BYTE_ENABLE.LMBE_LC_9_13_4  (
            .in0(N__5183),
            .in1(N__5264),
            .in2(N__5235),
            .in3(N__5315),
            .lcout(\U712_BYTE_ENABLE.LMBE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_LC_9_13_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_LC_9_13_7 .LUT_INIT=16'b0110000001100100;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_LC_9_13_7  (
            .in0(N__5190),
            .in1(N__5316),
            .in2(N__5268),
            .in3(N__5232),
            .lcout(\U712_BYTE_ENABLE.UMBE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UUBE_LC_9_14_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UUBE_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UUBE_LC_9_14_2 .LUT_INIT=16'b0101010010101000;
    LogicCell40 \U712_BYTE_ENABLE.UUBE_LC_9_14_2  (
            .in0(N__5313),
            .in1(N__5262),
            .in2(N__5233),
            .in3(N__5181),
            .lcout(\U712_BYTE_ENABLE.UUBE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_4_3 .LUT_INIT=16'b0000000001100111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_10_4_3  (
            .in0(N__8615),
            .in1(N__8835),
            .in2(N__8987),
            .in3(N__8537),
            .lcout(\U712_CHIP_RAM.un1_CMA31_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_4_6 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_10_4_6  (
            .in0(N__6609),
            .in1(N__8616),
            .in2(N__8375),
            .in3(N__8019),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_4_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_4_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_10_4_7  (
            .in0(N__8346),
            .in1(N__5559),
            .in2(N__5541),
            .in3(N__5538),
            .lcout(\U712_CHIP_RAM.N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_5_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_10_5_0  (
            .in0(N__8834),
            .in1(N__8962),
            .in2(N__8641),
            .in3(N__8535),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_5_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_5_2  (
            .in0(N__7994),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5504),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_78_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_5_3 .LUT_INIT=16'b1010101000000011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_5_3  (
            .in0(N__8536),
            .in1(N__5763),
            .in2(N__5511),
            .in3(N__5495),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9488),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_5_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_5_5  (
            .in0(N__5679),
            .in1(N__5748),
            .in2(_gnd_net_),
            .in3(N__7993),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_76_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_5_6 .LUT_INIT=16'b1010101100000001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_5_6  (
            .in0(N__5494),
            .in1(N__5784),
            .in2(N__5508),
            .in3(N__8963),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9488),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_5_7 .LUT_INIT=16'b1111000001110111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_5_7  (
            .in0(N__5505),
            .in1(N__7992),
            .in2(N__8881),
            .in3(N__5493),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9488),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_6_0 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_10_6_0  (
            .in0(N__6129),
            .in1(N__5478),
            .in2(N__6264),
            .in3(N__5802),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9495),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_6_1  (
            .in0(N__5778),
            .in1(N__5614),
            .in2(N__5682),
            .in3(N__6860),
            .lcout(\U712_CHIP_RAM.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_10_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_10_6_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_10_6_2  (
            .in0(N__7991),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6010),
            .lcout(\U712_CHIP_RAM.N_99 ),
            .ltout(\U712_CHIP_RAM.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_6_3 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_6_3  (
            .in0(N__5677),
            .in1(_gnd_net_),
            .in2(N__5766),
            .in3(N__5613),
            .lcout(\U712_CHIP_RAM.N_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_6_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIUFRT_3_LC_10_6_5  (
            .in0(_gnd_net_),
            .in1(N__6128),
            .in2(_gnd_net_),
            .in3(N__5611),
            .lcout(\U712_CHIP_RAM.N_93_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_6_6 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_6_6  (
            .in0(N__8836),
            .in1(N__8633),
            .in2(_gnd_net_),
            .in3(N__8967),
            .lcout(\U712_CHIP_RAM.CMA_5_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMT791_LC_10_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMT791_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMT791_LC_10_6_7 .LUT_INIT=16'b1000100001010101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIMT791_LC_10_6_7  (
            .in0(N__5897),
            .in1(N__5612),
            .in2(_gnd_net_),
            .in3(N__5733),
            .lcout(\U712_CHIP_RAM.N_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_10_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_10_7_0 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_10_7_0  (
            .in0(N__5730),
            .in1(N__6316),
            .in2(_gnd_net_),
            .in3(N__6291),
            .lcout(\U712_CHIP_RAM.N_54 ),
            .ltout(\U712_CHIP_RAM.N_54_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_10_7_1 .LUT_INIT=16'b0000001000000001;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_RNO_1_LC_10_7_1  (
            .in0(N__5886),
            .in1(N__5678),
            .in2(N__5637),
            .in3(N__5631),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNO_0_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNO_0_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_RNO_0_LC_10_7_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_RNO_0_LC_10_7_2  (
            .in0(N__6333),
            .in1(N__6072),
            .in2(_gnd_net_),
            .in3(N__8357),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH_CYCLE_START_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_10_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_10_7_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_10_7_3  (
            .in0(N__7229),
            .in1(N__6904),
            .in2(N__6321),
            .in3(N__7998),
            .lcout(\U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9498),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_10_7_6 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_RNO_0_LC_10_7_6  (
            .in0(N__5961),
            .in1(N__6317),
            .in2(_gnd_net_),
            .in3(N__6292),
            .lcout(),
            .ltout(\U712_CHIP_RAM.REFRESH_CYCLE_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_CYCLE_LC_10_7_7 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_CYCLE_LC_10_7_7  (
            .in0(N__6293),
            .in1(N__7997),
            .in2(N__6303),
            .in3(N__6300),
            .lcout(\U712_CHIP_RAM.REFRESH_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9498),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_8_2 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_RNO_0_LC_10_8_2  (
            .in0(N__6276),
            .in1(N__6259),
            .in2(N__6180),
            .in3(N__6156),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER53_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_8_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_8_4  (
            .in0(N__6586),
            .in1(N__6894),
            .in2(N__6071),
            .in3(N__6493),
            .lcout(\U712_CHIP_RAM.N_40 ),
            .ltout(\U712_CHIP_RAM.N_40_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_10_8_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNI3EN62_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6018),
            .in3(N__6011),
            .lcout(\U712_CHIP_RAM.N_59 ),
            .ltout(\U712_CHIP_RAM.N_59_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_8_6 .LUT_INIT=16'b0001000101010100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_8_6  (
            .in0(N__9359),
            .in1(N__5888),
            .in2(N__5970),
            .in3(N__5967),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9505),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_10_9_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_10_9_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_10_9_2  (
            .in0(N__9357),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5808),
            .lcout(\U712_CYCLE_TERM.N_45_0_0_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_9_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__9356),
            .in2(_gnd_net_),
            .in3(N__6600),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.DBR_SYNC_1_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_10_10_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.DBR_SYNC_1_LC_10_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.DBR_SYNC_1_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6492),
            .lcout(U712_REG_SM_DBR_SYNC_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9516),
            .ce(),
            .sr(N__9271));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_10_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_10_6 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_10_10_6 .LUT_INIT=16'b0101010001010000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_10_10_6  (
            .in0(N__6563),
            .in1(N__6830),
            .in2(N__6543),
            .in3(N__6528),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9516),
            .ce(),
            .sr(N__9271));
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_10_11_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_10_11_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBR_SYNC_0_LC_10_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DBR_SYNC_0_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6522),
            .lcout(U712_REG_SM_DBR_SYNC_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9518),
            .ce(),
            .sr(N__9268));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_LC_10_12_2 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_LC_10_12_2 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_LC_10_12_2  (
            .in0(N__6419),
            .in1(N__7386),
            .in2(N__8391),
            .in3(N__6462),
            .lcout(CUMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_LC_10_12_5 .LUT_INIT=16'b1100010011110101;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_LC_10_12_5  (
            .in0(N__8390),
            .in1(N__7337),
            .in2(N__6432),
            .in3(N__6420),
            .lcout(CUUBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_10_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDS_OUT_RNIL31J_LC_10_14_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.LDS_OUT_RNIL31J_LC_10_14_0  (
            .in0(N__6390),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7277),
            .lcout(U712_REG_SM_un1_LDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_11_3_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_11_3_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_11_3_5 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_11_3_5  (
            .in0(N__8890),
            .in1(N__9005),
            .in2(_gnd_net_),
            .in3(N__6639),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9479),
            .ce(N__9081),
            .sr(N__9313));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_3_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_11_3_6 .LUT_INIT=16'b1010101010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_11_3_6  (
            .in0(N__6765),
            .in1(_gnd_net_),
            .in2(N__9021),
            .in3(N__8891),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9479),
            .ce(N__9081),
            .sr(N__9313));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_4_3 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_11_4_3  (
            .in0(N__6747),
            .in1(N__6633),
            .in2(N__6729),
            .in3(N__8345),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_35_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_11_4_4 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_11_4_4  (
            .in0(N__8854),
            .in1(_gnd_net_),
            .in2(N__6705),
            .in3(N__8986),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9482),
            .ce(N__9064),
            .sr(N__9310));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_4_5 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_4_5  (
            .in0(N__6618),
            .in1(N__8343),
            .in2(N__8710),
            .in3(N__8415),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_4_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_11_4_6  (
            .in0(N__8344),
            .in1(N__6678),
            .in2(N__6660),
            .in3(N__6657),
            .lcout(\U712_CHIP_RAM.N_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_5_1 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_11_5_1  (
            .in0(N__7494),
            .in1(N__8377),
            .in2(N__6627),
            .in3(N__8666),
            .lcout(\U712_CHIP_RAM.CMA_5_3_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_11_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_11_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_11_6_0  (
            .in0(N__7487),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9489),
            .ce(N__7409),
            .sr(N__9295));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_11_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_11_6_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_11_6_2  (
            .in0(N__7517),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9489),
            .ce(N__7409),
            .sr(N__9295));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_11_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_11_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8454),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9489),
            .ce(N__7409),
            .sr(N__9295));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_11_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_11_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8055),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9489),
            .ce(N__7409),
            .sr(N__9295));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_11_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_11_7_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__9358),
            .in2(_gnd_net_),
            .in3(N__6779),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESS4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_7_6 .LUT_INIT=16'b0000001111110101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_11_7_6  (
            .in0(N__7065),
            .in1(N__9144),
            .in2(N__8378),
            .in3(N__8694),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_7_7  (
            .in0(N__8356),
            .in1(N__7059),
            .in2(N__7041),
            .in3(N__7038),
            .lcout(\U712_CHIP_RAM.N_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DBENn_RNO_0_LC_11_8_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.DBENn_RNO_0_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__7425),
            .in2(_gnd_net_),
            .in3(N__6895),
            .lcout(\U712_CHIP_RAM.DBENn_7_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_8_5 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_11_8_5  (
            .in0(N__7225),
            .in1(N__6896),
            .in2(N__6783),
            .in3(N__7982),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9499),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_11_9_3 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_11_9_3  (
            .in0(N__7014),
            .in1(N__6962),
            .in2(_gnd_net_),
            .in3(N__6903),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9506),
            .ce(N__6843),
            .sr(N__9272));
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_11_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_EN_i_ess_LC_11_10_0 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_i_ess_LC_11_10_0  (
            .in0(N__7937),
            .in1(N__6834),
            .in2(_gnd_net_),
            .in3(N__6819),
            .lcout(TACK_EN_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9513),
            .ce(N__6789),
            .sr(N__9269));
    defparam \U712_CHIP_RAM.CAS_SYNC_RNILUVG_1_LC_11_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNILUVG_1_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_SYNC_RNILUVG_1_LC_11_11_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_RNILUVG_1_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(N__7299),
            .in2(_gnd_net_),
            .in3(N__7310),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESS4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_12_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_12_1 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_11_12_1  (
            .in0(N__7385),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7336),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9519),
            .ce(),
            .sr(N__9264));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_12_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_11_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7311),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9519),
            .ce(),
            .sr(N__9264));
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_11_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDS_OUT_RNIUP9B_LC_11_13_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \U712_REG_SM.UDS_OUT_RNIUP9B_LC_11_13_1  (
            .in0(N__7293),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7278),
            .lcout(U712_REG_SM_un1_UDSn_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_DRDENn_LC_11_13_2 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_DRDENn_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_DRDENn_LC_11_13_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_DRDENn_LC_11_13_2  (
            .in0(N__7239),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7184),
            .lcout(DRDENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_4_3 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_12_4_3  (
            .in0(N__7419),
            .in1(N__8373),
            .in2(N__8709),
            .in3(N__7449),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_4_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_4_4  (
            .in0(N__8374),
            .in1(N__7110),
            .in2(N__7092),
            .in3(N__7089),
            .lcout(\U712_CHIP_RAM.N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_4_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_4_6  (
            .in0(N__9360),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7074),
            .lcout(\U712_CHIP_RAM.un1_CMA31_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7518),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9481),
            .ce(N__8774),
            .sr(N__9292));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7488),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9481),
            .ce(N__8774),
            .sr(N__9292));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_12_6_1 .LUT_INIT=16'b1110111100000001;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_12_6_1  (
            .in0(N__8897),
            .in1(N__9019),
            .in2(N__8718),
            .in3(N__7443),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9484),
            .ce(N__9080),
            .sr(N__9283));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_12_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_12_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_12_7_0  (
            .in0(N__8097),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9487),
            .ce(N__7410),
            .sr(N__9276));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_12_7_1  (
            .in0(N__9171),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9487),
            .ce(N__7410),
            .sr(N__9276));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_12_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_12_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_12_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8126),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9487),
            .ce(N__7410),
            .sr(N__9276));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_12_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_12_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_12_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_12_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8487),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9487),
            .ce(N__7410),
            .sr(N__9276));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_12_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_12_7_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_12_7_7  (
            .in0(N__8169),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9487),
            .ce(N__7410),
            .sr(N__9276));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_5 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_8_5  (
            .in0(N__7392),
            .in1(N__8314),
            .in2(N__8698),
            .in3(N__8460),
            .lcout(\U712_CHIP_RAM.CMA_5_3_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_0.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_0.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7897),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_3_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_3_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_13_3_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_13_3_0  (
            .in0(N__7698),
            .in1(N__8895),
            .in2(_gnd_net_),
            .in3(N__9018),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9480),
            .ce(N__9096),
            .sr(N__9314));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_3_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_3_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_13_3_3 .LUT_INIT=16'b1110111100000001;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_13_3_3  (
            .in0(N__9017),
            .in1(N__8896),
            .in2(N__8714),
            .in3(N__7785),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9480),
            .ce(N__9096),
            .sr(N__9314));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_4_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_4_3 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_13_4_3  (
            .in0(N__7755),
            .in1(N__8369),
            .in2(N__8716),
            .in3(N__8064),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_4_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_4_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_4_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_4_4  (
            .in0(N__8370),
            .in1(N__7746),
            .in2(N__7725),
            .in3(N__7722),
            .lcout(\U712_CHIP_RAM.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_5_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_5_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_13_5_1 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_13_5_1  (
            .in0(N__7692),
            .in1(N__7635),
            .in2(N__8142),
            .in3(N__8379),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9485),
            .ce(N__9091),
            .sr(N__9302));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_6_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_13_6_4  (
            .in0(N__7524),
            .in1(N__8901),
            .in2(_gnd_net_),
            .in3(N__9020),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9490),
            .ce(N__9095),
            .sr(N__9296));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_13_6_6 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_13_6_6  (
            .in0(N__9585),
            .in1(N__7634),
            .in2(N__7614),
            .in3(N__8380),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9490),
            .ce(N__9095),
            .sr(N__9296));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_4 .LUT_INIT=16'b1110001000110011;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_4  (
            .in0(N__7575),
            .in1(N__7554),
            .in2(N__7548),
            .in3(N__8376),
            .lcout(\U712_CHIP_RAM.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_8_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_8_1  (
            .in0(N__8483),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9500),
            .ce(N__8765),
            .sr(N__9279));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_8_4  (
            .in0(N__8450),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9500),
            .ce(N__8765),
            .sr(N__9279));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_14_4_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_14_4_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_14_4_5 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_14_4_5  (
            .in0(N__8403),
            .in1(N__8371),
            .in2(N__8715),
            .in3(N__8103),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_5_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_4_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_4_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_4_6 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_4_6  (
            .in0(N__8372),
            .in1(N__8202),
            .in2(N__8187),
            .in3(N__8184),
            .lcout(\U712_CHIP_RAM.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_5_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_5_3  (
            .in0(N__8168),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9491),
            .ce(N__8775),
            .sr(N__9311));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_5_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_5_4  (
            .in0(N__8133),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9491),
            .ce(N__8775),
            .sr(N__9311));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_6_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_6_4  (
            .in0(N__8093),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9496),
            .ce(N__8770),
            .sr(N__9303));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8048),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9496),
            .ce(N__8770),
            .sr(N__9303));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9167),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9501),
            .ce(N__8769),
            .sr(N__9297));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_4_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_4_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_15_4_1 .LUT_INIT=16'b1100100011001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_15_4_1  (
            .in0(N__8899),
            .in1(N__9135),
            .in2(N__9030),
            .in3(_gnd_net_),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9492),
            .ce(N__9065),
            .sr(N__9318));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_15_4_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_15_4_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_15_4_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_15_4_3  (
            .in0(N__8898),
            .in1(N__8708),
            .in2(N__9029),
            .in3(N__8550),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9492),
            .ce(N__9065),
            .sr(N__9318));
    defparam \U712_CHIP_RAM.WEn_LC_16_1_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_16_1_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_16_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_16_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9028),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9483),
            .ce(),
            .sr(N__9321));
    defparam \U712_CHIP_RAM.RASn_LC_16_3_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_16_3_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_16_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_16_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8900),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9493),
            .ce(),
            .sr(N__9319));
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_8_2 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_16_8_2  (
            .in0(N__9361),
            .in1(N__9543),
            .in2(_gnd_net_),
            .in3(N__9554),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESS5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_17_1_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_17_1_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_17_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_17_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8717),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9486),
            .ce(),
            .sr(N__9322));
    defparam \U712_CHIP_RAM.CRCSn_LC_17_4_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_17_4_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_17_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_17_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8549),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9502),
            .ce(),
            .sr(N__9320));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_8_2 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_8_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_17_8_2  (
            .in0(N__8499),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9581),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9520),
            .ce(),
            .sr(N__9312));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_17_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_17_8_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_17_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9555),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__9520),
            .ce(),
            .sr(N__9312));
endmodule // U712_TOP
